-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     Jun 1 2022 09:54:43

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : inout std_logic_vector(15 downto 0);
    port_data : inout std_logic_vector(7 downto 0);
    debug : out std_logic_vector(1 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    led : out std_logic_vector(7 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : inout std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__44416\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44377\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44296\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44287\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44125\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44107\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44027\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44008\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43999\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43989\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43906\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43731\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43692\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43659\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43653\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43548\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43503\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43440\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43326\ : std_logic;
signal \N__43323\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43197\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43191\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43061\ : std_logic;
signal \N__43058\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43049\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42750\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42732\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42544\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42541\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42520\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42496\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42415\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42407\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42398\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42355\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42304\ : std_logic;
signal \N__42301\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42211\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42130\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42124\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42107\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42059\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42056\ : std_logic;
signal \N__42055\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41644\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41421\ : std_logic;
signal \N__41418\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41398\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41386\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41152\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41134\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41131\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40816\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40727\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40677\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40452\ : std_logic;
signal \N__40449\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40207\ : std_logic;
signal \N__40204\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40180\ : std_logic;
signal \N__40177\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39871\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39784\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39461\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39250\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38608\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38063\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37020\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35263\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \VCCG0\ : std_logic;
signal \this_vga_signals.N_1307_0\ : std_logic;
signal \N_428\ : std_logic;
signal \N_842\ : std_logic;
signal rgb_c_4 : std_logic;
signal \M_vcounter_q_esr_RNIQ82H7_9\ : std_logic;
signal \M_this_oam_ram_read_data_13\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_13\ : std_logic;
signal rgb_c_2 : std_logic;
signal rgb_c_5 : std_logic;
signal \this_ppu.oam_cache.N_561_0\ : std_logic;
signal \this_ppu.oam_cache.mem_17\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_17\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_16\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_17\ : std_logic;
signal \M_this_ppu_spr_addr_4\ : std_logic;
signal \this_ppu.offset_y_cry_0\ : std_logic;
signal \this_ppu.offset_y_cry_1\ : std_logic;
signal \M_this_ppu_spr_addr_5\ : std_logic;
signal \this_ppu.oam_cache.mem_16\ : std_logic;
signal \this_ppu.oam_cache.mem_18\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_18\ : std_logic;
signal port_clk_c : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_0\ : std_logic;
signal \M_this_oam_ram_read_data_12\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_12\ : std_logic;
signal \this_ppu.oam_cache.N_579_0\ : std_logic;
signal \M_this_oam_ram_read_data_26\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_26\ : std_logic;
signal \N_84\ : std_logic;
signal rgb_c_0 : std_logic;
signal \M_this_oam_ram_read_data_15\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_15\ : std_logic;
signal \this_ppu.oam_cache.N_577_0\ : std_logic;
signal \this_ppu.oam_cache.N_567_0\ : std_logic;
signal \M_this_oam_ram_read_data_8\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_8\ : std_logic;
signal \M_this_oam_ram_read_data_9\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_9\ : std_logic;
signal \M_this_oam_ram_read_data_10\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_10\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_16\ : std_logic;
signal \this_ppu.oam_cache.mem_4\ : std_logic;
signal \this_ppu.N_985_0\ : std_logic;
signal \this_ppu.N_671_0\ : std_logic;
signal \this_ppu.N_426_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_oam_curr_q_1_c2_cascade_\ : std_logic;
signal \this_ppu.N_986_0\ : std_logic;
signal \this_ppu.un1_M_oam_curr_q_1_c4_cascade_\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_cascade_\ : std_logic;
signal \this_ppu.N_841_0\ : std_logic;
signal \this_ppu.N_841_0_cascade_\ : std_logic;
signal \this_ppu.N_669_0\ : std_logic;
signal \this_ppu.m18_i_o2_1_cascade_\ : std_logic;
signal \this_ppu.N_426_0\ : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal \this_ppu.oam_cache.mem_2\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_21\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_22\ : std_logic;
signal \M_this_oam_ram_read_data_3\ : std_logic;
signal \M_this_oam_ram_read_data_6\ : std_logic;
signal \M_this_oam_ram_read_data_25\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_25\ : std_logic;
signal \M_this_warmup_qZ0Z_1\ : std_logic;
signal \M_this_warmup_qZ0Z_0\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \M_this_warmup_qZ0Z_2\ : std_logic;
signal \un1_M_this_warmup_d_cry_1\ : std_logic;
signal \M_this_warmup_qZ0Z_3\ : std_logic;
signal \un1_M_this_warmup_d_cry_2\ : std_logic;
signal \M_this_warmup_qZ0Z_4\ : std_logic;
signal \un1_M_this_warmup_d_cry_3\ : std_logic;
signal \M_this_warmup_qZ0Z_5\ : std_logic;
signal \un1_M_this_warmup_d_cry_4\ : std_logic;
signal \M_this_warmup_qZ0Z_6\ : std_logic;
signal \un1_M_this_warmup_d_cry_5\ : std_logic;
signal \M_this_warmup_qZ0Z_7\ : std_logic;
signal \un1_M_this_warmup_d_cry_6\ : std_logic;
signal \M_this_warmup_qZ0Z_8\ : std_logic;
signal \un1_M_this_warmup_d_cry_7\ : std_logic;
signal \un1_M_this_warmup_d_cry_8\ : std_logic;
signal \M_this_warmup_qZ0Z_9\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \M_this_warmup_qZ0Z_10\ : std_logic;
signal \un1_M_this_warmup_d_cry_9\ : std_logic;
signal \M_this_warmup_qZ0Z_11\ : std_logic;
signal \un1_M_this_warmup_d_cry_10\ : std_logic;
signal \M_this_warmup_qZ0Z_12\ : std_logic;
signal \un1_M_this_warmup_d_cry_11\ : std_logic;
signal \M_this_warmup_qZ0Z_13\ : std_logic;
signal \un1_M_this_warmup_d_cry_12\ : std_logic;
signal \M_this_warmup_qZ0Z_14\ : std_logic;
signal \un1_M_this_warmup_d_cry_13\ : std_logic;
signal \M_this_warmup_qZ0Z_15\ : std_logic;
signal \un1_M_this_warmup_d_cry_14\ : std_logic;
signal \M_this_warmup_qZ0Z_16\ : std_logic;
signal \un1_M_this_warmup_d_cry_15\ : std_logic;
signal \un1_M_this_warmup_d_cry_16\ : std_logic;
signal \M_this_warmup_qZ0Z_17\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \M_this_warmup_qZ0Z_18\ : std_logic;
signal \un1_M_this_warmup_d_cry_17\ : std_logic;
signal \M_this_warmup_qZ0Z_19\ : std_logic;
signal \un1_M_this_warmup_d_cry_18\ : std_logic;
signal \M_this_warmup_qZ0Z_20\ : std_logic;
signal \un1_M_this_warmup_d_cry_19\ : std_logic;
signal \M_this_warmup_qZ0Z_21\ : std_logic;
signal \un1_M_this_warmup_d_cry_20\ : std_logic;
signal \M_this_warmup_qZ0Z_22\ : std_logic;
signal \un1_M_this_warmup_d_cry_21\ : std_logic;
signal \M_this_warmup_qZ0Z_23\ : std_logic;
signal \un1_M_this_warmup_d_cry_22\ : std_logic;
signal \M_this_warmup_qZ0Z_24\ : std_logic;
signal \un1_M_this_warmup_d_cry_23\ : std_logic;
signal \un1_M_this_warmup_d_cry_24\ : std_logic;
signal \M_this_warmup_qZ0Z_25\ : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal \M_this_warmup_qZ0Z_26\ : std_logic;
signal \un1_M_this_warmup_d_cry_25\ : std_logic;
signal \un1_M_this_warmup_d_cry_26\ : std_logic;
signal \M_this_warmup_qZ0Z_27\ : std_logic;
signal \M_this_oam_ram_write_data_18\ : std_logic;
signal \M_this_oam_ram_write_data_23\ : std_logic;
signal \M_this_oam_ram_write_data_20\ : std_logic;
signal \M_this_oam_ram_write_data_19\ : std_logic;
signal \M_this_oam_ram_write_data_17\ : std_logic;
signal rgb_c_1 : std_logic;
signal \M_this_oam_ram_read_data_0\ : std_logic;
signal \this_ppu.oam_cache.N_586_0\ : std_logic;
signal \this_ppu.oam_cache.mem_10\ : std_logic;
signal \this_ppu.N_844_0\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_10\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_0\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_1\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_2\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_3\ : std_logic;
signal \this_ppu.oam_cache.mem_7\ : std_logic;
signal \N_41_0\ : std_logic;
signal \M_this_ppu_oam_addr_1\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_qZ0Z_4\ : std_logic;
signal \this_ppu.m62_0_a2_0_o2_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_oam_curr_q_1_c4\ : std_logic;
signal \this_ppu.M_oam_curr_qc_0_1\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_CO\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_qZ0Z_1\ : std_logic;
signal \this_ppu.m62_0_a2_0_o2_1\ : std_logic;
signal \M_this_ppu_oam_addr_3\ : std_logic;
signal \M_this_ppu_oam_addr_2\ : std_logic;
signal \M_this_ppu_oam_addr_4\ : std_logic;
signal \this_ppu.un1_M_oam_curr_q_1_c2\ : std_logic;
signal \this_ppu.un1_M_oam_curr_q_1_c5\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_CO\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_qZ0Z_3\ : std_logic;
signal \M_this_oam_ram_read_data_24\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_24\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_1\ : std_logic;
signal \M_this_oam_ram_read_data_7\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.haddress_1_0\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m2\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3\ : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb1\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_qZ1Z_0\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal \M_this_oam_ram_read_data_16\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_i_16\ : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_i_17\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_0\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_i_18\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_1\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_2\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_3\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_4\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_5\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_3_c_RNIT7IDZ0\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_2_c_RNIR4HDZ0\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_6\ : std_logic;
signal \this_ppu.m28_e_i_o3_2\ : std_logic;
signal \M_this_oam_ram_read_data_18\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_18\ : std_logic;
signal \M_this_oam_ram_write_data_5\ : std_logic;
signal \M_this_oam_ram_read_data_22\ : std_logic;
signal \M_this_oam_ram_read_data_i_22\ : std_logic;
signal \M_this_oam_ram_read_data_29\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_29\ : std_logic;
signal \M_this_oam_ram_read_data_21\ : std_logic;
signal \M_this_oam_ram_read_data_i_21\ : std_logic;
signal \M_this_oam_ram_read_data_31\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_31\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_19\ : std_logic;
signal \M_this_oam_ram_read_data_19\ : std_logic;
signal \M_this_oam_ram_read_data_i_19\ : std_logic;
signal \M_this_oam_ram_write_data_10\ : std_logic;
signal \N_260\ : std_logic;
signal \M_this_oam_ram_read_data_28\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_28\ : std_logic;
signal \M_this_oam_ram_write_data_9\ : std_logic;
signal \M_this_oam_ram_read_data_i_20\ : std_logic;
signal \M_this_oam_ram_write_data_28\ : std_logic;
signal \M_this_oam_ram_write_data_8\ : std_logic;
signal \M_this_oam_ram_write_data_31\ : std_logic;
signal \M_this_oam_ram_write_data_16\ : std_logic;
signal \M_this_oam_ram_write_data_24\ : std_logic;
signal \this_vga_signals.hsync_1_i_0_0_1\ : std_logic;
signal \M_this_oam_ram_read_data_14\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_14\ : std_logic;
signal \this_vga_signals.hsync_1_i_0_0_a3_0_0\ : std_logic;
signal \this_vga_signals.N_811_0\ : std_logic;
signal rgb_c_3 : std_logic;
signal \M_this_ppu_oam_addr_5\ : std_logic;
signal \M_this_ppu_oam_addr_0\ : std_logic;
signal \this_ppu.m35_i_0_a3_1_3\ : std_logic;
signal \this_ppu.N_1394\ : std_logic;
signal \M_this_oam_ram_read_data_2\ : std_logic;
signal \this_ppu.m28_e_i_a3_4\ : std_logic;
signal \this_ppu.m28_e_i_a3_3\ : std_logic;
signal \this_ppu.N_1184_7_cascade_\ : std_logic;
signal \this_ppu.m18_i_1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0_2\ : std_logic;
signal \this_ppu.oam_cache.mem_12\ : std_logic;
signal \M_this_oam_ram_read_data_5\ : std_logic;
signal \this_ppu.oam_cache.N_569_0\ : std_logic;
signal \M_this_oam_ram_read_data_4\ : std_logic;
signal \this_ppu.oam_cache.N_575_0\ : std_logic;
signal \this_ppu.N_1182\ : std_logic;
signal \this_vga_signals.if_N_9_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c2_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_8_i\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_2\ : std_logic;
signal \M_this_oam_ram_read_data_27\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_27\ : std_logic;
signal \this_ppu.oam_cache.mem_0\ : std_logic;
signal \this_ppu.un1_oam_data_1_axb_7\ : std_logic;
signal \M_this_oam_ram_write_data_6\ : std_logic;
signal \M_this_data_tmp_qZ0Z_6\ : std_logic;
signal \M_this_oam_ram_write_data_7\ : std_logic;
signal \M_this_data_tmp_qZ0Z_7\ : std_logic;
signal \M_this_oam_ram_read_data_17\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_17\ : std_logic;
signal \M_this_data_tmp_qZ0Z_10\ : std_logic;
signal \M_this_data_tmp_qZ0Z_8\ : std_logic;
signal \M_this_data_tmp_qZ0Z_9\ : std_logic;
signal \M_this_oam_ram_write_data_26\ : std_logic;
signal \M_this_oam_ram_write_data_27\ : std_logic;
signal \M_this_oam_ram_write_data_30\ : std_logic;
signal \M_this_data_tmp_qZ0Z_15\ : std_logic;
signal \M_this_oam_ram_write_data_15\ : std_logic;
signal \M_this_data_tmp_qZ0Z_16\ : std_logic;
signal \M_this_data_tmp_qZ0Z_17\ : std_logic;
signal \M_this_data_tmp_qZ0Z_19\ : std_logic;
signal \M_this_data_tmp_qZ0Z_20\ : std_logic;
signal \M_this_data_tmp_qZ0Z_18\ : std_logic;
signal \M_this_oam_ram_write_data_0\ : std_logic;
signal \this_vga_ramdac.N_852_i_reto\ : std_logic;
signal \this_vga_signals.N_298_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_d7_0_i_0_o3_0_o3_4_a2_0\ : std_logic;
signal \this_vga_signals.N_1044_0_cascade_\ : std_logic;
signal \this_vga_signals.N_298_0\ : std_logic;
signal \this_vga_signals.hsync_1_i_0_0_a3_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_3_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_0_0_tz\ : std_logic;
signal \this_ppu.N_1184_7\ : std_logic;
signal \this_ppu.un1_M_state_q_7_i_0\ : std_logic;
signal \M_this_oam_ram_read_data_11\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_11\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_12\ : std_logic;
signal \this_ppu.oam_cache.mem_15\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.N_968\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.N_968_cascade_\ : std_logic;
signal \this_vga_signals.N_291_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb2\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_0\ : std_logic;
signal \M_this_oam_ram_read_data_20\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_20\ : std_logic;
signal \this_ppu.oam_cache.mem_13\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal \N_852_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \M_this_oam_ram_write_data_3\ : std_logic;
signal \M_this_data_tmp_qZ0Z_3\ : std_logic;
signal \M_this_oam_ram_write_data_4\ : std_logic;
signal \M_this_data_tmp_qZ0Z_4\ : std_logic;
signal \M_this_data_tmp_qZ0Z_5\ : std_logic;
signal \M_this_oam_ram_write_data_29\ : std_logic;
signal \M_this_oam_ram_write_data_21\ : std_logic;
signal \M_this_oam_ram_write_data_1\ : std_logic;
signal \M_this_oam_ram_write_data_25\ : std_logic;
signal \M_this_data_tmp_qZ0Z_21\ : std_logic;
signal \M_this_data_tmp_qZ0Z_23\ : std_logic;
signal \M_this_data_tmp_qZ0Z_0\ : std_logic;
signal \this_vga_ramdac.N_3856_reto\ : std_logic;
signal \this_vga_ramdac.i2_mux_cascade_\ : std_logic;
signal \this_vga_ramdac.N_3858_reto\ : std_logic;
signal \this_vga_ramdac.N_24_mux\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \this_vga_ramdac.m6_cascade_\ : std_logic;
signal \this_vga_ramdac.N_3857_reto\ : std_logic;
signal \this_ppu.oam_cache.mem_9\ : std_logic;
signal \this_vga_signals.M_pcounter_q_ret_RNIB85CZ0Z3_cascade_\ : std_logic;
signal \this_vga_signals.N_3_0_cascade_\ : std_logic;
signal \this_vga_ramdac.m16\ : std_logic;
signal \M_pcounter_q_ret_1_RNIOILK7_cascade_\ : std_logic;
signal \this_vga_ramdac.N_3859_reto\ : std_logic;
signal \this_vga_signals.N_2_0\ : std_logic;
signal \this_vga_signals.N_2_0_cascade_\ : std_logic;
signal \this_vga_ramdac.m19\ : std_logic;
signal \this_vga_ramdac.N_3860_reto\ : std_logic;
signal \this_ppu.oam_cache.mem_14\ : std_logic;
signal \this_ppu.m35_i_0_a3_0_cascade_\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_9\ : std_logic;
signal \this_ppu.oam_cache.mem_11\ : std_logic;
signal \this_ppu.oam_cache.mem_1\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_14\ : std_logic;
signal \this_ppu.N_1196_1\ : std_logic;
signal \this_ppu.M_oam_curr_qZ0Z_6\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_13\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNIRSG13Z0Z_9\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNIRSG13Z0Z_9_cascade_\ : std_logic;
signal \this_vga_signals.N_1307_1\ : std_logic;
signal \this_ppu.oam_cache.mem_8\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_11\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc1_0\ : std_logic;
signal \this_pixel_clk_M_counter_q_0\ : std_logic;
signal \this_pixel_clk_M_counter_q_i_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_2\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_3\ : std_logic;
signal \this_vga_signals.M_hcounter_q_RNII1437Z0Z_3\ : std_logic;
signal \M_this_oam_ram_read_data_30\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_30\ : std_logic;
signal \this_ppu.oam_cache.mem_3\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_1\ : std_logic;
signal \read_data_RNI5QFJ1_1\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_16\ : std_logic;
signal \M_this_ppu_spr_addr_3\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_2\ : std_logic;
signal \read_data_RNI6RFJ1_2\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_3\ : std_logic;
signal \read_data_RNI7SFJ1_3\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_4\ : std_logic;
signal \read_data_RNI9TFJ1_4\ : std_logic;
signal \this_vga_signals.M_pcounter_q_0Z0Z_1\ : std_logic;
signal \M_this_data_tmp_qZ0Z_11\ : std_logic;
signal \M_this_oam_ram_write_data_11\ : std_logic;
signal \M_this_oam_ram_write_data_12\ : std_logic;
signal \M_this_oam_ram_write_data_13\ : std_logic;
signal \M_this_oam_ram_write_data_14\ : std_logic;
signal \M_this_data_tmp_qZ0Z_12\ : std_logic;
signal \M_this_data_tmp_qZ0Z_14\ : std_logic;
signal \M_this_data_tmp_qZ0Z_1\ : std_logic;
signal \M_this_oam_ram_write_data_22\ : std_logic;
signal \M_this_data_tmp_qZ0Z_22\ : std_logic;
signal \M_this_map_ram_read_data_1\ : std_logic;
signal \N_724_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \this_vga_signals.N_1417\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_0\ : std_logic;
signal \this_vga_ramdac.i2_mux_0\ : std_logic;
signal \M_pcounter_q_ret_1_RNIOILK7\ : std_logic;
signal \this_vga_ramdac.N_3861_reto\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_ac0_11\ : std_logic;
signal \M_this_ppu_spr_addr_0\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_8\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_8\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_9\ : std_logic;
signal \M_this_ppu_spr_addr_1\ : std_logic;
signal \this_ppu.offset_x_cry_0\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_10\ : std_logic;
signal \M_this_ppu_spr_addr_2\ : std_logic;
signal \this_ppu.offset_x_cry_1\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_11\ : std_logic;
signal \this_ppu.m68_0_o2_0\ : std_logic;
signal \this_ppu.offset_x_cry_2\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_12\ : std_logic;
signal \this_ppu.offset_x_4\ : std_logic;
signal \this_ppu.offset_x_cry_3\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_13\ : std_logic;
signal \this_ppu.offset_x_5\ : std_logic;
signal \this_ppu.offset_x_cry_4\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_14\ : std_logic;
signal \M_this_ppu_map_addr_3\ : std_logic;
signal \this_ppu.offset_x_6\ : std_logic;
signal \this_ppu.offset_x_cry_5\ : std_logic;
signal \GNDG0\ : std_logic;
signal \this_ppu.offset_x_cry_6\ : std_logic;
signal \this_ppu.offset_x_cry_6_THRU_CRY_0_THRU_CO\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_15\ : std_logic;
signal \M_this_ppu_map_addr_4\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \this_ppu.offset_x_7\ : std_logic;
signal \this_ppu.m13_0_i_1\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \this_ppu.offset_y\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO\ : std_logic;
signal \this_ppu.M_screen_y_q_esr_RNI453Q6Z0Z_1\ : std_logic;
signal \this_ppu.M_surface_y_qZ0Z_1\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_0\ : std_logic;
signal \this_ppu.M_surface_y_qZ0Z_2\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_1\ : std_logic;
signal \M_this_ppu_map_addr_5\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_2\ : std_logic;
signal \this_ppu.M_screen_y_q_RNI8FJF7Z0Z_4\ : std_logic;
signal \M_this_ppu_map_addr_6\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_3\ : std_logic;
signal \M_this_ppu_map_addr_7\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_4\ : std_logic;
signal \M_this_ppu_map_addr_8\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_5\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_6\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \M_this_ppu_map_addr_9\ : std_logic;
signal \this_ppu.M_screen_y_q_esr_RNI563Q6Z0Z_2\ : std_logic;
signal \M_this_oam_ram_read_data_23\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_23\ : std_logic;
signal \M_this_oam_ram_read_data_1\ : std_logic;
signal \this_ppu.oam_cache.N_581_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_13\ : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal \M_this_data_count_q_cry_0\ : std_logic;
signal \M_this_data_count_q_cry_1\ : std_logic;
signal \M_this_data_count_q_cry_2\ : std_logic;
signal \M_this_data_count_q_cry_3\ : std_logic;
signal \M_this_data_count_q_cry_4\ : std_logic;
signal \M_this_data_count_q_cry_5\ : std_logic;
signal \M_this_data_count_q_cry_6\ : std_logic;
signal \M_this_data_count_q_cry_7\ : std_logic;
signal \bfn_14_25_0_\ : std_logic;
signal \M_this_data_count_q_cry_8\ : std_logic;
signal \M_this_data_count_q_cry_9\ : std_logic;
signal \M_this_data_count_q_cry_10\ : std_logic;
signal \M_this_data_count_q_cry_11\ : std_logic;
signal \M_this_data_count_q_cry_12\ : std_logic;
signal \M_this_oam_address_qZ0Z_7\ : std_logic;
signal \IO_port_data_write_i_m2_i_m2_0\ : std_logic;
signal \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\ : std_logic;
signal \this_ppu.M_state_qZ0Z_8\ : std_logic;
signal \this_ppu.N_762_0\ : std_logic;
signal \this_ppu.N_91_0\ : std_logic;
signal \this_ppu.N_91_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c3\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c3_cascade_\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c6\ : std_logic;
signal \this_ppu.N_1202\ : std_logic;
signal \this_ppu.M_state_qZ0Z_1\ : std_logic;
signal \M_this_status_flags_qZ0Z_0\ : std_logic;
signal \this_ppu.N_1201\ : std_logic;
signal \this_ppu.M_state_qZ0Z_4\ : std_logic;
signal \this_ppu.M_state_q_srsts_1_8\ : std_logic;
signal \this_ppu.N_1145\ : std_logic;
signal \this_ppu.M_screen_y_qZ0Z_7\ : std_logic;
signal \this_ppu.M_screen_y_qZ0Z_1\ : std_logic;
signal \this_ppu.un3_M_screen_y_d_0_c2\ : std_logic;
signal \this_ppu.un3_M_screen_y_d_0_c2_cascade_\ : std_logic;
signal \this_ppu.un3_M_screen_y_d_0_c4_cascade_\ : std_logic;
signal \this_ppu.un3_M_screen_y_d_0_c6\ : std_logic;
signal \N_861_0_cascade_\ : std_logic;
signal \this_ppu.M_screen_y_qZ0Z_2\ : std_logic;
signal \this_ppu.un3_M_screen_y_d_a_2\ : std_logic;
signal \M_this_ppu_vram_addr_7\ : std_logic;
signal \this_ppu.M_screen_y_q_RNIQ9FQ6Z0Z_0\ : std_logic;
signal \this_ppu.un1_M_screen_x_q_c4_cascade_\ : std_logic;
signal \this_ppu.un1_M_screen_x_q_c4\ : std_logic;
signal \M_this_ppu_vram_addr_4\ : std_logic;
signal \this_ppu.un1_M_screen_x_q_c5_cascade_\ : std_logic;
signal \M_this_ppu_vram_addr_5\ : std_logic;
signal \M_this_ppu_vram_addr_6\ : std_logic;
signal \M_this_ppu_vram_addr_2\ : std_logic;
signal \M_this_scroll_qZ0Z_0\ : std_logic;
signal \M_this_scroll_qZ0Z_1\ : std_logic;
signal \M_this_scroll_qZ0Z_2\ : std_logic;
signal \M_this_scroll_qZ0Z_4\ : std_logic;
signal \M_this_scroll_qZ0Z_7\ : std_logic;
signal this_vga_signals_vsync_1_i : std_logic;
signal \M_this_data_count_qZ0Z_0\ : std_logic;
signal \M_this_data_count_q_cry_0_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_1\ : std_logic;
signal \M_this_data_count_q_cry_1_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_2\ : std_logic;
signal \M_this_data_count_q_cry_2_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_3\ : std_logic;
signal \M_this_data_count_q_cry_3_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_4_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_5_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_10_THRU_CO\ : std_logic;
signal \M_this_data_count_q_s_10\ : std_logic;
signal \M_this_data_count_q_cry_11_THRU_CO\ : std_logic;
signal \M_this_data_count_q_s_13\ : std_logic;
signal \M_this_data_count_qZ0Z_12\ : std_logic;
signal \M_this_data_count_qZ0Z_11\ : std_logic;
signal \M_this_data_count_qZ0Z_13\ : std_logic;
signal \M_this_data_count_qZ0Z_10\ : std_logic;
signal \M_this_data_count_q_s_8\ : std_logic;
signal \M_this_data_count_qZ0Z_8\ : std_logic;
signal \M_this_data_count_qZ0Z_5\ : std_logic;
signal \M_this_data_count_qZ0Z_4\ : std_logic;
signal \un1_M_this_oam_address_q_c6\ : std_logic;
signal \this_vga_signals.g0_1\ : std_logic;
signal \this_vga_signals.N_3_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_2_1\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_CO\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_lcounter_q_e_1_0_cascade_\ : std_logic;
signal \N_26\ : std_logic;
signal \this_ppu.N_1198\ : std_logic;
signal \this_ppu.N_1198_cascade_\ : std_logic;
signal \M_this_ppu_map_addr_1\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c2_cascade_\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c5_cascade_\ : std_logic;
signal \M_this_ppu_map_addr_2\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c2\ : std_logic;
signal \this_ppu.offset_x\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c1\ : std_logic;
signal \M_this_ppu_map_addr_0\ : std_logic;
signal \this_ppu.M_surface_x_qZ0Z_2\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c1_cascade_\ : std_logic;
signal \this_ppu.M_surface_x_qZ0Z_1\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c4\ : std_logic;
signal \this_ppu.M_state_qZ0Z_2\ : std_logic;
signal \this_ppu.M_state_qZ0Z_10\ : std_logic;
signal \M_this_ppu_vram_addr_3\ : std_logic;
signal \this_ppu.N_798_0_cascade_\ : std_logic;
signal \M_this_ppu_vram_data_0\ : std_logic;
signal \this_ppu.N_1182_1\ : std_logic;
signal \this_ppu.M_state_qZ0Z_5\ : std_logic;
signal \this_vga_signals.g0_2\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \this_ppu.M_state_qZ0Z_6\ : std_logic;
signal \this_ppu.N_82_0\ : std_logic;
signal \this_ppu.N_1659_0\ : std_logic;
signal \this_ppu.M_screen_y_qZ0Z_3\ : std_logic;
signal \M_this_scroll_qZ0Z_3\ : std_logic;
signal \this_ppu.M_screen_y_q_esr_RNIF77F7Z0Z_3\ : std_logic;
signal \this_ppu.M_state_qZ0Z_9\ : std_logic;
signal \this_ppu.M_state_qZ0Z_7\ : std_logic;
signal \this_ppu.N_61_0\ : std_logic;
signal \M_this_ppu_vram_addr_1\ : std_logic;
signal \this_ppu.N_61_0_cascade_\ : std_logic;
signal \M_this_ppu_vram_addr_0\ : std_logic;
signal \this_ppu.un1_M_screen_x_q_c2\ : std_logic;
signal \this_ppu.M_state_d30_i_i_o2_3\ : std_logic;
signal \this_ppu.N_79_0\ : std_logic;
signal \this_ppu.N_79_0_cascade_\ : std_logic;
signal \this_ppu.M_pixel_cnt_q_600_1\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_d_1_sqmuxa_0_i_0_0\ : std_logic;
signal \this_ppu.N_999_0\ : std_logic;
signal \this_ppu.N_838_0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_0\ : std_logic;
signal \this_ppu.N_1042_0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_11\ : std_logic;
signal \this_ppu.M_state_qZ0Z_3\ : std_logic;
signal \this_ppu.N_1042_0_cascade_\ : std_logic;
signal \this_ppu.un30_0_a2_i_0\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ0Z_0\ : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ0Z_3\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ0Z_7\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_6_s1\ : std_logic;
signal \this_ppu.N_1205\ : std_logic;
signal \this_ppu.M_state_d30_i_i_o2_4\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ0Z_1\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ0Z_2\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ0Z_5\ : std_logic;
signal \this_ppu.N_1301_cascade_\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ0Z_6\ : std_logic;
signal \this_ppu.N_1730_0\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1_THRU_CO\ : std_logic;
signal \this_ppu.N_677_0\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ0Z_4\ : std_logic;
signal \M_this_data_count_q_cry_6_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_8_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_9\ : std_logic;
signal \N_231\ : std_logic;
signal \M_this_data_tmp_qZ0Z_2\ : std_logic;
signal \M_this_oam_ram_write_data_2\ : std_logic;
signal \M_this_data_count_qZ0Z_7\ : std_logic;
signal \M_this_data_count_qZ0Z_6\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_16\ : std_logic;
signal \N_1709_0\ : std_logic;
signal \N_1693_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNI01JU6Z0Z_9\ : std_logic;
signal \this_ppu.N_1269_cascade_\ : std_logic;
signal \this_ppu.N_1006_0\ : std_logic;
signal \this_vga_signals.N_1264_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_4_1_0_x0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_4_1_0_x1\ : std_logic;
signal \M_this_scroll_qZ0Z_10\ : std_logic;
signal \M_this_scroll_qZ0Z_11\ : std_logic;
signal \M_this_scroll_qZ0Z_12\ : std_logic;
signal \M_this_scroll_qZ0Z_13\ : std_logic;
signal \M_this_scroll_qZ0Z_14\ : std_logic;
signal \M_this_scroll_qZ0Z_15\ : std_logic;
signal \M_this_scroll_qZ0Z_8\ : std_logic;
signal \M_this_scroll_qZ0Z_9\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_2_cascade_\ : std_logic;
signal \this_vga_signals.N_4_0\ : std_logic;
signal \this_vga_signals.if_m1_0_x2_1\ : std_logic;
signal \this_vga_signals.r_N_2_i_0\ : std_logic;
signal \this_vga_signals.N_836_0\ : std_logic;
signal \this_vga_signals.N_1043_cascade_\ : std_logic;
signal \this_vga_signals_M_lcounter_q_0\ : std_logic;
signal \N_792_0\ : std_logic;
signal \this_vga_signals_M_lcounter_q_1\ : std_logic;
signal \this_ppu.M_last_q_0\ : std_logic;
signal \N_771_0\ : std_logic;
signal \N_771_0_cascade_\ : std_logic;
signal \this_ppu.N_774_0\ : std_logic;
signal \this_vga_signals.g1_0_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_6_0_0_0\ : std_logic;
signal \this_vga_signals.g1_0_0\ : std_logic;
signal \this_vga_signals.N_27_0_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_1_0_cascade_\ : std_logic;
signal \M_this_reset_cond_out_0\ : std_logic;
signal \N_782_0\ : std_logic;
signal \N_1725_0\ : std_logic;
signal \N_1717_0\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_12\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_3\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_16\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_16\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_a2_10Z0Z_16\ : std_logic;
signal \N_778_0_cascade_\ : std_logic;
signal \N_1701_0\ : std_logic;
signal \un1_M_this_oam_address_q_c5\ : std_logic;
signal \M_this_oam_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_oam_address_q_c5_cascade_\ : std_logic;
signal \M_this_oam_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_oam_address_q_c2\ : std_logic;
signal \M_this_oam_address_qZ0Z_2\ : std_logic;
signal \M_this_oam_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_oam_address_q_c3\ : std_logic;
signal \M_this_oam_address_qZ0Z_4\ : std_logic;
signal \M_this_oam_address_qZ0Z_1\ : std_logic;
signal \M_this_oam_address_qZ0Z_0\ : std_logic;
signal \N_778_0\ : std_logic;
signal \M_this_oam_ram_write_data_0_sqmuxa\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb2_i\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_2_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0\ : std_logic;
signal \this_ppu.N_1115\ : std_logic;
signal \this_vga_signals.g0_33_N_3L4\ : std_logic;
signal \this_vga_signals.g0_33_N_4L6\ : std_logic;
signal \this_vga_signals.g0_33_N_5L8\ : std_logic;
signal \this_vga_signals.M_hcounter_d7_0_i_0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \bfn_18_21_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_1\ : std_logic;
signal \G_535\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7\ : std_logic;
signal \bfn_18_22_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8\ : std_logic;
signal \this_vga_signals.g0_0_0\ : std_logic;
signal \this_vga_signals.IO_port_data_write_0_a2_i_o2_2Z0Z_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.vsync_1_0_a3_0_a3_5\ : std_logic;
signal \M_this_state_qZ0Z_12\ : std_logic;
signal \this_ppu.N_430_1_0_cascade_\ : std_logic;
signal \M_this_state_q_fastZ0Z_13\ : std_logic;
signal \this_vga_signals.N_38_i_0_a2_3Z0Z_0_cascade_\ : std_logic;
signal \this_vga_signals.N_38_i_0_a2_3_xZ0Z1_cascade_\ : std_logic;
signal \this_vga_signals.N_38_i_0_a2_3_cascade_\ : std_logic;
signal \this_vga_signals.N_38_i_0_a2_0_3\ : std_logic;
signal port_enb_c : std_logic;
signal \this_start_data_delay_M_last_q\ : std_logic;
signal \M_this_delay_clk_out_0\ : std_logic;
signal \N_765_0_cascade_\ : std_logic;
signal \this_ppu.N_229_1_0\ : std_logic;
signal \this_ppu.N_229_1_0_cascade_\ : std_logic;
signal \N_229\ : std_logic;
signal \N_1423\ : std_logic;
signal \this_vga_signals.SUM_2_i_i_1_0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_x1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_0_0_ns_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_0_1_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_0_1_1\ : std_logic;
signal \this_vga_signals.if_m5_s_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m5_d\ : std_logic;
signal \this_vga_signals.if_m5_d_cascade_\ : std_logic;
signal \this_vga_signals.N_2840_0_0\ : std_logic;
signal \this_vga_signals.N_27_0_0\ : std_logic;
signal \this_vga_signals.vaddress_7_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3\ : std_logic;
signal \this_vga_signals.g1_2_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m6_i_x2_3\ : std_logic;
signal \this_vga_signals.g1_3\ : std_logic;
signal \this_vga_signals_CO0_0_i_i\ : std_logic;
signal \this_vga_signals_CO0_0_i_i_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_8\ : std_logic;
signal \this_vga_signals.g1\ : std_logic;
signal \this_vga_signals.N_39_0\ : std_logic;
signal \this_vga_signals.vaddress_7\ : std_logic;
signal \this_vga_signals.N_38_i_0_a2_0_4Z0Z_1\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_17_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_17\ : std_logic;
signal \this_vga_signals.vsync_1_0_a3_0_a3_0\ : std_logic;
signal \M_this_state_qZ0Z_18\ : std_logic;
signal \this_ppu_M_this_map_address_d_4_sqmuxa_0_a3_i_o3_i_a3_0\ : std_logic;
signal \this_ppu.N_1322_cascade_\ : std_logic;
signal \M_this_spr_ram_write_data_0\ : std_logic;
signal \this_vga_signals.N_1247\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0_cascade_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_9\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_0_1_1_1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.M_vcounter_q_5_repZ0Z1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c2_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_4\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_4_3\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_x1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1\ : std_logic;
signal \this_vga_signals.N_27_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_x0\ : std_logic;
signal \this_vga_signals.if_N_7_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_d_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_1_3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_1_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_d\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.N_3_1_0_1\ : std_logic;
signal \this_vga_signals.g0_2_1\ : std_logic;
signal \this_vga_signals.g0_5\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0\ : std_logic;
signal \this_vga_signals.g0_1_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c2_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_0_3_1\ : std_logic;
signal \this_vga_signals.g0_0_3\ : std_logic;
signal \this_vga_signals.g1_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_0_1\ : std_logic;
signal \this_vga_signals.g0_2_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.vaddress_9\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_0_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_i\ : std_logic;
signal \this_vga_signals.g0_0_x2\ : std_logic;
signal \this_vga_signals.if_m5_i_0_0_0\ : std_logic;
signal \this_ppu.N_1002_0\ : std_logic;
signal \this_ppu.N_235_2_0\ : std_logic;
signal \this_ppu.N_235_2_0_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_7\ : std_logic;
signal \this_ppu.N_1162\ : std_logic;
signal \M_this_state_qZ0Z_9\ : std_logic;
signal \M_this_state_qZ0Z_11\ : std_logic;
signal \this_ppu.N_1301\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_i_0_0Z0Z_15\ : std_logic;
signal \M_this_state_qZ0Z_15\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_7\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_11\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_8\ : std_logic;
signal \this_ppu.N_807_0_cascade_\ : std_logic;
signal \this_ppu.N_1341\ : std_logic;
signal \M_this_spr_ram_write_data_2\ : std_logic;
signal \this_ppu.oam_cache.mem_5\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_1_3\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_0_3_cascade_\ : std_logic;
signal \this_vga_signals.N_7\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_2_3\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_3_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_2_0_3\ : std_logic;
signal \this_ppu.m18_i_o2_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_0_3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0\ : std_logic;
signal \N_814_0_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_2_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_2_2\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_0_2_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_x1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_x0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3\ : std_logic;
signal \this_vga_signals.g1_0\ : std_logic;
signal \this_vga_signals.g0_0_1\ : std_logic;
signal \this_vga_signals.g0_3_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c2_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_9_repZ0Z1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_4_1_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_8_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_7_repZ0Z1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_3_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.SUM_2_i_i_1_0_3\ : std_logic;
signal \this_vga_signals.N_5_0_0\ : std_logic;
signal \this_vga_signals.g1_0_1\ : std_logic;
signal \this_vga_signals.N_39_0_0\ : std_logic;
signal \this_vga_signals.g1_3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.N_4_1\ : std_logic;
signal \this_vga_signals.g3_cascade_\ : std_logic;
signal \this_vga_signals.N_5_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_0_0_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_0_0_1\ : std_logic;
signal \this_vga_signals.N_1264\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\ : std_logic;
signal \this_vga_signals_M_vcounter_q_8\ : std_logic;
signal \N_1001_0\ : std_logic;
signal \N_814_0\ : std_logic;
signal \N_1001_0_cascade_\ : std_logic;
signal \this_vga_signals_M_vcounter_q_9\ : std_logic;
signal \this_vga_signals.g4\ : std_logic;
signal \this_ppu.N_1278_cascade_\ : std_logic;
signal \this_ppu.N_767_0\ : std_logic;
signal \this_ppu.N_1425\ : std_logic;
signal \this_ppu.N_1149_cascade_\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_0_a3_1_2_1Z0Z_0\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_0_0_tz_0_0\ : std_logic;
signal \M_this_state_qZ0Z_8\ : std_logic;
signal \N_815_0\ : std_logic;
signal led_c_7 : std_logic;
signal \this_ppu.N_807_0\ : std_logic;
signal \M_this_state_qZ0Z_16\ : std_logic;
signal \N_1415\ : std_logic;
signal \N_1415_cascade_\ : std_logic;
signal \this_ppu.N_1278\ : std_logic;
signal \this_ppu.N_1166\ : std_logic;
signal \this_ppu.N_1263_cascade_\ : std_logic;
signal \this_ppu.N_1176_1\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_3\ : std_logic;
signal \this_ppu.N_893\ : std_logic;
signal \this_ppu.N_969\ : std_logic;
signal \un1_M_this_state_q_11_0_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_this_state_q_11_0_0Z0Z_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_this_state_q_11_0_0Z0Z_1\ : std_logic;
signal \this_ppu.N_430_1_0\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_2\ : std_logic;
signal \this_ppu.N_1158_cascade_\ : std_logic;
signal \this_ppu.N_1263\ : std_logic;
signal port_address_in_4 : std_logic;
signal port_address_in_0 : std_logic;
signal port_rw_in : std_logic;
signal \N_1422\ : std_logic;
signal \M_this_spr_address_qZ0Z_0\ : std_logic;
signal \bfn_22_14_0_\ : std_logic;
signal \M_this_spr_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_spr_address_q_cry_0\ : std_logic;
signal \M_this_spr_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_spr_address_q_cry_1\ : std_logic;
signal \M_this_spr_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_spr_address_q_cry_2\ : std_logic;
signal \M_this_spr_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_spr_address_q_cry_3\ : std_logic;
signal \M_this_spr_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_spr_address_q_cry_4\ : std_logic;
signal \M_this_spr_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_spr_address_q_cry_5\ : std_logic;
signal \M_this_spr_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_spr_address_q_cry_6\ : std_logic;
signal \un1_M_this_spr_address_q_cry_7\ : std_logic;
signal \M_this_spr_address_qZ0Z_8\ : std_logic;
signal \bfn_22_15_0_\ : std_logic;
signal \M_this_spr_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_spr_address_q_cry_8\ : std_logic;
signal \M_this_spr_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_spr_address_q_cry_9\ : std_logic;
signal \un1_M_this_spr_address_q_cry_10\ : std_logic;
signal \un1_M_this_spr_address_q_cry_11\ : std_logic;
signal \N_1005_0\ : std_logic;
signal \un1_M_this_spr_address_q_cry_12\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_5\ : std_logic;
signal \this_ppu.oam_cache.mem_6\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_6\ : std_logic;
signal \this_spr_ram.mem_out_bus4_2\ : std_logic;
signal \this_spr_ram.mem_out_bus0_2\ : std_logic;
signal \this_spr_ram.mem_mem_0_1_RNIM6VFZ0_cascade_\ : std_logic;
signal \this_spr_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\ : std_logic;
signal \M_this_spr_ram_read_data_2_cascade_\ : std_logic;
signal \M_this_ppu_vram_data_2\ : std_logic;
signal \this_spr_ram.mem_out_bus5_0\ : std_logic;
signal \this_spr_ram.mem_out_bus1_0\ : std_logic;
signal \this_spr_ram.mem_out_bus4_1\ : std_logic;
signal \this_spr_ram.mem_out_bus0_1\ : std_logic;
signal \this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0_cascade_\ : std_logic;
signal \this_spr_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\ : std_logic;
signal \M_this_spr_ram_read_data_2\ : std_logic;
signal \M_this_spr_ram_read_data_1_cascade_\ : std_logic;
signal \this_ppu.N_1000_0\ : std_logic;
signal \M_this_spr_ram_read_data_1\ : std_logic;
signal \M_this_ppu_vram_data_1\ : std_logic;
signal \this_spr_ram.mem_mem_1_0_RNIMA1GZ0\ : std_logic;
signal \M_this_spr_ram_read_data_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\ : std_logic;
signal \this_vga_signals.N_1307_0_g\ : std_logic;
signal \this_vga_signals.N_1637_g\ : std_logic;
signal \this_vga_signals.N_5_i_0\ : std_logic;
signal \this_vga_signals.N_5_i_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_0_1\ : std_logic;
signal \this_vga_signals.g0_21_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_ns\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_3\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_1_1\ : std_logic;
signal \this_vga_signals.vaddress_6\ : std_logic;
signal \this_vga_signals.vaddress_5\ : std_logic;
signal \this_vga_signals.g2_1_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_4\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_2_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1\ : std_logic;
signal \this_vga_signals.if_N_7_0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_d_0_0\ : std_logic;
signal \this_vga_signals_M_vcounter_q_4\ : std_logic;
signal \this_vga_signals_M_vcounter_q_7\ : std_logic;
signal \this_vga_signals_M_vcounter_q_5\ : std_logic;
signal \this_vga_signals_M_vcounter_q_6\ : std_logic;
signal \this_vga_signals.vaddress_0_0_7\ : std_logic;
signal \M_this_scroll_qZ0Z_6\ : std_logic;
signal \this_ppu.M_screen_y_q_esr_RNILD7F7Z0Z_6\ : std_logic;
signal \M_this_spr_ram_write_data_3\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_0_a2_1_xZ0Z_0\ : std_logic;
signal \this_ppu.N_798_0\ : std_logic;
signal \this_ppu.N_1426\ : std_logic;
signal \M_this_ppu_vram_data_3\ : std_logic;
signal \this_ppu.N_1257\ : std_logic;
signal \this_ppu.N_1322\ : std_logic;
signal \M_this_spr_ram_write_data_1\ : std_logic;
signal led_c_1 : std_logic;
signal \N_1416_cascade_\ : std_logic;
signal \N_1151_3\ : std_logic;
signal \this_ppu.N_787_0\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_0_a2_1_sxZ0Z_0\ : std_logic;
signal \M_this_state_qZ0Z_14\ : std_logic;
signal \M_this_state_qZ0Z_13\ : std_logic;
signal \M_this_spr_ram_write_en_0_i_1_0\ : std_logic;
signal \M_this_state_qZ0Z_3\ : std_logic;
signal port_address_in_2 : std_logic;
signal port_address_in_1 : std_logic;
signal \M_this_substate_qZ0\ : std_logic;
signal \this_ppu_M_this_substate_d_0_sqmuxa_3_0_a3_0_a3_1\ : std_logic;
signal \M_this_map_address_qc_3_0_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_10\ : std_logic;
signal \N_169_0\ : std_logic;
signal \N_1048_i\ : std_logic;
signal \this_spr_ram.mem_out_bus5_1\ : std_logic;
signal \this_spr_ram.mem_out_bus1_1\ : std_logic;
signal \this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0\ : std_logic;
signal \this_spr_ram.mem_out_bus5_2\ : std_logic;
signal \this_spr_ram.mem_out_bus1_2\ : std_logic;
signal \this_spr_ram.mem_mem_1_1_RNIOA1GZ0\ : std_logic;
signal \this_spr_ram.mem_out_bus6_0\ : std_logic;
signal \this_spr_ram.mem_out_bus2_0\ : std_logic;
signal \this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_\ : std_logic;
signal \this_spr_ram.mem_DOUT_7_i_m2_ns_1_0\ : std_logic;
signal \this_spr_ram.mem_WE_0\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_7\ : std_logic;
signal \this_spr_ram.mem_out_bus6_2\ : std_logic;
signal \this_spr_ram.mem_out_bus2_2\ : std_logic;
signal \this_spr_ram.mem_mem_2_1_RNIQE3GZ0\ : std_logic;
signal \this_spr_ram.mem_out_bus4_3\ : std_logic;
signal \this_spr_ram.mem_out_bus0_3\ : std_logic;
signal \this_ppu.N_753_0\ : std_logic;
signal \this_ppu.M_screen_y_qZ0Z_6\ : std_logic;
signal \this_ppu.M_screen_y_qZ0Z_4\ : std_logic;
signal \this_ppu.un3_M_screen_y_d_0_c4\ : std_logic;
signal \N_861_0\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_0\ : std_logic;
signal \this_ppu.M_screen_y_qZ0Z_5\ : std_logic;
signal \M_this_scroll_qZ0Z_5\ : std_logic;
signal \this_ppu.M_screen_y_q_esr_RNIJB7F7Z0Z_5\ : std_logic;
signal \this_spr_ram.mem_radregZ0Z_12\ : std_logic;
signal \this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0\ : std_logic;
signal \this_spr_ram.mem_radregZ0Z_11\ : std_logic;
signal \this_spr_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\ : std_logic;
signal \M_this_spr_ram_read_data_3\ : std_logic;
signal \this_spr_ram.mem_out_bus5_3\ : std_logic;
signal \this_spr_ram.mem_out_bus1_3\ : std_logic;
signal \this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0\ : std_logic;
signal \this_spr_ram.mem_out_bus6_3\ : std_logic;
signal \this_spr_ram.mem_out_bus2_3\ : std_logic;
signal \this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0\ : std_logic;
signal \this_spr_ram.mem_out_bus7_0\ : std_logic;
signal \this_spr_ram.mem_out_bus3_0\ : std_logic;
signal \this_spr_ram.mem_mem_3_0_RNIQI5GZ0\ : std_logic;
signal \this_spr_ram.mem_out_bus7_1\ : std_logic;
signal \this_spr_ram.mem_out_bus3_1\ : std_logic;
signal \this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0\ : std_logic;
signal \this_spr_ram.mem_out_bus7_2\ : std_logic;
signal \this_spr_ram.mem_out_bus3_2\ : std_logic;
signal \this_spr_ram.mem_mem_3_1_RNISI5GZ0\ : std_logic;
signal \this_spr_ram.mem_out_bus7_3\ : std_logic;
signal \this_spr_ram.mem_out_bus3_3\ : std_logic;
signal \this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0\ : std_logic;
signal \M_this_ctrl_flags_qZ0Z_7\ : std_logic;
signal \M_this_state_qZ0Z_2\ : std_logic;
signal \N_38_i_0\ : std_logic;
signal \N_38_i_0_i\ : std_logic;
signal \this_ppu.N_856_0\ : std_logic;
signal \this_ppu_un1_M_this_state_q_7_i_0_0_0_cascade_\ : std_logic;
signal \N_816_0\ : std_logic;
signal \N_1416\ : std_logic;
signal \M_this_state_qZ0Z_5\ : std_logic;
signal led_c_6 : std_logic;
signal \M_this_state_qZ0Z_6\ : std_logic;
signal \this_ppu_un1_M_this_state_q_7_i_0_0_0\ : std_logic;
signal \un1_M_this_state_q_7_i_0_a3_0_0_cascade_\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0\ : std_logic;
signal \M_this_map_ram_read_data_0\ : std_logic;
signal \this_ppu.N_785_0\ : std_logic;
signal \read_data_RNI4PFJ1_0\ : std_logic;
signal \N_1058\ : std_logic;
signal \N_1062_cascade_\ : std_logic;
signal \M_this_map_address_qc_5_0\ : std_logic;
signal \N_1066\ : std_logic;
signal \M_this_map_address_qc_6_0_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_4\ : std_logic;
signal \N_794_0\ : std_logic;
signal \M_this_map_address_qc_4_0\ : std_logic;
signal \N_918_0\ : std_logic;
signal m5_i_a2_i_o3_i_a3 : std_logic;
signal \N_1048_i_0\ : std_logic;
signal \this_spr_ram.mem_WE_12\ : std_logic;
signal \this_spr_ram.mem_WE_8\ : std_logic;
signal \this_spr_ram.mem_WE_14\ : std_logic;
signal \this_spr_ram.mem_WE_10\ : std_logic;
signal \this_spr_ram.mem_out_bus4_0\ : std_logic;
signal \this_spr_ram.mem_out_bus0_0\ : std_logic;
signal \this_spr_ram.mem_mem_0_0_RNIK6VFZ0\ : std_logic;
signal \this_spr_ram.mem_out_bus2_1\ : std_logic;
signal \this_spr_ram.mem_radregZ0Z_13\ : std_logic;
signal \this_spr_ram.mem_out_bus6_1\ : std_logic;
signal \this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0\ : std_logic;
signal \M_this_map_ram_read_data_7\ : std_logic;
signal \IO_port_data_write_i_m2_i_m2_7\ : std_logic;
signal \this_spr_ram.mem_WE_6\ : std_logic;
signal \this_spr_ram.mem_WE_4\ : std_logic;
signal \M_this_spr_address_qZ0Z_12\ : std_logic;
signal \M_this_spr_address_qZ0Z_11\ : std_logic;
signal \M_this_spr_address_qZ0Z_13\ : std_logic;
signal \M_this_spr_ram_write_en_0_i_1_0_0\ : std_logic;
signal \this_spr_ram.mem_WE_2\ : std_logic;
signal \N_842_0\ : std_logic;
signal \M_this_status_flags_qZ0Z_7\ : std_logic;
signal \M_this_map_address_qc_3_1\ : std_logic;
signal \un1_M_this_map_address_q_cry_0_c_RNOZ0\ : std_logic;
signal \bfn_24_23_0_\ : std_logic;
signal \M_this_map_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_map_address_q_cry_0_THRU_CO\ : std_logic;
signal \un1_M_this_map_address_q_cry_0\ : std_logic;
signal \M_this_map_address_qZ0Z_2\ : std_logic;
signal \M_this_map_address_q_RNO_1Z0Z_2\ : std_logic;
signal \un1_M_this_map_address_q_cry_1\ : std_logic;
signal \M_this_map_address_qZ0Z_3\ : std_logic;
signal \M_this_map_address_q_RNO_1Z0Z_3\ : std_logic;
signal \un1_M_this_map_address_q_cry_2\ : std_logic;
signal \M_this_map_address_qZ0Z_4\ : std_logic;
signal \M_this_map_address_q_RNO_1Z0Z_4\ : std_logic;
signal \un1_M_this_map_address_q_cry_3\ : std_logic;
signal \un1_M_this_state_q_7_i_0_a3_0_0\ : std_logic;
signal \un1_M_this_map_address_q_cry_4\ : std_logic;
signal \un1_M_this_map_address_q_cry_5\ : std_logic;
signal \un1_M_this_map_address_q_cry_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_7\ : std_logic;
signal \bfn_24_24_0_\ : std_logic;
signal \un1_M_this_map_address_q_cry_8\ : std_logic;
signal \un1_M_this_map_address_q_cry_5_THRU_CO\ : std_logic;
signal port_data_in_1 : std_logic;
signal \M_this_map_address_qc_8_1_cascade_\ : std_logic;
signal \M_this_map_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_7_THRU_CO\ : std_logic;
signal \un1_M_this_map_address_q_axb_0\ : std_logic;
signal \M_this_map_address_qc_2_0\ : std_logic;
signal \N_1097\ : std_logic;
signal \M_this_map_address_qZ0Z_0\ : std_logic;
signal \N_921_0\ : std_logic;
signal \N_919_0\ : std_logic;
signal \N_923_0\ : std_logic;
signal \N_920_0\ : std_logic;
signal \N_922_0\ : std_logic;
signal \N_296_0\ : std_logic;
signal \N_924_0\ : std_logic;
signal port_data_in_5 : std_logic;
signal \M_this_ctrl_flags_qZ0Z_5\ : std_logic;
signal port_data_in_7 : std_logic;
signal \M_this_ctrl_flags_qZ0Z_6\ : std_logic;
signal port_data_in_6 : std_logic;
signal \N_247\ : std_logic;
signal \M_this_ext_address_qZ0Z_0\ : std_logic;
signal \bfn_26_21_0_\ : std_logic;
signal \un1_M_this_ext_address_q_cry_0\ : std_logic;
signal \M_this_ext_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_ext_address_q_cry_1_THRU_CO\ : std_logic;
signal \un1_M_this_ext_address_q_cry_1\ : std_logic;
signal \un1_M_this_ext_address_q_cry_2\ : std_logic;
signal \un1_M_this_ext_address_q_cry_3\ : std_logic;
signal \un1_M_this_ext_address_q_cry_4\ : std_logic;
signal \un1_M_this_ext_address_q_cry_5\ : std_logic;
signal \un1_M_this_ext_address_q_cry_6\ : std_logic;
signal \un1_M_this_ext_address_q_cry_7\ : std_logic;
signal \bfn_26_22_0_\ : std_logic;
signal \M_this_ext_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_ext_address_q_cry_8_c_RNIS45FZ0\ : std_logic;
signal \un1_M_this_ext_address_q_cry_8\ : std_logic;
signal \un1_M_this_ext_address_q_cry_9\ : std_logic;
signal \un1_M_this_ext_address_q_cry_10\ : std_logic;
signal \un1_M_this_ext_address_q_cry_11\ : std_logic;
signal \M_this_ext_address_qZ0Z_13\ : std_logic;
signal \un1_M_this_ext_address_q_cry_12_c_RNIIMQAZ0\ : std_logic;
signal \un1_M_this_ext_address_q_cry_12\ : std_logic;
signal \M_this_ext_address_qZ0Z_14\ : std_logic;
signal \un1_M_this_ext_address_q_cry_13_c_RNIKPRAZ0\ : std_logic;
signal \un1_M_this_ext_address_q_cry_13\ : std_logic;
signal \M_this_ext_address_qZ0Z_15\ : std_logic;
signal \un1_M_this_ext_address_q_cry_14\ : std_logic;
signal \un1_M_this_ext_address_q_cry_14_c_RNIMSSAZ0\ : std_logic;
signal \un1_M_this_ext_address_q_cry_9_c_RNI55NHZ0\ : std_logic;
signal \M_this_ext_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_ext_address_q_cry_6_THRU_CO\ : std_logic;
signal \M_this_ext_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_ext_address_q_cry_10_c_RNIEGOAZ0\ : std_logic;
signal \M_this_ext_address_qZ0Z_11\ : std_logic;
signal \un1_M_this_ext_address_q_cry_11_c_RNIGJPAZ0\ : std_logic;
signal \M_this_ext_address_qZ0Z_12\ : std_logic;
signal \M_this_state_qZ0Z_1\ : std_logic;
signal \M_this_ctrl_flags_qZ0Z_4\ : std_logic;
signal \M_this_map_address_qZ0Z_9\ : std_logic;
signal port_data_in_4 : std_logic;
signal \N_1081_cascade_\ : std_logic;
signal \M_this_map_address_qc_1_1\ : std_logic;
signal \M_this_map_address_qZ0Z_8\ : std_logic;
signal port_data_in_3 : std_logic;
signal \N_1078_cascade_\ : std_logic;
signal \M_this_map_address_qc_0_1\ : std_logic;
signal \M_this_map_ram_read_data_2\ : std_logic;
signal \N_726_0\ : std_logic;
signal \un1_M_this_ext_address_q_cry_7_c_RNIQ14FZ0\ : std_logic;
signal \M_this_ext_address_qZ0Z_8\ : std_logic;
signal \un1_M_this_ext_address_q_cry_0_THRU_CO\ : std_logic;
signal \M_this_ext_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_ext_address_q_cry_2_THRU_CO\ : std_logic;
signal \M_this_ext_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_ext_address_q_cry_3_THRU_CO\ : std_logic;
signal \M_this_ext_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_ext_address_q_cry_4_THRU_CO\ : std_logic;
signal \M_this_ext_address_qZ0Z_5\ : std_logic;
signal \N_773_0\ : std_logic;
signal \N_765_0\ : std_logic;
signal \un1_M_this_ext_address_q_cry_5_THRU_CO\ : std_logic;
signal \M_this_ext_address_qZ0Z_6\ : std_logic;
signal \M_this_reset_cond_out_g_0\ : std_logic;
signal \un1_M_this_map_address_q_cry_6_THRU_CO\ : std_logic;
signal \M_this_map_address_qZ0Z_7\ : std_logic;
signal \N_801_0\ : std_logic;
signal port_data_in_2 : std_logic;
signal \N_1075_cascade_\ : std_logic;
signal \M_this_map_address_qc_1_0\ : std_logic;
signal port_address_in_3 : std_logic;
signal \N_459_0\ : std_logic;
signal \N_1276\ : std_logic;
signal \N_1242\ : std_logic;
signal port_data_in_0 : std_logic;
signal \N_1068\ : std_logic;
signal \M_this_map_address_qc_7_1\ : std_logic;
signal \M_this_map_address_q_RNO_1Z0Z_5\ : std_logic;
signal \N_1258\ : std_logic;
signal \M_this_map_address_qZ0Z_5\ : std_logic;
signal clk_0_c_g : std_logic;
signal \N_620_g\ : std_logic;
signal \M_this_map_ram_read_data_6\ : std_logic;
signal \N_734_0\ : std_logic;
signal \M_this_map_ram_read_data_5\ : std_logic;
signal \N_996_0\ : std_logic;
signal port_address_in_6 : std_logic;
signal port_address_in_5 : std_logic;
signal port_address_in_7 : std_logic;
signal \M_this_substate_d_0_sqmuxa_3_0_o2_x\ : std_logic;
signal \M_this_map_ram_read_data_4\ : std_logic;
signal \N_730_0\ : std_logic;
signal \this_vga_signals.N_834_0\ : std_logic;
signal \M_this_map_ram_read_data_3\ : std_logic;
signal \N_728_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic_vector(1 downto 0);
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal led_wire : std_logic_vector(7 downto 0);
signal port_clk_wire : std_logic;
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_map_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    led <= led_wire;
    port_clk_wire <= port_clk;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \M_this_map_ram_read_data_3\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_2\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_1\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_0\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&\N__21724\&\N__21343\&\N__21388\&\N__21427\&\N__21475\&\N__21187\&\N__21259\&\N__22924\&\N__23008\&\N__23416\;
    \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&\N__40825\&\N__41560\&\N__42886\&\N__39646\&\N__42190\&\N__39244\&\N__39289\&\N__39331\&\N__39388\&\N__39574\;
    \this_map_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&\N__40171\&'0'&'0'&'0'&\N__40186\&'0'&'0'&'0'&\N__38494\&'0'&'0'&'0'&\N__36076\&'0';
    \M_this_map_ram_read_data_7\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_6\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_5\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_4\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&\N__21718\&\N__21337\&\N__21382\&\N__21420\&\N__21469\&\N__21181\&\N__21253\&\N__22918\&\N__23001\&\N__23410\;
    \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&\N__40819\&\N__41554\&\N__42880\&\N__39640\&\N__42184\&\N__39238\&\N__39283\&\N__39325\&\N__39382\&\N__39568\;
    \this_map_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&\N__40075\&'0'&'0'&'0'&\N__40180\&'0'&'0'&'0'&\N__40165\&'0'&'0'&'0'&\N__39520\&'0';
    \M_this_oam_ram_read_data_15\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(15);
    \M_this_oam_ram_read_data_14\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(14);
    \M_this_oam_ram_read_data_13\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_oam_ram_read_data_12\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(12);
    \M_this_oam_ram_read_data_11\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \M_this_oam_ram_read_data_10\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(10);
    \M_this_oam_ram_read_data_9\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_oam_ram_read_data_8\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(8);
    \M_this_oam_ram_read_data_7\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(7);
    \M_this_oam_ram_read_data_6\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(6);
    \M_this_oam_ram_read_data_5\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_oam_ram_read_data_4\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(4);
    \M_this_oam_ram_read_data_3\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_oam_ram_read_data_2\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_oam_ram_read_data_1\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_0\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__16678\&\N__15631\&\N__15757\&\N__15694\&\N__15451\&\N__16639\;
    \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__21814\&\N__26470\&\N__26521\&\N__26932\&\N__26998\&\N__26413\;
    \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ <= \N__17098\&\N__19276\&\N__19285\&\N__19294\&\N__19303\&\N__16318\&\N__16549\&\N__16519\&\N__17029\&\N__17050\&\N__16147\&\N__18010\&\N__18028\&\N__25327\&\N__18190\&\N__17230\;
    \M_this_oam_ram_read_data_31\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(15);
    \M_this_oam_ram_read_data_30\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(14);
    \M_this_oam_ram_read_data_29\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(13);
    \M_this_oam_ram_read_data_28\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(12);
    \M_this_oam_ram_read_data_27\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \M_this_oam_ram_read_data_26\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(10);
    \M_this_oam_ram_read_data_25\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(9);
    \M_this_oam_ram_read_data_24\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(8);
    \M_this_oam_ram_read_data_23\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(7);
    \M_this_oam_ram_read_data_22\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(6);
    \M_this_oam_ram_read_data_21\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_oam_ram_read_data_20\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(4);
    \M_this_oam_ram_read_data_19\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \M_this_oam_ram_read_data_18\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(2);
    \M_this_oam_ram_read_data_17\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_16\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__16672\&\N__15625\&\N__15751\&\N__15688\&\N__15445\&\N__16633\;
    \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__21808\&\N__26464\&\N__26515\&\N__26926\&\N__26992\&\N__26407\;
    \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ <= \N__16507\&\N__17113\&\N__17980\&\N__16528\&\N__17122\&\N__17131\&\N__18178\&\N__16489\&\N__15373\&\N__20221\&\N__17971\&\N__15367\&\N__15361\&\N__15205\&\N__15355\&\N__16498\;
    \this_ppu.oam_cache.mem_15\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(15);
    \this_ppu.oam_cache.mem_14\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(14);
    \this_ppu.oam_cache.mem_13\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(13);
    \this_ppu.oam_cache.mem_12\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(12);
    \this_ppu.oam_cache.mem_11\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_ppu.oam_cache.mem_10\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(10);
    \this_ppu.oam_cache.mem_9\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(9);
    \this_ppu.oam_cache.mem_8\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(8);
    \this_ppu.oam_cache.mem_7\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(7);
    \this_ppu.oam_cache.mem_6\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(6);
    \this_ppu.oam_cache.mem_5\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(5);
    \this_ppu.oam_cache.mem_4\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(4);
    \this_ppu.oam_cache.mem_3\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_ppu.oam_cache.mem_2\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(2);
    \this_ppu.oam_cache.mem_1\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(1);
    \this_ppu.oam_cache.mem_0\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_ppu.oam_cache.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__14788\&\N__14809\&\N__14824\&\N__14875\;
    \this_ppu.oam_cache.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__15535\&\N__22657\&\N__15805\&\N__16060\;
    \this_ppu.oam_cache.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_ppu.oam_cache.mem_mem_0_0_physical_WDATA_wire\ <= \N__14737\&\N__16450\&\N__13990\&\N__14614\&\N__17476\&\N__14668\&\N__14689\&\N__14707\&\N__14530\&\N__14725\&\N__16765\&\N__16732\&\N__14731\&\N__14602\&\N__21613\&\N__15301\;
    \this_ppu.oam_cache.mem_18\ <= \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\(2);
    \this_ppu.oam_cache.mem_17\ <= \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\(1);
    \this_ppu.oam_cache.mem_16\ <= \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\(0);
    \this_ppu.oam_cache.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__14782\&\N__14803\&\N__14818\&\N__14869\;
    \this_ppu.oam_cache.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__15529\&\N__22650\&\N__15799\&\N__16054\;
    \this_ppu.oam_cache.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_ppu.oam_cache.mem_mem_0_1_physical_WDATA_wire\ <= \N__16363\&\N__18964\&\N__16420\&\N__16282\&\N__16888\&\N__14578\&\N__14974\&\N__15946\&\N__21655\&\N__15031\&\N__15037\&\N__17566\&\N__16351\&\N__16159\&\N__16987\&\N__14662\;
    \this_spr_ram.mem_out_bus0_1\ <= \this_spr_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus0_0\ <= \this_spr_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_0_0_physical_RADDR_wire\ <= \N__19517\&\N__19715\&\N__19939\&\N__18921\&\N__38080\&\N__14283\&\N__14482\&\N__20129\&\N__20653\&\N__20878\&\N__21111\;
    \this_spr_ram.mem_mem_0_0_physical_WADDR_wire\ <= \N__33419\&\N__33607\&\N__33891\&\N__31338\&\N__31544\&\N__31713\&\N__31971\&\N__32172\&\N__32390\&\N__32601\&\N__32845\;
    \this_spr_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__35965\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28126\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus0_3\ <= \this_spr_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus0_2\ <= \this_spr_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_0_1_physical_RADDR_wire\ <= \N__19516\&\N__19714\&\N__19938\&\N__18922\&\N__38079\&\N__14284\&\N__14466\&\N__20128\&\N__20605\&\N__20874\&\N__21112\;
    \this_spr_ram.mem_mem_0_1_physical_WADDR_wire\ <= \N__33443\&\N__33673\&\N__33881\&\N__31337\&\N__31543\&\N__31712\&\N__31962\&\N__32171\&\N__32380\&\N__32602\&\N__32839\;
    \this_spr_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__34577\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__29428\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus1_1\ <= \this_spr_ram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus1_0\ <= \this_spr_ram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_1_0_physical_RADDR_wire\ <= \N__19501\&\N__19717\&\N__19929\&\N__18917\&\N__38105\&\N__14282\&\N__14409\&\N__20140\&\N__20665\&\N__20867\&\N__21132\;
    \this_spr_ram.mem_mem_1_0_physical_WADDR_wire\ <= \N__33386\&\N__33658\&\N__33860\&\N__31316\&\N__31526\&\N__31735\&\N__31945\&\N__32150\&\N__32365\&\N__32631\&\N__32823\;
    \this_spr_ram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__35960\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28122\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus1_3\ <= \this_spr_ram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus1_2\ <= \this_spr_ram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_1_1_physical_RADDR_wire\ <= \N__19500\&\N__19713\&\N__19928\&\N__18906\&\N__38104\&\N__14280\&\N__14494\&\N__20139\&\N__20661\&\N__20857\&\N__21103\;
    \this_spr_ram.mem_mem_1_1_physical_WADDR_wire\ <= \N__33423\&\N__33633\&\N__33830\&\N__31315\&\N__31525\&\N__31708\&\N__31921\&\N__32149\&\N__32342\&\N__32632\&\N__32796\;
    \this_spr_ram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__34576\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__29423\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus2_1\ <= \this_spr_ram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus2_0\ <= \this_spr_ram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_2_0_physical_RADDR_wire\ <= \N__19522\&\N__19709\&\N__19905\&\N__18905\&\N__38090\&\N__14269\&\N__14490\&\N__20132\&\N__20654\&\N__20845\&\N__21104\;
    \this_spr_ram.mem_mem_2_0_physical_WADDR_wire\ <= \N__33372\&\N__33597\&\N__33794\&\N__31282\&\N__31492\&\N__31707\&\N__31888\&\N__32116\&\N__32313\&\N__32579\&\N__32761\;
    \this_spr_ram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__35950\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28115\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus2_3\ <= \this_spr_ram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus2_2\ <= \this_spr_ram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_2_1_physical_RADDR_wire\ <= \N__19499\&\N__19685\&\N__19869\&\N__18904\&\N__38053\&\N__14268\&\N__14483\&\N__20118\&\N__20642\&\N__20833\&\N__21134\;
    \this_spr_ram.mem_mem_2_1_physical_WADDR_wire\ <= \N__33432\&\N__33616\&\N__33813\&\N__31241\&\N__31424\&\N__31648\&\N__31830\&\N__32055\&\N__32259\&\N__32537\&\N__32702\;
    \this_spr_ram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__34553\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__29411\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus3_1\ <= \this_spr_ram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus3_0\ <= \this_spr_ram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_3_0_physical_RADDR_wire\ <= \N__19518\&\N__19684\&\N__19937\&\N__18903\&\N__38069\&\N__14267\&\N__14470\&\N__20117\&\N__20620\&\N__20817\&\N__21133\;
    \this_spr_ram.mem_mem_3_0_physical_WADDR_wire\ <= \N__33403\&\N__33576\&\N__33773\&\N__31242\&\N__31475\&\N__31694\&\N__31869\&\N__32099\&\N__32296\&\N__32613\&\N__32742\;
    \this_spr_ram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__35936\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28105\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus3_3\ <= \this_spr_ram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus3_2\ <= \this_spr_ram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_3_1_physical_RADDR_wire\ <= \N__19498\&\N__19683\&\N__19924\&\N__18916\&\N__38040\&\N__14276\&\N__14446\&\N__20116\&\N__20609\&\N__20790\&\N__21126\;
    \this_spr_ram.mem_mem_3_1_physical_WADDR_wire\ <= \N__33433\&\N__33649\&\N__33814\&\N__31258\&\N__31476\&\N__31727\&\N__31909\&\N__32100\&\N__32297\&\N__32633\&\N__32782\;
    \this_spr_ram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__34565\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__29427\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus4_1\ <= \this_spr_ram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus4_0\ <= \this_spr_ram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_4_0_physical_RADDR_wire\ <= \N__19509\&\N__19682\&\N__19922\&\N__18899\&\N__38039\&\N__14262\&\N__14364\&\N__20115\&\N__20572\&\N__20757\&\N__21116\;
    \this_spr_ram.mem_mem_4_0_physical_WADDR_wire\ <= \N__33402\&\N__33620\&\N__33849\&\N__31295\&\N__31514\&\N__31728\&\N__31910\&\N__32138\&\N__32331\&\N__32609\&\N__32783\;
    \this_spr_ram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__35918\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28093\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus4_3\ <= \this_spr_ram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus4_2\ <= \this_spr_ram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_4_1_physical_RADDR_wire\ <= \N__19485\&\N__19681\&\N__19886\&\N__18895\&\N__38037\&\N__14263\&\N__14458\&\N__20111\&\N__20610\&\N__20802\&\N__21135\;
    \this_spr_ram.mem_mem_4_1_physical_WADDR_wire\ <= \N__33431\&\N__33650\&\N__33876\&\N__31296\&\N__31515\&\N__31746\&\N__31911\&\N__32139\&\N__32332\&\N__32641\&\N__32815\;
    \this_spr_ram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__34528\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__29418\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus5_1\ <= \this_spr_ram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus5_0\ <= \this_spr_ram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_5_0_physical_RADDR_wire\ <= \N__19486\&\N__19692\&\N__19918\&\N__18896\&\N__37997\&\N__14264\&\N__14459\&\N__20112\&\N__20639\&\N__20803\&\N__21084\;
    \this_spr_ram.mem_mem_5_0_physical_WADDR_wire\ <= \N__33430\&\N__33651\&\N__33856\&\N__31323\&\N__31538\&\N__31747\&\N__31940\&\N__32166\&\N__32360\&\N__32637\&\N__32816\;
    \this_spr_ram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__35914\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28081\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus5_3\ <= \this_spr_ram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus5_2\ <= \this_spr_ram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_5_1_physical_RADDR_wire\ <= \N__19496\&\N__19693\&\N__19923\&\N__18897\&\N__38038\&\N__14265\&\N__14480\&\N__20113\&\N__20640\&\N__20829\&\N__21083\;
    \this_spr_ram.mem_mem_5_1_physical_WADDR_wire\ <= \N__33453\&\N__33669\&\N__33890\&\N__31324\&\N__31539\&\N__31714\&\N__31941\&\N__32170\&\N__32361\&\N__32630\&\N__32837\;
    \this_spr_ram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__34566\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__29375\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus6_1\ <= \this_spr_ram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus6_0\ <= \this_spr_ram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_6_0_physical_RADDR_wire\ <= \N__19497\&\N__19694\&\N__19936\&\N__18898\&\N__38068\&\N__14266\&\N__14481\&\N__20114\&\N__20641\&\N__20830\&\N__21082\;
    \this_spr_ram.mem_mem_6_0_physical_WADDR_wire\ <= \N__33444\&\N__33678\&\N__33880\&\N__31339\&\N__31546\&\N__31736\&\N__31961\&\N__32182\&\N__32379\&\N__32623\&\N__32838\;
    \this_spr_ram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__35949\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28080\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus6_3\ <= \this_spr_ram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus6_2\ <= \this_spr_ram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_6_1_physical_RADDR_wire\ <= \N__19480\&\N__19704\&\N__19843\&\N__18850\&\N__38097\&\N__14257\&\N__14385\&\N__20104\&\N__20632\&\N__20810\&\N__21127\;
    \this_spr_ram.mem_mem_6_1_physical_WADDR_wire\ <= \N__33452\&\N__33662\&\N__33885\&\N__31340\&\N__31533\&\N__31748\&\N__31966\&\N__32183\&\N__32372\&\N__32634\&\N__32830\;
    \this_spr_ram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__34578\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__29407\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus7_1\ <= \this_spr_ram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus7_0\ <= \this_spr_ram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_7_0_physical_RADDR_wire\ <= \N__19481\&\N__19705\&\N__19844\&\N__18894\&\N__38106\&\N__14258\&\N__14386\&\N__20130\&\N__20565\&\N__20831\&\N__21128\;
    \this_spr_ram.mem_mem_7_0_physical_WADDR_wire\ <= \N__33448\&\N__33674\&\N__33886\&\N__31347\&\N__31534\&\N__31755\&\N__31970\&\N__32187\&\N__32391\&\N__32635\&\N__32843\;
    \this_spr_ram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__35964\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28114\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus7_3\ <= \this_spr_ram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus7_2\ <= \this_spr_ram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_7_1_physical_RADDR_wire\ <= \N__19508\&\N__19716\&\N__19885\&\N__18854\&\N__38107\&\N__14281\&\N__14416\&\N__20131\&\N__20652\&\N__20832\&\N__21139\;
    \this_spr_ram.mem_mem_7_1_physical_WADDR_wire\ <= \N__33454\&\N__33679\&\N__33892\&\N__31348\&\N__31545\&\N__31756\&\N__31972\&\N__32188\&\N__32395\&\N__32636\&\N__32844\;
    \this_spr_ram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__34582\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__29422\&'0'&'0'&'0';
    \M_this_vram_read_data_3\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_vram_read_data_2\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_vram_read_data_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_vram_read_data_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__23854\&\N__15466\&\N__18043\&\N__17539\&\N__16012\&\N__14839\&\N__16078\&\N__15883\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__22411\&\N__22267\&\N__22294\&\N__22330\&\N__23179\&\N__22243\&\N__23545\&\N__23512\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__34405\&\N__33979\&\N__34330\&\N__23125\;

    \this_map_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42140\,
            RE => \N__25236\,
            WCLKE => \N__40149\,
            WCLK => \N__42141\,
            WE => \N__25255\
        );

    \this_map_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42144\,
            RE => \N__25259\,
            WCLKE => \N__40156\,
            WCLK => \N__42145\,
            WE => \N__25264\
        );

    \this_oam_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42117\,
            RE => \N__24986\,
            WCLKE => \N__26758\,
            WCLK => \N__42118\,
            WE => \N__24991\
        );

    \this_oam_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42127\,
            RE => \N__24987\,
            WCLKE => \N__26757\,
            WCLK => \N__42128\,
            WE => \N__25133\
        );

    \this_ppu.oam_cache.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_ppu.oam_cache.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_ppu.oam_cache.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_ppu.oam_cache.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_ppu.oam_cache.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42060\,
            RE => \N__24833\,
            WCLKE => \N__24184\,
            WCLK => \N__42061\,
            WE => \N__24906\
        );

    \this_ppu.oam_cache.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_ppu.oam_cache.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_ppu.oam_cache.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_ppu.oam_cache.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_ppu.oam_cache.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42084\,
            RE => \N__24852\,
            WCLKE => \N__24141\,
            WCLK => \N__42085\,
            WE => \N__24907\
        );

    \this_spr_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__41984\,
            RE => \N__25263\,
            WCLKE => \N__38323\,
            WCLK => \N__41985\,
            WE => \N__25262\
        );

    \this_spr_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__41986\,
            RE => \N__25261\,
            WCLKE => \N__38322\,
            WCLK => \N__41987\,
            WE => \N__25247\
        );

    \this_spr_ram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__41988\,
            RE => \N__25251\,
            WCLKE => \N__38365\,
            WCLK => \N__41989\,
            WE => \N__25243\
        );

    \this_spr_ram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__41996\,
            RE => \N__25138\,
            WCLKE => \N__38364\,
            WCLK => \N__41995\,
            WE => \N__25220\
        );

    \this_spr_ram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42013\,
            RE => \N__25206\,
            WCLKE => \N__39184\,
            WCLK => \N__42014\,
            WE => \N__25219\
        );

    \this_spr_ram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42029\,
            RE => \N__25205\,
            WCLKE => \N__39180\,
            WCLK => \N__42030\,
            WE => \N__25164\
        );

    \this_spr_ram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42047\,
            RE => \N__25083\,
            WCLKE => \N__38346\,
            WCLK => \N__42048\,
            WE => \N__25142\
        );

    \this_spr_ram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42071\,
            RE => \N__25076\,
            WCLKE => \N__38347\,
            WCLK => \N__42072\,
            WE => \N__25084\
        );

    \this_spr_ram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42094\,
            RE => \N__25203\,
            WCLKE => \N__38961\,
            WCLK => \N__42095\,
            WE => \N__25110\
        );

    \this_spr_ram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42110\,
            RE => \N__25204\,
            WCLKE => \N__38962\,
            WCLK => \N__42111\,
            WE => \N__25176\
        );

    \this_spr_ram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42121\,
            RE => \N__25059\,
            WCLKE => \N__38943\,
            WCLK => \N__42122\,
            WE => \N__25177\
        );

    \this_spr_ram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42130\,
            RE => \N__25060\,
            WCLKE => \N__38944\,
            WCLK => \N__42131\,
            WE => \N__25227\
        );

    \this_spr_ram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42135\,
            RE => \N__25235\,
            WCLKE => \N__38646\,
            WCLK => \N__42136\,
            WE => \N__25228\
        );

    \this_spr_ram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42133\,
            RE => \N__24999\,
            WCLKE => \N__38650\,
            WCLK => \N__42134\,
            WE => \N__25134\
        );

    \this_spr_ram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42138\,
            RE => \N__25061\,
            WCLKE => \N__36702\,
            WCLK => \N__42139\,
            WE => \N__25071\
        );

    \this_spr_ram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42142\,
            RE => \N__25072\,
            WCLKE => \N__36706\,
            WCLK => \N__42143\,
            WE => \N__25199\
        );

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__42103\,
            RE => \N__24923\,
            WCLKE => \N__23035\,
            WCLK => \N__42104\,
            WE => \N__24870\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__44414\,
            GLOBALBUFFEROUTPUT => clk_0_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44416\,
            DIN => \N__44415\,
            DOUT => \N__44414\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__44416\,
            PADOUT => \N__44415\,
            PADIN => \N__44414\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44405\,
            DIN => \N__44404\,
            DOUT => \N__44403\,
            PACKAGEPIN => debug_wire(0)
        );

    \debug_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44405\,
            PADOUT => \N__44404\,
            PADIN => \N__44403\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44396\,
            DIN => \N__44395\,
            DOUT => \N__44394\,
            PACKAGEPIN => debug_wire(1)
        );

    \debug_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44396\,
            PADOUT => \N__44395\,
            PADIN => \N__44394\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44387\,
            DIN => \N__44386\,
            DOUT => \N__44385\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44387\,
            PADOUT => \N__44386\,
            PADIN => \N__44385\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14569\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44378\,
            DIN => \N__44377\,
            DOUT => \N__44376\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44378\,
            PADOUT => \N__44377\,
            PADIN => \N__44376\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__16306\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44369\,
            DIN => \N__44368\,
            DOUT => \N__44367\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44369\,
            PADOUT => \N__44368\,
            PADIN => \N__44367\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__25260\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44360\,
            DIN => \N__44359\,
            DOUT => \N__44358\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44360\,
            PADOUT => \N__44359\,
            PADIN => \N__44358\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__35863\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44351\,
            DIN => \N__44350\,
            DOUT => \N__44349\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44351\,
            PADOUT => \N__44350\,
            PADIN => \N__44349\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44342\,
            DIN => \N__44341\,
            DOUT => \N__44340\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44342\,
            PADOUT => \N__44341\,
            PADIN => \N__44340\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44333\,
            DIN => \N__44332\,
            DOUT => \N__44331\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44333\,
            PADOUT => \N__44332\,
            PADIN => \N__44331\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44324\,
            DIN => \N__44323\,
            DOUT => \N__44322\,
            PACKAGEPIN => led_wire(5)
        );

    \led_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44324\,
            PADOUT => \N__44323\,
            PADIN => \N__44322\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__36064\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44315\,
            DIN => \N__44314\,
            DOUT => \N__44313\,
            PACKAGEPIN => led_wire(6)
        );

    \led_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44315\,
            PADOUT => \N__44314\,
            PADIN => \N__44313\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37360\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44306\,
            DIN => \N__44305\,
            DOUT => \N__44304\,
            PACKAGEPIN => led_wire(7)
        );

    \led_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44306\,
            PADOUT => \N__44305\,
            PADIN => \N__44304\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__30871\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44297\,
            DIN => \N__44296\,
            DOUT => \N__44295\,
            PACKAGEPIN => port_address(0)
        );

    \port_address_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44297\,
            PADOUT => \N__44296\,
            PADIN => \N__44295\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__40291\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37607\
        );

    \port_address_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44288\,
            DIN => \N__44287\,
            DOUT => \N__44286\,
            PACKAGEPIN => port_address(1)
        );

    \port_address_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44288\,
            PADOUT => \N__44287\,
            PADIN => \N__44286\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__41305\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37585\
        );

    \port_address_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44279\,
            DIN => \N__44278\,
            DOUT => \N__44277\,
            PACKAGEPIN => port_address(2)
        );

    \port_address_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44279\,
            PADOUT => \N__44278\,
            PADIN => \N__44277\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__40246\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37576\
        );

    \port_address_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44270\,
            DIN => \N__44269\,
            DOUT => \N__44268\,
            PACKAGEPIN => port_address(3)
        );

    \port_address_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44270\,
            PADOUT => \N__44269\,
            PADIN => \N__44268\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__41266\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37622\
        );

    \port_address_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44261\,
            DIN => \N__44260\,
            DOUT => \N__44259\,
            PACKAGEPIN => port_address(4)
        );

    \port_address_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44261\,
            PADOUT => \N__44260\,
            PADIN => \N__44259\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__41227\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37611\
        );

    \port_address_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44252\,
            DIN => \N__44251\,
            DOUT => \N__44250\,
            PACKAGEPIN => port_address(5)
        );

    \port_address_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44252\,
            PADOUT => \N__44251\,
            PADIN => \N__44250\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__41191\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37561\
        );

    \port_address_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44243\,
            DIN => \N__44242\,
            DOUT => \N__44241\,
            PACKAGEPIN => port_address(6)
        );

    \port_address_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44243\,
            PADOUT => \N__44242\,
            PADIN => \N__44241\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__43279\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37606\
        );

    \port_address_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44234\,
            DIN => \N__44233\,
            DOUT => \N__44232\,
            PACKAGEPIN => port_address(7)
        );

    \port_address_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44234\,
            PADOUT => \N__44233\,
            PADIN => \N__44232\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__40984\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37639\
        );

    \port_address_obuft_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44225\,
            DIN => \N__44224\,
            DOUT => \N__44223\,
            PACKAGEPIN => port_address(10)
        );

    \port_address_obuft_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44225\,
            PADOUT => \N__44224\,
            PADIN => \N__44223\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__41020\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37577\
        );

    \port_address_obuft_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44216\,
            DIN => \N__44215\,
            DOUT => \N__44214\,
            PACKAGEPIN => port_address(11)
        );

    \port_address_obuft_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44216\,
            PADOUT => \N__44215\,
            PADIN => \N__44214\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__40942\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37609\
        );

    \port_address_obuft_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44207\,
            DIN => \N__44206\,
            DOUT => \N__44205\,
            PACKAGEPIN => port_address(12)
        );

    \port_address_obuft_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44207\,
            PADOUT => \N__44206\,
            PADIN => \N__44205\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__40912\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37612\
        );

    \port_address_obuft_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44198\,
            DIN => \N__44197\,
            DOUT => \N__44196\,
            PACKAGEPIN => port_address(13)
        );

    \port_address_obuft_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44198\,
            PADOUT => \N__44197\,
            PADIN => \N__44196\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__40582\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37562\
        );

    \port_address_obuft_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44189\,
            DIN => \N__44188\,
            DOUT => \N__44187\,
            PACKAGEPIN => port_address(14)
        );

    \port_address_obuft_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44189\,
            PADOUT => \N__44188\,
            PADIN => \N__44187\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__40543\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37623\
        );

    \port_address_obuft_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44180\,
            DIN => \N__44179\,
            DOUT => \N__44178\,
            PACKAGEPIN => port_address(15)
        );

    \port_address_obuft_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44180\,
            PADOUT => \N__44179\,
            PADIN => \N__44178\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__40507\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37635\
        );

    \port_address_obuft_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44171\,
            DIN => \N__44170\,
            DOUT => \N__44169\,
            PACKAGEPIN => port_address(8)
        );

    \port_address_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44171\,
            PADOUT => \N__44170\,
            PADIN => \N__44169\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__41335\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37608\
        );

    \port_address_obuft_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44162\,
            DIN => \N__44161\,
            DOUT => \N__44160\,
            PACKAGEPIN => port_address(9)
        );

    \port_address_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44162\,
            PADOUT => \N__44161\,
            PADIN => \N__44160\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__40636\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37584\
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44153\,
            DIN => \N__44152\,
            DOUT => \N__44151\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__44153\,
            PADOUT => \N__44152\,
            PADIN => \N__44151\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44144\,
            DIN => \N__44143\,
            DOUT => \N__44142\,
            PACKAGEPIN => port_data(0)
        );

    \port_data_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44144\,
            PADOUT => \N__44143\,
            PADIN => \N__44142\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__21787\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__38437\
        );

    \port_data_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44135\,
            DIN => \N__44134\,
            DOUT => \N__44133\,
            PACKAGEPIN => port_data(1)
        );

    \port_data_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44135\,
            PADOUT => \N__44134\,
            PADIN => \N__44133\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__20173\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__38438\
        );

    \port_data_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44126\,
            DIN => \N__44125\,
            DOUT => \N__44124\,
            PACKAGEPIN => port_data(2)
        );

    \port_data_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44126\,
            PADOUT => \N__44125\,
            PADIN => \N__44124\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__41350\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__38401\
        );

    \port_data_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44117\,
            DIN => \N__44116\,
            DOUT => \N__44115\,
            PACKAGEPIN => port_data(3)
        );

    \port_data_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44117\,
            PADOUT => \N__44116\,
            PADIN => \N__44115\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__43588\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__38413\
        );

    \port_data_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44108\,
            DIN => \N__44107\,
            DOUT => \N__44106\,
            PACKAGEPIN => port_data(4)
        );

    \port_data_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44108\,
            PADOUT => \N__44107\,
            PADIN => \N__44106\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__43714\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__38431\
        );

    \port_data_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44099\,
            DIN => \N__44098\,
            DOUT => \N__44097\,
            PACKAGEPIN => port_data(5)
        );

    \port_data_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44099\,
            PADOUT => \N__44098\,
            PADIN => \N__44097\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__43903\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__38445\
        );

    \port_data_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44090\,
            DIN => \N__44089\,
            DOUT => \N__44088\,
            PACKAGEPIN => port_data(6)
        );

    \port_data_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44090\,
            PADOUT => \N__44089\,
            PADIN => \N__44088\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__41575\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__38457\
        );

    \port_data_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44081\,
            DIN => \N__44080\,
            DOUT => \N__44079\,
            PACKAGEPIN => port_data(7)
        );

    \port_data_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44081\,
            PADOUT => \N__44080\,
            PADIN => \N__44079\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__38983\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__38461\
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44072\,
            DIN => \N__44071\,
            DOUT => \N__44070\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44072\,
            PADOUT => \N__44071\,
            PADIN => \N__44070\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14062\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44063\,
            DIN => \N__44062\,
            DOUT => \N__44061\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44063\,
            PADOUT => \N__44062\,
            PADIN => \N__44061\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37762\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44054\,
            DIN => \N__44053\,
            DOUT => \N__44052\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__44054\,
            PADOUT => \N__44053\,
            PADIN => \N__44052\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44045\,
            DIN => \N__44044\,
            DOUT => \N__44043\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44045\,
            PADOUT => \N__44044\,
            PADIN => \N__44043\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14020\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44036\,
            DIN => \N__44035\,
            DOUT => \N__44034\,
            PACKAGEPIN => port_rw
        );

    \port_rw_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__44036\,
            PADOUT => \N__44035\,
            PADIN => \N__44034\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_in,
            DIN1 => OPEN,
            DOUT0 => \N__24869\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__37610\
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44027\,
            DIN => \N__44026\,
            DOUT => \N__44025\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44027\,
            PADOUT => \N__44026\,
            PADIN => \N__44025\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14770\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44018\,
            DIN => \N__44017\,
            DOUT => \N__44016\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44018\,
            PADOUT => \N__44017\,
            PADIN => \N__44016\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__15349\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44009\,
            DIN => \N__44008\,
            DOUT => \N__44007\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44009\,
            PADOUT => \N__44008\,
            PADIN => \N__44007\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13978\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__44000\,
            DIN => \N__43999\,
            DOUT => \N__43998\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__44000\,
            PADOUT => \N__43999\,
            PADIN => \N__43998\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__16699\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__43991\,
            DIN => \N__43990\,
            DOUT => \N__43989\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__43991\,
            PADOUT => \N__43990\,
            PADIN => \N__43989\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14044\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__43982\,
            DIN => \N__43981\,
            DOUT => \N__43980\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__43982\,
            PADOUT => \N__43981\,
            PADIN => \N__43980\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14551\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__43973\,
            DIN => \N__43972\,
            DOUT => \N__43971\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__43973\,
            PADOUT => \N__43972\,
            PADIN => \N__43971\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__43964\,
            DIN => \N__43963\,
            DOUT => \N__43962\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__43964\,
            PADOUT => \N__43963\,
            PADIN => \N__43962\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14056\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__43955\,
            DIN => \N__43954\,
            DOUT => \N__43953\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__43955\,
            PADOUT => \N__43954\,
            PADIN => \N__43953\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__22441\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__11033\ : InMux
    port map (
            O => \N__43936\,
            I => \N__43932\
        );

    \I__11032\ : InMux
    port map (
            O => \N__43935\,
            I => \N__43929\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__43932\,
            I => \N__43926\
        );

    \I__11030\ : LocalMux
    port map (
            O => \N__43929\,
            I => \N__43923\
        );

    \I__11029\ : Span4Mux_v
    port map (
            O => \N__43926\,
            I => \N__43920\
        );

    \I__11028\ : Span4Mux_h
    port map (
            O => \N__43923\,
            I => \N__43917\
        );

    \I__11027\ : Span4Mux_h
    port map (
            O => \N__43920\,
            I => \N__43912\
        );

    \I__11026\ : Span4Mux_v
    port map (
            O => \N__43917\,
            I => \N__43912\
        );

    \I__11025\ : Span4Mux_v
    port map (
            O => \N__43912\,
            I => \N__43909\
        );

    \I__11024\ : Span4Mux_v
    port map (
            O => \N__43909\,
            I => \N__43906\
        );

    \I__11023\ : Odrv4
    port map (
            O => \N__43906\,
            I => \M_this_map_ram_read_data_5\
        );

    \I__11022\ : IoInMux
    port map (
            O => \N__43903\,
            I => \N__43900\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__43900\,
            I => \N__43897\
        );

    \I__11020\ : Odrv12
    port map (
            O => \N__43897\,
            I => \N_996_0\
        );

    \I__11019\ : CascadeMux
    port map (
            O => \N__43894\,
            I => \N__43891\
        );

    \I__11018\ : InMux
    port map (
            O => \N__43891\,
            I => \N__43888\
        );

    \I__11017\ : LocalMux
    port map (
            O => \N__43888\,
            I => \N__43884\
        );

    \I__11016\ : CascadeMux
    port map (
            O => \N__43887\,
            I => \N__43881\
        );

    \I__11015\ : Span4Mux_h
    port map (
            O => \N__43884\,
            I => \N__43878\
        );

    \I__11014\ : InMux
    port map (
            O => \N__43881\,
            I => \N__43875\
        );

    \I__11013\ : Span4Mux_h
    port map (
            O => \N__43878\,
            I => \N__43869\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__43875\,
            I => \N__43869\
        );

    \I__11011\ : InMux
    port map (
            O => \N__43874\,
            I => \N__43866\
        );

    \I__11010\ : Sp12to4
    port map (
            O => \N__43869\,
            I => \N__43861\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__43866\,
            I => \N__43861\
        );

    \I__11008\ : Span12Mux_v
    port map (
            O => \N__43861\,
            I => \N__43858\
        );

    \I__11007\ : Odrv12
    port map (
            O => \N__43858\,
            I => port_address_in_6
        );

    \I__11006\ : InMux
    port map (
            O => \N__43855\,
            I => \N__43851\
        );

    \I__11005\ : InMux
    port map (
            O => \N__43854\,
            I => \N__43848\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__43851\,
            I => \N__43844\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__43848\,
            I => \N__43841\
        );

    \I__11002\ : InMux
    port map (
            O => \N__43847\,
            I => \N__43838\
        );

    \I__11001\ : Span4Mux_v
    port map (
            O => \N__43844\,
            I => \N__43835\
        );

    \I__11000\ : Span4Mux_v
    port map (
            O => \N__43841\,
            I => \N__43832\
        );

    \I__10999\ : LocalMux
    port map (
            O => \N__43838\,
            I => \N__43829\
        );

    \I__10998\ : Sp12to4
    port map (
            O => \N__43835\,
            I => \N__43826\
        );

    \I__10997\ : Span4Mux_h
    port map (
            O => \N__43832\,
            I => \N__43823\
        );

    \I__10996\ : Span4Mux_v
    port map (
            O => \N__43829\,
            I => \N__43820\
        );

    \I__10995\ : Odrv12
    port map (
            O => \N__43826\,
            I => port_address_in_5
        );

    \I__10994\ : Odrv4
    port map (
            O => \N__43823\,
            I => port_address_in_5
        );

    \I__10993\ : Odrv4
    port map (
            O => \N__43820\,
            I => port_address_in_5
        );

    \I__10992\ : InMux
    port map (
            O => \N__43813\,
            I => \N__43810\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__43810\,
            I => \N__43807\
        );

    \I__10990\ : Span4Mux_v
    port map (
            O => \N__43807\,
            I => \N__43803\
        );

    \I__10989\ : InMux
    port map (
            O => \N__43806\,
            I => \N__43800\
        );

    \I__10988\ : Span4Mux_h
    port map (
            O => \N__43803\,
            I => \N__43796\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__43800\,
            I => \N__43793\
        );

    \I__10986\ : InMux
    port map (
            O => \N__43799\,
            I => \N__43790\
        );

    \I__10985\ : Span4Mux_v
    port map (
            O => \N__43796\,
            I => \N__43787\
        );

    \I__10984\ : Span4Mux_h
    port map (
            O => \N__43793\,
            I => \N__43784\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__43790\,
            I => \N__43781\
        );

    \I__10982\ : Sp12to4
    port map (
            O => \N__43787\,
            I => \N__43778\
        );

    \I__10981\ : Sp12to4
    port map (
            O => \N__43784\,
            I => \N__43775\
        );

    \I__10980\ : Span12Mux_v
    port map (
            O => \N__43781\,
            I => \N__43772\
        );

    \I__10979\ : Span12Mux_s2_h
    port map (
            O => \N__43778\,
            I => \N__43767\
        );

    \I__10978\ : Span12Mux_v
    port map (
            O => \N__43775\,
            I => \N__43767\
        );

    \I__10977\ : Span12Mux_v
    port map (
            O => \N__43772\,
            I => \N__43764\
        );

    \I__10976\ : Span12Mux_v
    port map (
            O => \N__43767\,
            I => \N__43761\
        );

    \I__10975\ : Odrv12
    port map (
            O => \N__43764\,
            I => port_address_in_7
        );

    \I__10974\ : Odrv12
    port map (
            O => \N__43761\,
            I => port_address_in_7
        );

    \I__10973\ : InMux
    port map (
            O => \N__43756\,
            I => \N__43753\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__43753\,
            I => \N__43750\
        );

    \I__10971\ : Odrv12
    port map (
            O => \N__43750\,
            I => \M_this_substate_d_0_sqmuxa_3_0_o2_x\
        );

    \I__10970\ : InMux
    port map (
            O => \N__43747\,
            I => \N__43743\
        );

    \I__10969\ : InMux
    port map (
            O => \N__43746\,
            I => \N__43740\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__43743\,
            I => \N__43737\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__43740\,
            I => \N__43734\
        );

    \I__10966\ : Span4Mux_h
    port map (
            O => \N__43737\,
            I => \N__43731\
        );

    \I__10965\ : Span4Mux_v
    port map (
            O => \N__43734\,
            I => \N__43728\
        );

    \I__10964\ : Sp12to4
    port map (
            O => \N__43731\,
            I => \N__43725\
        );

    \I__10963\ : Span4Mux_v
    port map (
            O => \N__43728\,
            I => \N__43722\
        );

    \I__10962\ : Span12Mux_v
    port map (
            O => \N__43725\,
            I => \N__43719\
        );

    \I__10961\ : Odrv4
    port map (
            O => \N__43722\,
            I => \M_this_map_ram_read_data_4\
        );

    \I__10960\ : Odrv12
    port map (
            O => \N__43719\,
            I => \M_this_map_ram_read_data_4\
        );

    \I__10959\ : IoInMux
    port map (
            O => \N__43714\,
            I => \N__43711\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__43711\,
            I => \N__43708\
        );

    \I__10957\ : Odrv12
    port map (
            O => \N__43708\,
            I => \N_730_0\
        );

    \I__10956\ : InMux
    port map (
            O => \N__43705\,
            I => \N__43700\
        );

    \I__10955\ : InMux
    port map (
            O => \N__43704\,
            I => \N__43697\
        );

    \I__10954\ : InMux
    port map (
            O => \N__43703\,
            I => \N__43692\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__43700\,
            I => \N__43687\
        );

    \I__10952\ : LocalMux
    port map (
            O => \N__43697\,
            I => \N__43687\
        );

    \I__10951\ : InMux
    port map (
            O => \N__43696\,
            I => \N__43682\
        );

    \I__10950\ : InMux
    port map (
            O => \N__43695\,
            I => \N__43682\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__43692\,
            I => \N__43678\
        );

    \I__10948\ : Span4Mux_v
    port map (
            O => \N__43687\,
            I => \N__43675\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__43682\,
            I => \N__43672\
        );

    \I__10946\ : InMux
    port map (
            O => \N__43681\,
            I => \N__43669\
        );

    \I__10945\ : Span4Mux_v
    port map (
            O => \N__43678\,
            I => \N__43666\
        );

    \I__10944\ : Span4Mux_v
    port map (
            O => \N__43675\,
            I => \N__43659\
        );

    \I__10943\ : Span4Mux_v
    port map (
            O => \N__43672\,
            I => \N__43659\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__43669\,
            I => \N__43656\
        );

    \I__10941\ : Span4Mux_h
    port map (
            O => \N__43666\,
            I => \N__43653\
        );

    \I__10940\ : InMux
    port map (
            O => \N__43665\,
            I => \N__43650\
        );

    \I__10939\ : InMux
    port map (
            O => \N__43664\,
            I => \N__43647\
        );

    \I__10938\ : Span4Mux_h
    port map (
            O => \N__43659\,
            I => \N__43642\
        );

    \I__10937\ : Span4Mux_v
    port map (
            O => \N__43656\,
            I => \N__43642\
        );

    \I__10936\ : Span4Mux_h
    port map (
            O => \N__43653\,
            I => \N__43639\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__43650\,
            I => \N__43636\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__43647\,
            I => \N__43633\
        );

    \I__10933\ : Sp12to4
    port map (
            O => \N__43642\,
            I => \N__43630\
        );

    \I__10932\ : Span4Mux_h
    port map (
            O => \N__43639\,
            I => \N__43623\
        );

    \I__10931\ : Span4Mux_v
    port map (
            O => \N__43636\,
            I => \N__43623\
        );

    \I__10930\ : Span4Mux_v
    port map (
            O => \N__43633\,
            I => \N__43623\
        );

    \I__10929\ : Span12Mux_h
    port map (
            O => \N__43630\,
            I => \N__43620\
        );

    \I__10928\ : Span4Mux_v
    port map (
            O => \N__43623\,
            I => \N__43617\
        );

    \I__10927\ : Odrv12
    port map (
            O => \N__43620\,
            I => \this_vga_signals.N_834_0\
        );

    \I__10926\ : Odrv4
    port map (
            O => \N__43617\,
            I => \this_vga_signals.N_834_0\
        );

    \I__10925\ : InMux
    port map (
            O => \N__43612\,
            I => \N__43609\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__43609\,
            I => \N__43605\
        );

    \I__10923\ : InMux
    port map (
            O => \N__43608\,
            I => \N__43602\
        );

    \I__10922\ : Span12Mux_v
    port map (
            O => \N__43605\,
            I => \N__43599\
        );

    \I__10921\ : LocalMux
    port map (
            O => \N__43602\,
            I => \N__43596\
        );

    \I__10920\ : Span12Mux_h
    port map (
            O => \N__43599\,
            I => \N__43593\
        );

    \I__10919\ : Odrv4
    port map (
            O => \N__43596\,
            I => \M_this_map_ram_read_data_3\
        );

    \I__10918\ : Odrv12
    port map (
            O => \N__43593\,
            I => \M_this_map_ram_read_data_3\
        );

    \I__10917\ : IoInMux
    port map (
            O => \N__43588\,
            I => \N__43585\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__43585\,
            I => \N__43582\
        );

    \I__10915\ : Span4Mux_s1_v
    port map (
            O => \N__43582\,
            I => \N__43579\
        );

    \I__10914\ : Odrv4
    port map (
            O => \N__43579\,
            I => \N_728_0\
        );

    \I__10913\ : CascadeMux
    port map (
            O => \N__43576\,
            I => \N__43569\
        );

    \I__10912\ : CascadeMux
    port map (
            O => \N__43575\,
            I => \N__43558\
        );

    \I__10911\ : CascadeMux
    port map (
            O => \N__43574\,
            I => \N__43555\
        );

    \I__10910\ : CascadeMux
    port map (
            O => \N__43573\,
            I => \N__43552\
        );

    \I__10909\ : CascadeMux
    port map (
            O => \N__43572\,
            I => \N__43549\
        );

    \I__10908\ : InMux
    port map (
            O => \N__43569\,
            I => \N__43530\
        );

    \I__10907\ : InMux
    port map (
            O => \N__43568\,
            I => \N__43530\
        );

    \I__10906\ : InMux
    port map (
            O => \N__43567\,
            I => \N__43530\
        );

    \I__10905\ : InMux
    port map (
            O => \N__43566\,
            I => \N__43530\
        );

    \I__10904\ : InMux
    port map (
            O => \N__43565\,
            I => \N__43530\
        );

    \I__10903\ : InMux
    port map (
            O => \N__43564\,
            I => \N__43530\
        );

    \I__10902\ : InMux
    port map (
            O => \N__43563\,
            I => \N__43517\
        );

    \I__10901\ : InMux
    port map (
            O => \N__43562\,
            I => \N__43517\
        );

    \I__10900\ : InMux
    port map (
            O => \N__43561\,
            I => \N__43517\
        );

    \I__10899\ : InMux
    port map (
            O => \N__43558\,
            I => \N__43517\
        );

    \I__10898\ : InMux
    port map (
            O => \N__43555\,
            I => \N__43517\
        );

    \I__10897\ : InMux
    port map (
            O => \N__43552\,
            I => \N__43504\
        );

    \I__10896\ : InMux
    port map (
            O => \N__43549\,
            I => \N__43504\
        );

    \I__10895\ : InMux
    port map (
            O => \N__43548\,
            I => \N__43504\
        );

    \I__10894\ : InMux
    port map (
            O => \N__43547\,
            I => \N__43504\
        );

    \I__10893\ : InMux
    port map (
            O => \N__43546\,
            I => \N__43504\
        );

    \I__10892\ : InMux
    port map (
            O => \N__43545\,
            I => \N__43504\
        );

    \I__10891\ : InMux
    port map (
            O => \N__43544\,
            I => \N__43496\
        );

    \I__10890\ : InMux
    port map (
            O => \N__43543\,
            I => \N__43493\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__43530\,
            I => \N__43490\
        );

    \I__10888\ : CascadeMux
    port map (
            O => \N__43529\,
            I => \N__43481\
        );

    \I__10887\ : InMux
    port map (
            O => \N__43528\,
            I => \N__43478\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__43517\,
            I => \N__43475\
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__43504\,
            I => \N__43472\
        );

    \I__10884\ : InMux
    port map (
            O => \N__43503\,
            I => \N__43467\
        );

    \I__10883\ : InMux
    port map (
            O => \N__43502\,
            I => \N__43464\
        );

    \I__10882\ : InMux
    port map (
            O => \N__43501\,
            I => \N__43461\
        );

    \I__10881\ : InMux
    port map (
            O => \N__43500\,
            I => \N__43457\
        );

    \I__10880\ : InMux
    port map (
            O => \N__43499\,
            I => \N__43454\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__43496\,
            I => \N__43447\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__43493\,
            I => \N__43447\
        );

    \I__10877\ : Span4Mux_h
    port map (
            O => \N__43490\,
            I => \N__43447\
        );

    \I__10876\ : InMux
    port map (
            O => \N__43489\,
            I => \N__43440\
        );

    \I__10875\ : InMux
    port map (
            O => \N__43488\,
            I => \N__43440\
        );

    \I__10874\ : InMux
    port map (
            O => \N__43487\,
            I => \N__43440\
        );

    \I__10873\ : InMux
    port map (
            O => \N__43486\,
            I => \N__43433\
        );

    \I__10872\ : InMux
    port map (
            O => \N__43485\,
            I => \N__43433\
        );

    \I__10871\ : InMux
    port map (
            O => \N__43484\,
            I => \N__43433\
        );

    \I__10870\ : InMux
    port map (
            O => \N__43481\,
            I => \N__43428\
        );

    \I__10869\ : LocalMux
    port map (
            O => \N__43478\,
            I => \N__43425\
        );

    \I__10868\ : Span4Mux_v
    port map (
            O => \N__43475\,
            I => \N__43420\
        );

    \I__10867\ : Span4Mux_h
    port map (
            O => \N__43472\,
            I => \N__43420\
        );

    \I__10866\ : InMux
    port map (
            O => \N__43471\,
            I => \N__43417\
        );

    \I__10865\ : InMux
    port map (
            O => \N__43470\,
            I => \N__43412\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__43467\,
            I => \N__43405\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__43464\,
            I => \N__43405\
        );

    \I__10862\ : LocalMux
    port map (
            O => \N__43461\,
            I => \N__43405\
        );

    \I__10861\ : InMux
    port map (
            O => \N__43460\,
            I => \N__43402\
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__43457\,
            I => \N__43398\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__43454\,
            I => \N__43389\
        );

    \I__10858\ : Span4Mux_v
    port map (
            O => \N__43447\,
            I => \N__43389\
        );

    \I__10857\ : LocalMux
    port map (
            O => \N__43440\,
            I => \N__43389\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__43433\,
            I => \N__43389\
        );

    \I__10855\ : InMux
    port map (
            O => \N__43432\,
            I => \N__43384\
        );

    \I__10854\ : InMux
    port map (
            O => \N__43431\,
            I => \N__43384\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__43428\,
            I => \N__43381\
        );

    \I__10852\ : Span4Mux_v
    port map (
            O => \N__43425\,
            I => \N__43378\
        );

    \I__10851\ : Span4Mux_h
    port map (
            O => \N__43420\,
            I => \N__43373\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__43417\,
            I => \N__43373\
        );

    \I__10849\ : InMux
    port map (
            O => \N__43416\,
            I => \N__43366\
        );

    \I__10848\ : InMux
    port map (
            O => \N__43415\,
            I => \N__43366\
        );

    \I__10847\ : LocalMux
    port map (
            O => \N__43412\,
            I => \N__43362\
        );

    \I__10846\ : Span4Mux_v
    port map (
            O => \N__43405\,
            I => \N__43357\
        );

    \I__10845\ : LocalMux
    port map (
            O => \N__43402\,
            I => \N__43357\
        );

    \I__10844\ : InMux
    port map (
            O => \N__43401\,
            I => \N__43351\
        );

    \I__10843\ : Span4Mux_v
    port map (
            O => \N__43398\,
            I => \N__43344\
        );

    \I__10842\ : Span4Mux_v
    port map (
            O => \N__43389\,
            I => \N__43344\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__43384\,
            I => \N__43344\
        );

    \I__10840\ : Span4Mux_v
    port map (
            O => \N__43381\,
            I => \N__43341\
        );

    \I__10839\ : Span4Mux_h
    port map (
            O => \N__43378\,
            I => \N__43338\
        );

    \I__10838\ : Span4Mux_h
    port map (
            O => \N__43373\,
            I => \N__43335\
        );

    \I__10837\ : InMux
    port map (
            O => \N__43372\,
            I => \N__43332\
        );

    \I__10836\ : InMux
    port map (
            O => \N__43371\,
            I => \N__43329\
        );

    \I__10835\ : LocalMux
    port map (
            O => \N__43366\,
            I => \N__43326\
        );

    \I__10834\ : InMux
    port map (
            O => \N__43365\,
            I => \N__43323\
        );

    \I__10833\ : Span4Mux_h
    port map (
            O => \N__43362\,
            I => \N__43318\
        );

    \I__10832\ : Span4Mux_h
    port map (
            O => \N__43357\,
            I => \N__43318\
        );

    \I__10831\ : InMux
    port map (
            O => \N__43356\,
            I => \N__43311\
        );

    \I__10830\ : InMux
    port map (
            O => \N__43355\,
            I => \N__43311\
        );

    \I__10829\ : InMux
    port map (
            O => \N__43354\,
            I => \N__43311\
        );

    \I__10828\ : LocalMux
    port map (
            O => \N__43351\,
            I => \N__43306\
        );

    \I__10827\ : Span4Mux_h
    port map (
            O => \N__43344\,
            I => \N__43306\
        );

    \I__10826\ : Odrv4
    port map (
            O => \N__43341\,
            I => \N_765_0\
        );

    \I__10825\ : Odrv4
    port map (
            O => \N__43338\,
            I => \N_765_0\
        );

    \I__10824\ : Odrv4
    port map (
            O => \N__43335\,
            I => \N_765_0\
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__43332\,
            I => \N_765_0\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__43329\,
            I => \N_765_0\
        );

    \I__10821\ : Odrv4
    port map (
            O => \N__43326\,
            I => \N_765_0\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__43323\,
            I => \N_765_0\
        );

    \I__10819\ : Odrv4
    port map (
            O => \N__43318\,
            I => \N_765_0\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__43311\,
            I => \N_765_0\
        );

    \I__10817\ : Odrv4
    port map (
            O => \N__43306\,
            I => \N_765_0\
        );

    \I__10816\ : InMux
    port map (
            O => \N__43285\,
            I => \N__43282\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__43282\,
            I => \un1_M_this_ext_address_q_cry_5_THRU_CO\
        );

    \I__10814\ : IoInMux
    port map (
            O => \N__43279\,
            I => \N__43276\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__43276\,
            I => \N__43272\
        );

    \I__10812\ : CascadeMux
    port map (
            O => \N__43275\,
            I => \N__43268\
        );

    \I__10811\ : Span12Mux_s5_h
    port map (
            O => \N__43272\,
            I => \N__43265\
        );

    \I__10810\ : InMux
    port map (
            O => \N__43271\,
            I => \N__43262\
        );

    \I__10809\ : InMux
    port map (
            O => \N__43268\,
            I => \N__43259\
        );

    \I__10808\ : Odrv12
    port map (
            O => \N__43265\,
            I => \M_this_ext_address_qZ0Z_6\
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__43262\,
            I => \M_this_ext_address_qZ0Z_6\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__43259\,
            I => \M_this_ext_address_qZ0Z_6\
        );

    \I__10805\ : CascadeMux
    port map (
            O => \N__43252\,
            I => \N__43245\
        );

    \I__10804\ : CascadeMux
    port map (
            O => \N__43251\,
            I => \N__43229\
        );

    \I__10803\ : InMux
    port map (
            O => \N__43250\,
            I => \N__43212\
        );

    \I__10802\ : InMux
    port map (
            O => \N__43249\,
            I => \N__43212\
        );

    \I__10801\ : InMux
    port map (
            O => \N__43248\,
            I => \N__43209\
        );

    \I__10800\ : InMux
    port map (
            O => \N__43245\,
            I => \N__43206\
        );

    \I__10799\ : InMux
    port map (
            O => \N__43244\,
            I => \N__43203\
        );

    \I__10798\ : InMux
    port map (
            O => \N__43243\,
            I => \N__43200\
        );

    \I__10797\ : InMux
    port map (
            O => \N__43242\,
            I => \N__43197\
        );

    \I__10796\ : InMux
    port map (
            O => \N__43241\,
            I => \N__43194\
        );

    \I__10795\ : InMux
    port map (
            O => \N__43240\,
            I => \N__43191\
        );

    \I__10794\ : InMux
    port map (
            O => \N__43239\,
            I => \N__43186\
        );

    \I__10793\ : InMux
    port map (
            O => \N__43238\,
            I => \N__43186\
        );

    \I__10792\ : InMux
    port map (
            O => \N__43237\,
            I => \N__43183\
        );

    \I__10791\ : InMux
    port map (
            O => \N__43236\,
            I => \N__43180\
        );

    \I__10790\ : InMux
    port map (
            O => \N__43235\,
            I => \N__43177\
        );

    \I__10789\ : InMux
    port map (
            O => \N__43234\,
            I => \N__43174\
        );

    \I__10788\ : InMux
    port map (
            O => \N__43233\,
            I => \N__43171\
        );

    \I__10787\ : InMux
    port map (
            O => \N__43232\,
            I => \N__43166\
        );

    \I__10786\ : InMux
    port map (
            O => \N__43229\,
            I => \N__43166\
        );

    \I__10785\ : InMux
    port map (
            O => \N__43228\,
            I => \N__43163\
        );

    \I__10784\ : InMux
    port map (
            O => \N__43227\,
            I => \N__43158\
        );

    \I__10783\ : InMux
    port map (
            O => \N__43226\,
            I => \N__43158\
        );

    \I__10782\ : InMux
    port map (
            O => \N__43225\,
            I => \N__43153\
        );

    \I__10781\ : InMux
    port map (
            O => \N__43224\,
            I => \N__43153\
        );

    \I__10780\ : InMux
    port map (
            O => \N__43223\,
            I => \N__43150\
        );

    \I__10779\ : InMux
    port map (
            O => \N__43222\,
            I => \N__43147\
        );

    \I__10778\ : InMux
    port map (
            O => \N__43221\,
            I => \N__43144\
        );

    \I__10777\ : InMux
    port map (
            O => \N__43220\,
            I => \N__43141\
        );

    \I__10776\ : InMux
    port map (
            O => \N__43219\,
            I => \N__43138\
        );

    \I__10775\ : InMux
    port map (
            O => \N__43218\,
            I => \N__43135\
        );

    \I__10774\ : InMux
    port map (
            O => \N__43217\,
            I => \N__43132\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__43212\,
            I => \N__43094\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__43209\,
            I => \N__43091\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__43206\,
            I => \N__43088\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__43203\,
            I => \N__43085\
        );

    \I__10769\ : LocalMux
    port map (
            O => \N__43200\,
            I => \N__43082\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__43197\,
            I => \N__43079\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__43194\,
            I => \N__43076\
        );

    \I__10766\ : LocalMux
    port map (
            O => \N__43191\,
            I => \N__43073\
        );

    \I__10765\ : LocalMux
    port map (
            O => \N__43186\,
            I => \N__43070\
        );

    \I__10764\ : LocalMux
    port map (
            O => \N__43183\,
            I => \N__43067\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__43180\,
            I => \N__43064\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__43177\,
            I => \N__43061\
        );

    \I__10761\ : LocalMux
    port map (
            O => \N__43174\,
            I => \N__43058\
        );

    \I__10760\ : LocalMux
    port map (
            O => \N__43171\,
            I => \N__43055\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__43166\,
            I => \N__43052\
        );

    \I__10758\ : LocalMux
    port map (
            O => \N__43163\,
            I => \N__43049\
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__43158\,
            I => \N__43046\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__43153\,
            I => \N__43043\
        );

    \I__10755\ : LocalMux
    port map (
            O => \N__43150\,
            I => \N__43040\
        );

    \I__10754\ : LocalMux
    port map (
            O => \N__43147\,
            I => \N__43037\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__43144\,
            I => \N__43034\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__43141\,
            I => \N__43031\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__43138\,
            I => \N__43028\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__43135\,
            I => \N__43025\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__43132\,
            I => \N__43022\
        );

    \I__10748\ : SRMux
    port map (
            O => \N__43131\,
            I => \N__42901\
        );

    \I__10747\ : SRMux
    port map (
            O => \N__43130\,
            I => \N__42901\
        );

    \I__10746\ : SRMux
    port map (
            O => \N__43129\,
            I => \N__42901\
        );

    \I__10745\ : SRMux
    port map (
            O => \N__43128\,
            I => \N__42901\
        );

    \I__10744\ : SRMux
    port map (
            O => \N__43127\,
            I => \N__42901\
        );

    \I__10743\ : SRMux
    port map (
            O => \N__43126\,
            I => \N__42901\
        );

    \I__10742\ : SRMux
    port map (
            O => \N__43125\,
            I => \N__42901\
        );

    \I__10741\ : SRMux
    port map (
            O => \N__43124\,
            I => \N__42901\
        );

    \I__10740\ : SRMux
    port map (
            O => \N__43123\,
            I => \N__42901\
        );

    \I__10739\ : SRMux
    port map (
            O => \N__43122\,
            I => \N__42901\
        );

    \I__10738\ : SRMux
    port map (
            O => \N__43121\,
            I => \N__42901\
        );

    \I__10737\ : SRMux
    port map (
            O => \N__43120\,
            I => \N__42901\
        );

    \I__10736\ : SRMux
    port map (
            O => \N__43119\,
            I => \N__42901\
        );

    \I__10735\ : SRMux
    port map (
            O => \N__43118\,
            I => \N__42901\
        );

    \I__10734\ : SRMux
    port map (
            O => \N__43117\,
            I => \N__42901\
        );

    \I__10733\ : SRMux
    port map (
            O => \N__43116\,
            I => \N__42901\
        );

    \I__10732\ : SRMux
    port map (
            O => \N__43115\,
            I => \N__42901\
        );

    \I__10731\ : SRMux
    port map (
            O => \N__43114\,
            I => \N__42901\
        );

    \I__10730\ : SRMux
    port map (
            O => \N__43113\,
            I => \N__42901\
        );

    \I__10729\ : SRMux
    port map (
            O => \N__43112\,
            I => \N__42901\
        );

    \I__10728\ : SRMux
    port map (
            O => \N__43111\,
            I => \N__42901\
        );

    \I__10727\ : SRMux
    port map (
            O => \N__43110\,
            I => \N__42901\
        );

    \I__10726\ : SRMux
    port map (
            O => \N__43109\,
            I => \N__42901\
        );

    \I__10725\ : SRMux
    port map (
            O => \N__43108\,
            I => \N__42901\
        );

    \I__10724\ : SRMux
    port map (
            O => \N__43107\,
            I => \N__42901\
        );

    \I__10723\ : SRMux
    port map (
            O => \N__43106\,
            I => \N__42901\
        );

    \I__10722\ : SRMux
    port map (
            O => \N__43105\,
            I => \N__42901\
        );

    \I__10721\ : SRMux
    port map (
            O => \N__43104\,
            I => \N__42901\
        );

    \I__10720\ : SRMux
    port map (
            O => \N__43103\,
            I => \N__42901\
        );

    \I__10719\ : SRMux
    port map (
            O => \N__43102\,
            I => \N__42901\
        );

    \I__10718\ : SRMux
    port map (
            O => \N__43101\,
            I => \N__42901\
        );

    \I__10717\ : SRMux
    port map (
            O => \N__43100\,
            I => \N__42901\
        );

    \I__10716\ : SRMux
    port map (
            O => \N__43099\,
            I => \N__42901\
        );

    \I__10715\ : SRMux
    port map (
            O => \N__43098\,
            I => \N__42901\
        );

    \I__10714\ : SRMux
    port map (
            O => \N__43097\,
            I => \N__42901\
        );

    \I__10713\ : Glb2LocalMux
    port map (
            O => \N__43094\,
            I => \N__42901\
        );

    \I__10712\ : Glb2LocalMux
    port map (
            O => \N__43091\,
            I => \N__42901\
        );

    \I__10711\ : Glb2LocalMux
    port map (
            O => \N__43088\,
            I => \N__42901\
        );

    \I__10710\ : Glb2LocalMux
    port map (
            O => \N__43085\,
            I => \N__42901\
        );

    \I__10709\ : Glb2LocalMux
    port map (
            O => \N__43082\,
            I => \N__42901\
        );

    \I__10708\ : Glb2LocalMux
    port map (
            O => \N__43079\,
            I => \N__42901\
        );

    \I__10707\ : Glb2LocalMux
    port map (
            O => \N__43076\,
            I => \N__42901\
        );

    \I__10706\ : Glb2LocalMux
    port map (
            O => \N__43073\,
            I => \N__42901\
        );

    \I__10705\ : Glb2LocalMux
    port map (
            O => \N__43070\,
            I => \N__42901\
        );

    \I__10704\ : Glb2LocalMux
    port map (
            O => \N__43067\,
            I => \N__42901\
        );

    \I__10703\ : Glb2LocalMux
    port map (
            O => \N__43064\,
            I => \N__42901\
        );

    \I__10702\ : Glb2LocalMux
    port map (
            O => \N__43061\,
            I => \N__42901\
        );

    \I__10701\ : Glb2LocalMux
    port map (
            O => \N__43058\,
            I => \N__42901\
        );

    \I__10700\ : Glb2LocalMux
    port map (
            O => \N__43055\,
            I => \N__42901\
        );

    \I__10699\ : Glb2LocalMux
    port map (
            O => \N__43052\,
            I => \N__42901\
        );

    \I__10698\ : Glb2LocalMux
    port map (
            O => \N__43049\,
            I => \N__42901\
        );

    \I__10697\ : Glb2LocalMux
    port map (
            O => \N__43046\,
            I => \N__42901\
        );

    \I__10696\ : Glb2LocalMux
    port map (
            O => \N__43043\,
            I => \N__42901\
        );

    \I__10695\ : Glb2LocalMux
    port map (
            O => \N__43040\,
            I => \N__42901\
        );

    \I__10694\ : Glb2LocalMux
    port map (
            O => \N__43037\,
            I => \N__42901\
        );

    \I__10693\ : Glb2LocalMux
    port map (
            O => \N__43034\,
            I => \N__42901\
        );

    \I__10692\ : Glb2LocalMux
    port map (
            O => \N__43031\,
            I => \N__42901\
        );

    \I__10691\ : Glb2LocalMux
    port map (
            O => \N__43028\,
            I => \N__42901\
        );

    \I__10690\ : Glb2LocalMux
    port map (
            O => \N__43025\,
            I => \N__42901\
        );

    \I__10689\ : Glb2LocalMux
    port map (
            O => \N__43022\,
            I => \N__42901\
        );

    \I__10688\ : GlobalMux
    port map (
            O => \N__42901\,
            I => \N__42898\
        );

    \I__10687\ : gio2CtrlBuf
    port map (
            O => \N__42898\,
            I => \M_this_reset_cond_out_g_0\
        );

    \I__10686\ : InMux
    port map (
            O => \N__42895\,
            I => \N__42892\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__42892\,
            I => \N__42889\
        );

    \I__10684\ : Odrv12
    port map (
            O => \N__42889\,
            I => \un1_M_this_map_address_q_cry_6_THRU_CO\
        );

    \I__10683\ : CascadeMux
    port map (
            O => \N__42886\,
            I => \N__42883\
        );

    \I__10682\ : CascadeBuf
    port map (
            O => \N__42883\,
            I => \N__42880\
        );

    \I__10681\ : CascadeMux
    port map (
            O => \N__42880\,
            I => \N__42877\
        );

    \I__10680\ : InMux
    port map (
            O => \N__42877\,
            I => \N__42874\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__42874\,
            I => \N__42871\
        );

    \I__10678\ : Span4Mux_h
    port map (
            O => \N__42871\,
            I => \N__42866\
        );

    \I__10677\ : CascadeMux
    port map (
            O => \N__42870\,
            I => \N__42863\
        );

    \I__10676\ : InMux
    port map (
            O => \N__42869\,
            I => \N__42860\
        );

    \I__10675\ : Span4Mux_v
    port map (
            O => \N__42866\,
            I => \N__42856\
        );

    \I__10674\ : InMux
    port map (
            O => \N__42863\,
            I => \N__42853\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__42860\,
            I => \N__42850\
        );

    \I__10672\ : InMux
    port map (
            O => \N__42859\,
            I => \N__42847\
        );

    \I__10671\ : Span4Mux_v
    port map (
            O => \N__42856\,
            I => \N__42844\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__42853\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__10669\ : Odrv4
    port map (
            O => \N__42850\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__10668\ : LocalMux
    port map (
            O => \N__42847\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__10667\ : Odrv4
    port map (
            O => \N__42844\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__10666\ : InMux
    port map (
            O => \N__42835\,
            I => \N__42831\
        );

    \I__10665\ : InMux
    port map (
            O => \N__42834\,
            I => \N__42825\
        );

    \I__10664\ : LocalMux
    port map (
            O => \N__42831\,
            I => \N__42822\
        );

    \I__10663\ : InMux
    port map (
            O => \N__42830\,
            I => \N__42817\
        );

    \I__10662\ : InMux
    port map (
            O => \N__42829\,
            I => \N__42817\
        );

    \I__10661\ : InMux
    port map (
            O => \N__42828\,
            I => \N__42814\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__42825\,
            I => \N__42807\
        );

    \I__10659\ : Span4Mux_v
    port map (
            O => \N__42822\,
            I => \N__42807\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__42817\,
            I => \N__42807\
        );

    \I__10657\ : LocalMux
    port map (
            O => \N__42814\,
            I => \N__42804\
        );

    \I__10656\ : Span4Mux_h
    port map (
            O => \N__42807\,
            I => \N__42801\
        );

    \I__10655\ : Odrv12
    port map (
            O => \N__42804\,
            I => \N_801_0\
        );

    \I__10654\ : Odrv4
    port map (
            O => \N__42801\,
            I => \N_801_0\
        );

    \I__10653\ : InMux
    port map (
            O => \N__42796\,
            I => \N__42793\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__42793\,
            I => \N__42788\
        );

    \I__10651\ : InMux
    port map (
            O => \N__42792\,
            I => \N__42785\
        );

    \I__10650\ : InMux
    port map (
            O => \N__42791\,
            I => \N__42782\
        );

    \I__10649\ : Span4Mux_h
    port map (
            O => \N__42788\,
            I => \N__42775\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__42785\,
            I => \N__42775\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__42782\,
            I => \N__42775\
        );

    \I__10646\ : Span4Mux_v
    port map (
            O => \N__42775\,
            I => \N__42769\
        );

    \I__10645\ : InMux
    port map (
            O => \N__42774\,
            I => \N__42766\
        );

    \I__10644\ : InMux
    port map (
            O => \N__42773\,
            I => \N__42761\
        );

    \I__10643\ : InMux
    port map (
            O => \N__42772\,
            I => \N__42758\
        );

    \I__10642\ : Span4Mux_h
    port map (
            O => \N__42769\,
            I => \N__42754\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__42766\,
            I => \N__42751\
        );

    \I__10640\ : InMux
    port map (
            O => \N__42765\,
            I => \N__42747\
        );

    \I__10639\ : InMux
    port map (
            O => \N__42764\,
            I => \N__42744\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__42761\,
            I => \N__42741\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__42758\,
            I => \N__42738\
        );

    \I__10636\ : CascadeMux
    port map (
            O => \N__42757\,
            I => \N__42735\
        );

    \I__10635\ : Span4Mux_h
    port map (
            O => \N__42754\,
            I => \N__42732\
        );

    \I__10634\ : Span4Mux_v
    port map (
            O => \N__42751\,
            I => \N__42729\
        );

    \I__10633\ : InMux
    port map (
            O => \N__42750\,
            I => \N__42726\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__42747\,
            I => \N__42723\
        );

    \I__10631\ : LocalMux
    port map (
            O => \N__42744\,
            I => \N__42720\
        );

    \I__10630\ : Span4Mux_v
    port map (
            O => \N__42741\,
            I => \N__42717\
        );

    \I__10629\ : Span4Mux_v
    port map (
            O => \N__42738\,
            I => \N__42714\
        );

    \I__10628\ : InMux
    port map (
            O => \N__42735\,
            I => \N__42711\
        );

    \I__10627\ : Span4Mux_h
    port map (
            O => \N__42732\,
            I => \N__42703\
        );

    \I__10626\ : Span4Mux_v
    port map (
            O => \N__42729\,
            I => \N__42703\
        );

    \I__10625\ : LocalMux
    port map (
            O => \N__42726\,
            I => \N__42703\
        );

    \I__10624\ : Span12Mux_v
    port map (
            O => \N__42723\,
            I => \N__42698\
        );

    \I__10623\ : Span12Mux_h
    port map (
            O => \N__42720\,
            I => \N__42698\
        );

    \I__10622\ : IoSpan4Mux
    port map (
            O => \N__42717\,
            I => \N__42695\
        );

    \I__10621\ : Sp12to4
    port map (
            O => \N__42714\,
            I => \N__42692\
        );

    \I__10620\ : LocalMux
    port map (
            O => \N__42711\,
            I => \N__42689\
        );

    \I__10619\ : InMux
    port map (
            O => \N__42710\,
            I => \N__42686\
        );

    \I__10618\ : Span4Mux_h
    port map (
            O => \N__42703\,
            I => \N__42683\
        );

    \I__10617\ : Span12Mux_h
    port map (
            O => \N__42698\,
            I => \N__42680\
        );

    \I__10616\ : IoSpan4Mux
    port map (
            O => \N__42695\,
            I => \N__42677\
        );

    \I__10615\ : Span12Mux_h
    port map (
            O => \N__42692\,
            I => \N__42670\
        );

    \I__10614\ : Sp12to4
    port map (
            O => \N__42689\,
            I => \N__42670\
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__42686\,
            I => \N__42670\
        );

    \I__10612\ : Span4Mux_v
    port map (
            O => \N__42683\,
            I => \N__42667\
        );

    \I__10611\ : Odrv12
    port map (
            O => \N__42680\,
            I => port_data_in_2
        );

    \I__10610\ : Odrv4
    port map (
            O => \N__42677\,
            I => port_data_in_2
        );

    \I__10609\ : Odrv12
    port map (
            O => \N__42670\,
            I => port_data_in_2
        );

    \I__10608\ : Odrv4
    port map (
            O => \N__42667\,
            I => port_data_in_2
        );

    \I__10607\ : CascadeMux
    port map (
            O => \N__42658\,
            I => \N_1075_cascade_\
        );

    \I__10606\ : InMux
    port map (
            O => \N__42655\,
            I => \N__42652\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__42652\,
            I => \M_this_map_address_qc_1_0\
        );

    \I__10604\ : InMux
    port map (
            O => \N__42649\,
            I => \N__42645\
        );

    \I__10603\ : InMux
    port map (
            O => \N__42648\,
            I => \N__42642\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__42645\,
            I => \N__42637\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__42642\,
            I => \N__42637\
        );

    \I__10600\ : Span4Mux_v
    port map (
            O => \N__42637\,
            I => \N__42633\
        );

    \I__10599\ : InMux
    port map (
            O => \N__42636\,
            I => \N__42630\
        );

    \I__10598\ : Span4Mux_h
    port map (
            O => \N__42633\,
            I => \N__42625\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__42630\,
            I => \N__42625\
        );

    \I__10596\ : Span4Mux_h
    port map (
            O => \N__42625\,
            I => \N__42622\
        );

    \I__10595\ : Span4Mux_v
    port map (
            O => \N__42622\,
            I => \N__42619\
        );

    \I__10594\ : Odrv4
    port map (
            O => \N__42619\,
            I => port_address_in_3
        );

    \I__10593\ : InMux
    port map (
            O => \N__42616\,
            I => \N__42611\
        );

    \I__10592\ : InMux
    port map (
            O => \N__42615\,
            I => \N__42608\
        );

    \I__10591\ : InMux
    port map (
            O => \N__42614\,
            I => \N__42605\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__42611\,
            I => \N__42598\
        );

    \I__10589\ : LocalMux
    port map (
            O => \N__42608\,
            I => \N__42598\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__42605\,
            I => \N__42598\
        );

    \I__10587\ : Odrv12
    port map (
            O => \N__42598\,
            I => \N_459_0\
        );

    \I__10586\ : InMux
    port map (
            O => \N__42595\,
            I => \N__42589\
        );

    \I__10585\ : InMux
    port map (
            O => \N__42594\,
            I => \N__42585\
        );

    \I__10584\ : InMux
    port map (
            O => \N__42593\,
            I => \N__42582\
        );

    \I__10583\ : InMux
    port map (
            O => \N__42592\,
            I => \N__42579\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__42589\,
            I => \N__42576\
        );

    \I__10581\ : InMux
    port map (
            O => \N__42588\,
            I => \N__42573\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__42585\,
            I => \N__42568\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__42582\,
            I => \N__42568\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__42579\,
            I => \N__42565\
        );

    \I__10577\ : Span4Mux_h
    port map (
            O => \N__42576\,
            I => \N__42562\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__42573\,
            I => \N__42555\
        );

    \I__10575\ : Span4Mux_v
    port map (
            O => \N__42568\,
            I => \N__42555\
        );

    \I__10574\ : Span4Mux_h
    port map (
            O => \N__42565\,
            I => \N__42555\
        );

    \I__10573\ : Span4Mux_h
    port map (
            O => \N__42562\,
            I => \N__42552\
        );

    \I__10572\ : Span4Mux_h
    port map (
            O => \N__42555\,
            I => \N__42549\
        );

    \I__10571\ : Odrv4
    port map (
            O => \N__42552\,
            I => \N_1276\
        );

    \I__10570\ : Odrv4
    port map (
            O => \N__42549\,
            I => \N_1276\
        );

    \I__10569\ : InMux
    port map (
            O => \N__42544\,
            I => \N__42536\
        );

    \I__10568\ : InMux
    port map (
            O => \N__42543\,
            I => \N__42533\
        );

    \I__10567\ : CascadeMux
    port map (
            O => \N__42542\,
            I => \N__42530\
        );

    \I__10566\ : InMux
    port map (
            O => \N__42541\,
            I => \N__42526\
        );

    \I__10565\ : InMux
    port map (
            O => \N__42540\,
            I => \N__42523\
        );

    \I__10564\ : InMux
    port map (
            O => \N__42539\,
            I => \N__42520\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__42536\,
            I => \N__42517\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__42533\,
            I => \N__42514\
        );

    \I__10561\ : InMux
    port map (
            O => \N__42530\,
            I => \N__42509\
        );

    \I__10560\ : InMux
    port map (
            O => \N__42529\,
            I => \N__42509\
        );

    \I__10559\ : LocalMux
    port map (
            O => \N__42526\,
            I => \N__42500\
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__42523\,
            I => \N__42500\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__42520\,
            I => \N__42500\
        );

    \I__10556\ : Span12Mux_v
    port map (
            O => \N__42517\,
            I => \N__42496\
        );

    \I__10555\ : Span4Mux_v
    port map (
            O => \N__42514\,
            I => \N__42493\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__42509\,
            I => \N__42490\
        );

    \I__10553\ : InMux
    port map (
            O => \N__42508\,
            I => \N__42487\
        );

    \I__10552\ : InMux
    port map (
            O => \N__42507\,
            I => \N__42484\
        );

    \I__10551\ : Span12Mux_s10_h
    port map (
            O => \N__42500\,
            I => \N__42481\
        );

    \I__10550\ : InMux
    port map (
            O => \N__42499\,
            I => \N__42478\
        );

    \I__10549\ : Odrv12
    port map (
            O => \N__42496\,
            I => \N_1242\
        );

    \I__10548\ : Odrv4
    port map (
            O => \N__42493\,
            I => \N_1242\
        );

    \I__10547\ : Odrv4
    port map (
            O => \N__42490\,
            I => \N_1242\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__42487\,
            I => \N_1242\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__42484\,
            I => \N_1242\
        );

    \I__10544\ : Odrv12
    port map (
            O => \N__42481\,
            I => \N_1242\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__42478\,
            I => \N_1242\
        );

    \I__10542\ : CascadeMux
    port map (
            O => \N__42463\,
            I => \N__42460\
        );

    \I__10541\ : InMux
    port map (
            O => \N__42460\,
            I => \N__42456\
        );

    \I__10540\ : CascadeMux
    port map (
            O => \N__42459\,
            I => \N__42453\
        );

    \I__10539\ : LocalMux
    port map (
            O => \N__42456\,
            I => \N__42450\
        );

    \I__10538\ : InMux
    port map (
            O => \N__42453\,
            I => \N__42446\
        );

    \I__10537\ : Span4Mux_h
    port map (
            O => \N__42450\,
            I => \N__42440\
        );

    \I__10536\ : InMux
    port map (
            O => \N__42449\,
            I => \N__42436\
        );

    \I__10535\ : LocalMux
    port map (
            O => \N__42446\,
            I => \N__42433\
        );

    \I__10534\ : InMux
    port map (
            O => \N__42445\,
            I => \N__42430\
        );

    \I__10533\ : InMux
    port map (
            O => \N__42444\,
            I => \N__42426\
        );

    \I__10532\ : InMux
    port map (
            O => \N__42443\,
            I => \N__42423\
        );

    \I__10531\ : Span4Mux_h
    port map (
            O => \N__42440\,
            I => \N__42420\
        );

    \I__10530\ : InMux
    port map (
            O => \N__42439\,
            I => \N__42417\
        );

    \I__10529\ : LocalMux
    port map (
            O => \N__42436\,
            I => \N__42412\
        );

    \I__10528\ : Span4Mux_h
    port map (
            O => \N__42433\,
            I => \N__42407\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__42430\,
            I => \N__42407\
        );

    \I__10526\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42404\
        );

    \I__10525\ : LocalMux
    port map (
            O => \N__42426\,
            I => \N__42401\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__42423\,
            I => \N__42398\
        );

    \I__10523\ : Span4Mux_h
    port map (
            O => \N__42420\,
            I => \N__42393\
        );

    \I__10522\ : LocalMux
    port map (
            O => \N__42417\,
            I => \N__42393\
        );

    \I__10521\ : InMux
    port map (
            O => \N__42416\,
            I => \N__42390\
        );

    \I__10520\ : InMux
    port map (
            O => \N__42415\,
            I => \N__42387\
        );

    \I__10519\ : Span4Mux_v
    port map (
            O => \N__42412\,
            I => \N__42384\
        );

    \I__10518\ : Span4Mux_h
    port map (
            O => \N__42407\,
            I => \N__42381\
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__42404\,
            I => \N__42378\
        );

    \I__10516\ : Span4Mux_h
    port map (
            O => \N__42401\,
            I => \N__42374\
        );

    \I__10515\ : Span4Mux_v
    port map (
            O => \N__42398\,
            I => \N__42371\
        );

    \I__10514\ : Span4Mux_h
    port map (
            O => \N__42393\,
            I => \N__42368\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__42390\,
            I => \N__42363\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__42387\,
            I => \N__42363\
        );

    \I__10511\ : Span4Mux_v
    port map (
            O => \N__42384\,
            I => \N__42358\
        );

    \I__10510\ : Span4Mux_h
    port map (
            O => \N__42381\,
            I => \N__42358\
        );

    \I__10509\ : Span4Mux_v
    port map (
            O => \N__42378\,
            I => \N__42355\
        );

    \I__10508\ : InMux
    port map (
            O => \N__42377\,
            I => \N__42352\
        );

    \I__10507\ : Span4Mux_v
    port map (
            O => \N__42374\,
            I => \N__42347\
        );

    \I__10506\ : Span4Mux_h
    port map (
            O => \N__42371\,
            I => \N__42347\
        );

    \I__10505\ : Span4Mux_v
    port map (
            O => \N__42368\,
            I => \N__42342\
        );

    \I__10504\ : Span4Mux_h
    port map (
            O => \N__42363\,
            I => \N__42342\
        );

    \I__10503\ : Span4Mux_h
    port map (
            O => \N__42358\,
            I => \N__42339\
        );

    \I__10502\ : Sp12to4
    port map (
            O => \N__42355\,
            I => \N__42334\
        );

    \I__10501\ : LocalMux
    port map (
            O => \N__42352\,
            I => \N__42334\
        );

    \I__10500\ : Span4Mux_h
    port map (
            O => \N__42347\,
            I => \N__42329\
        );

    \I__10499\ : Span4Mux_v
    port map (
            O => \N__42342\,
            I => \N__42329\
        );

    \I__10498\ : Sp12to4
    port map (
            O => \N__42339\,
            I => \N__42324\
        );

    \I__10497\ : Span12Mux_h
    port map (
            O => \N__42334\,
            I => \N__42324\
        );

    \I__10496\ : Odrv4
    port map (
            O => \N__42329\,
            I => port_data_in_0
        );

    \I__10495\ : Odrv12
    port map (
            O => \N__42324\,
            I => port_data_in_0
        );

    \I__10494\ : InMux
    port map (
            O => \N__42319\,
            I => \N__42316\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__42316\,
            I => \N_1068\
        );

    \I__10492\ : InMux
    port map (
            O => \N__42313\,
            I => \N__42310\
        );

    \I__10491\ : LocalMux
    port map (
            O => \N__42310\,
            I => \M_this_map_address_qc_7_1\
        );

    \I__10490\ : InMux
    port map (
            O => \N__42307\,
            I => \N__42304\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__42304\,
            I => \N__42301\
        );

    \I__10488\ : Span4Mux_h
    port map (
            O => \N__42301\,
            I => \N__42298\
        );

    \I__10487\ : Odrv4
    port map (
            O => \N__42298\,
            I => \M_this_map_address_q_RNO_1Z0Z_5\
        );

    \I__10486\ : CascadeMux
    port map (
            O => \N__42295\,
            I => \N__42290\
        );

    \I__10485\ : InMux
    port map (
            O => \N__42294\,
            I => \N__42285\
        );

    \I__10484\ : InMux
    port map (
            O => \N__42293\,
            I => \N__42280\
        );

    \I__10483\ : InMux
    port map (
            O => \N__42290\,
            I => \N__42277\
        );

    \I__10482\ : InMux
    port map (
            O => \N__42289\,
            I => \N__42274\
        );

    \I__10481\ : InMux
    port map (
            O => \N__42288\,
            I => \N__42271\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__42285\,
            I => \N__42268\
        );

    \I__10479\ : InMux
    port map (
            O => \N__42284\,
            I => \N__42263\
        );

    \I__10478\ : InMux
    port map (
            O => \N__42283\,
            I => \N__42263\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__42280\,
            I => \N__42255\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__42277\,
            I => \N__42250\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__42274\,
            I => \N__42250\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__42271\,
            I => \N__42247\
        );

    \I__10473\ : Span4Mux_v
    port map (
            O => \N__42268\,
            I => \N__42244\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__42263\,
            I => \N__42241\
        );

    \I__10471\ : InMux
    port map (
            O => \N__42262\,
            I => \N__42237\
        );

    \I__10470\ : CascadeMux
    port map (
            O => \N__42261\,
            I => \N__42234\
        );

    \I__10469\ : InMux
    port map (
            O => \N__42260\,
            I => \N__42227\
        );

    \I__10468\ : InMux
    port map (
            O => \N__42259\,
            I => \N__42227\
        );

    \I__10467\ : InMux
    port map (
            O => \N__42258\,
            I => \N__42227\
        );

    \I__10466\ : Span4Mux_h
    port map (
            O => \N__42255\,
            I => \N__42220\
        );

    \I__10465\ : Span4Mux_v
    port map (
            O => \N__42250\,
            I => \N__42220\
        );

    \I__10464\ : Span4Mux_v
    port map (
            O => \N__42247\,
            I => \N__42220\
        );

    \I__10463\ : Span4Mux_h
    port map (
            O => \N__42244\,
            I => \N__42217\
        );

    \I__10462\ : Span4Mux_h
    port map (
            O => \N__42241\,
            I => \N__42214\
        );

    \I__10461\ : InMux
    port map (
            O => \N__42240\,
            I => \N__42211\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__42237\,
            I => \N__42208\
        );

    \I__10459\ : InMux
    port map (
            O => \N__42234\,
            I => \N__42205\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__42227\,
            I => \N_1258\
        );

    \I__10457\ : Odrv4
    port map (
            O => \N__42220\,
            I => \N_1258\
        );

    \I__10456\ : Odrv4
    port map (
            O => \N__42217\,
            I => \N_1258\
        );

    \I__10455\ : Odrv4
    port map (
            O => \N__42214\,
            I => \N_1258\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__42211\,
            I => \N_1258\
        );

    \I__10453\ : Odrv12
    port map (
            O => \N__42208\,
            I => \N_1258\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__42205\,
            I => \N_1258\
        );

    \I__10451\ : CascadeMux
    port map (
            O => \N__42190\,
            I => \N__42187\
        );

    \I__10450\ : CascadeBuf
    port map (
            O => \N__42187\,
            I => \N__42184\
        );

    \I__10449\ : CascadeMux
    port map (
            O => \N__42184\,
            I => \N__42180\
        );

    \I__10448\ : CascadeMux
    port map (
            O => \N__42183\,
            I => \N__42177\
        );

    \I__10447\ : InMux
    port map (
            O => \N__42180\,
            I => \N__42174\
        );

    \I__10446\ : InMux
    port map (
            O => \N__42177\,
            I => \N__42171\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__42174\,
            I => \N__42168\
        );

    \I__10444\ : LocalMux
    port map (
            O => \N__42171\,
            I => \N__42164\
        );

    \I__10443\ : Span4Mux_s2_v
    port map (
            O => \N__42168\,
            I => \N__42161\
        );

    \I__10442\ : InMux
    port map (
            O => \N__42167\,
            I => \N__42158\
        );

    \I__10441\ : Span4Mux_h
    port map (
            O => \N__42164\,
            I => \N__42155\
        );

    \I__10440\ : Span4Mux_v
    port map (
            O => \N__42161\,
            I => \N__42152\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__42158\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__10438\ : Odrv4
    port map (
            O => \N__42155\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__10437\ : Odrv4
    port map (
            O => \N__42152\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__10436\ : ClkMux
    port map (
            O => \N__42145\,
            I => \N__41659\
        );

    \I__10435\ : ClkMux
    port map (
            O => \N__42144\,
            I => \N__41659\
        );

    \I__10434\ : ClkMux
    port map (
            O => \N__42143\,
            I => \N__41659\
        );

    \I__10433\ : ClkMux
    port map (
            O => \N__42142\,
            I => \N__41659\
        );

    \I__10432\ : ClkMux
    port map (
            O => \N__42141\,
            I => \N__41659\
        );

    \I__10431\ : ClkMux
    port map (
            O => \N__42140\,
            I => \N__41659\
        );

    \I__10430\ : ClkMux
    port map (
            O => \N__42139\,
            I => \N__41659\
        );

    \I__10429\ : ClkMux
    port map (
            O => \N__42138\,
            I => \N__41659\
        );

    \I__10428\ : ClkMux
    port map (
            O => \N__42137\,
            I => \N__41659\
        );

    \I__10427\ : ClkMux
    port map (
            O => \N__42136\,
            I => \N__41659\
        );

    \I__10426\ : ClkMux
    port map (
            O => \N__42135\,
            I => \N__41659\
        );

    \I__10425\ : ClkMux
    port map (
            O => \N__42134\,
            I => \N__41659\
        );

    \I__10424\ : ClkMux
    port map (
            O => \N__42133\,
            I => \N__41659\
        );

    \I__10423\ : ClkMux
    port map (
            O => \N__42132\,
            I => \N__41659\
        );

    \I__10422\ : ClkMux
    port map (
            O => \N__42131\,
            I => \N__41659\
        );

    \I__10421\ : ClkMux
    port map (
            O => \N__42130\,
            I => \N__41659\
        );

    \I__10420\ : ClkMux
    port map (
            O => \N__42129\,
            I => \N__41659\
        );

    \I__10419\ : ClkMux
    port map (
            O => \N__42128\,
            I => \N__41659\
        );

    \I__10418\ : ClkMux
    port map (
            O => \N__42127\,
            I => \N__41659\
        );

    \I__10417\ : ClkMux
    port map (
            O => \N__42126\,
            I => \N__41659\
        );

    \I__10416\ : ClkMux
    port map (
            O => \N__42125\,
            I => \N__41659\
        );

    \I__10415\ : ClkMux
    port map (
            O => \N__42124\,
            I => \N__41659\
        );

    \I__10414\ : ClkMux
    port map (
            O => \N__42123\,
            I => \N__41659\
        );

    \I__10413\ : ClkMux
    port map (
            O => \N__42122\,
            I => \N__41659\
        );

    \I__10412\ : ClkMux
    port map (
            O => \N__42121\,
            I => \N__41659\
        );

    \I__10411\ : ClkMux
    port map (
            O => \N__42120\,
            I => \N__41659\
        );

    \I__10410\ : ClkMux
    port map (
            O => \N__42119\,
            I => \N__41659\
        );

    \I__10409\ : ClkMux
    port map (
            O => \N__42118\,
            I => \N__41659\
        );

    \I__10408\ : ClkMux
    port map (
            O => \N__42117\,
            I => \N__41659\
        );

    \I__10407\ : ClkMux
    port map (
            O => \N__42116\,
            I => \N__41659\
        );

    \I__10406\ : ClkMux
    port map (
            O => \N__42115\,
            I => \N__41659\
        );

    \I__10405\ : ClkMux
    port map (
            O => \N__42114\,
            I => \N__41659\
        );

    \I__10404\ : ClkMux
    port map (
            O => \N__42113\,
            I => \N__41659\
        );

    \I__10403\ : ClkMux
    port map (
            O => \N__42112\,
            I => \N__41659\
        );

    \I__10402\ : ClkMux
    port map (
            O => \N__42111\,
            I => \N__41659\
        );

    \I__10401\ : ClkMux
    port map (
            O => \N__42110\,
            I => \N__41659\
        );

    \I__10400\ : ClkMux
    port map (
            O => \N__42109\,
            I => \N__41659\
        );

    \I__10399\ : ClkMux
    port map (
            O => \N__42108\,
            I => \N__41659\
        );

    \I__10398\ : ClkMux
    port map (
            O => \N__42107\,
            I => \N__41659\
        );

    \I__10397\ : ClkMux
    port map (
            O => \N__42106\,
            I => \N__41659\
        );

    \I__10396\ : ClkMux
    port map (
            O => \N__42105\,
            I => \N__41659\
        );

    \I__10395\ : ClkMux
    port map (
            O => \N__42104\,
            I => \N__41659\
        );

    \I__10394\ : ClkMux
    port map (
            O => \N__42103\,
            I => \N__41659\
        );

    \I__10393\ : ClkMux
    port map (
            O => \N__42102\,
            I => \N__41659\
        );

    \I__10392\ : ClkMux
    port map (
            O => \N__42101\,
            I => \N__41659\
        );

    \I__10391\ : ClkMux
    port map (
            O => \N__42100\,
            I => \N__41659\
        );

    \I__10390\ : ClkMux
    port map (
            O => \N__42099\,
            I => \N__41659\
        );

    \I__10389\ : ClkMux
    port map (
            O => \N__42098\,
            I => \N__41659\
        );

    \I__10388\ : ClkMux
    port map (
            O => \N__42097\,
            I => \N__41659\
        );

    \I__10387\ : ClkMux
    port map (
            O => \N__42096\,
            I => \N__41659\
        );

    \I__10386\ : ClkMux
    port map (
            O => \N__42095\,
            I => \N__41659\
        );

    \I__10385\ : ClkMux
    port map (
            O => \N__42094\,
            I => \N__41659\
        );

    \I__10384\ : ClkMux
    port map (
            O => \N__42093\,
            I => \N__41659\
        );

    \I__10383\ : ClkMux
    port map (
            O => \N__42092\,
            I => \N__41659\
        );

    \I__10382\ : ClkMux
    port map (
            O => \N__42091\,
            I => \N__41659\
        );

    \I__10381\ : ClkMux
    port map (
            O => \N__42090\,
            I => \N__41659\
        );

    \I__10380\ : ClkMux
    port map (
            O => \N__42089\,
            I => \N__41659\
        );

    \I__10379\ : ClkMux
    port map (
            O => \N__42088\,
            I => \N__41659\
        );

    \I__10378\ : ClkMux
    port map (
            O => \N__42087\,
            I => \N__41659\
        );

    \I__10377\ : ClkMux
    port map (
            O => \N__42086\,
            I => \N__41659\
        );

    \I__10376\ : ClkMux
    port map (
            O => \N__42085\,
            I => \N__41659\
        );

    \I__10375\ : ClkMux
    port map (
            O => \N__42084\,
            I => \N__41659\
        );

    \I__10374\ : ClkMux
    port map (
            O => \N__42083\,
            I => \N__41659\
        );

    \I__10373\ : ClkMux
    port map (
            O => \N__42082\,
            I => \N__41659\
        );

    \I__10372\ : ClkMux
    port map (
            O => \N__42081\,
            I => \N__41659\
        );

    \I__10371\ : ClkMux
    port map (
            O => \N__42080\,
            I => \N__41659\
        );

    \I__10370\ : ClkMux
    port map (
            O => \N__42079\,
            I => \N__41659\
        );

    \I__10369\ : ClkMux
    port map (
            O => \N__42078\,
            I => \N__41659\
        );

    \I__10368\ : ClkMux
    port map (
            O => \N__42077\,
            I => \N__41659\
        );

    \I__10367\ : ClkMux
    port map (
            O => \N__42076\,
            I => \N__41659\
        );

    \I__10366\ : ClkMux
    port map (
            O => \N__42075\,
            I => \N__41659\
        );

    \I__10365\ : ClkMux
    port map (
            O => \N__42074\,
            I => \N__41659\
        );

    \I__10364\ : ClkMux
    port map (
            O => \N__42073\,
            I => \N__41659\
        );

    \I__10363\ : ClkMux
    port map (
            O => \N__42072\,
            I => \N__41659\
        );

    \I__10362\ : ClkMux
    port map (
            O => \N__42071\,
            I => \N__41659\
        );

    \I__10361\ : ClkMux
    port map (
            O => \N__42070\,
            I => \N__41659\
        );

    \I__10360\ : ClkMux
    port map (
            O => \N__42069\,
            I => \N__41659\
        );

    \I__10359\ : ClkMux
    port map (
            O => \N__42068\,
            I => \N__41659\
        );

    \I__10358\ : ClkMux
    port map (
            O => \N__42067\,
            I => \N__41659\
        );

    \I__10357\ : ClkMux
    port map (
            O => \N__42066\,
            I => \N__41659\
        );

    \I__10356\ : ClkMux
    port map (
            O => \N__42065\,
            I => \N__41659\
        );

    \I__10355\ : ClkMux
    port map (
            O => \N__42064\,
            I => \N__41659\
        );

    \I__10354\ : ClkMux
    port map (
            O => \N__42063\,
            I => \N__41659\
        );

    \I__10353\ : ClkMux
    port map (
            O => \N__42062\,
            I => \N__41659\
        );

    \I__10352\ : ClkMux
    port map (
            O => \N__42061\,
            I => \N__41659\
        );

    \I__10351\ : ClkMux
    port map (
            O => \N__42060\,
            I => \N__41659\
        );

    \I__10350\ : ClkMux
    port map (
            O => \N__42059\,
            I => \N__41659\
        );

    \I__10349\ : ClkMux
    port map (
            O => \N__42058\,
            I => \N__41659\
        );

    \I__10348\ : ClkMux
    port map (
            O => \N__42057\,
            I => \N__41659\
        );

    \I__10347\ : ClkMux
    port map (
            O => \N__42056\,
            I => \N__41659\
        );

    \I__10346\ : ClkMux
    port map (
            O => \N__42055\,
            I => \N__41659\
        );

    \I__10345\ : ClkMux
    port map (
            O => \N__42054\,
            I => \N__41659\
        );

    \I__10344\ : ClkMux
    port map (
            O => \N__42053\,
            I => \N__41659\
        );

    \I__10343\ : ClkMux
    port map (
            O => \N__42052\,
            I => \N__41659\
        );

    \I__10342\ : ClkMux
    port map (
            O => \N__42051\,
            I => \N__41659\
        );

    \I__10341\ : ClkMux
    port map (
            O => \N__42050\,
            I => \N__41659\
        );

    \I__10340\ : ClkMux
    port map (
            O => \N__42049\,
            I => \N__41659\
        );

    \I__10339\ : ClkMux
    port map (
            O => \N__42048\,
            I => \N__41659\
        );

    \I__10338\ : ClkMux
    port map (
            O => \N__42047\,
            I => \N__41659\
        );

    \I__10337\ : ClkMux
    port map (
            O => \N__42046\,
            I => \N__41659\
        );

    \I__10336\ : ClkMux
    port map (
            O => \N__42045\,
            I => \N__41659\
        );

    \I__10335\ : ClkMux
    port map (
            O => \N__42044\,
            I => \N__41659\
        );

    \I__10334\ : ClkMux
    port map (
            O => \N__42043\,
            I => \N__41659\
        );

    \I__10333\ : ClkMux
    port map (
            O => \N__42042\,
            I => \N__41659\
        );

    \I__10332\ : ClkMux
    port map (
            O => \N__42041\,
            I => \N__41659\
        );

    \I__10331\ : ClkMux
    port map (
            O => \N__42040\,
            I => \N__41659\
        );

    \I__10330\ : ClkMux
    port map (
            O => \N__42039\,
            I => \N__41659\
        );

    \I__10329\ : ClkMux
    port map (
            O => \N__42038\,
            I => \N__41659\
        );

    \I__10328\ : ClkMux
    port map (
            O => \N__42037\,
            I => \N__41659\
        );

    \I__10327\ : ClkMux
    port map (
            O => \N__42036\,
            I => \N__41659\
        );

    \I__10326\ : ClkMux
    port map (
            O => \N__42035\,
            I => \N__41659\
        );

    \I__10325\ : ClkMux
    port map (
            O => \N__42034\,
            I => \N__41659\
        );

    \I__10324\ : ClkMux
    port map (
            O => \N__42033\,
            I => \N__41659\
        );

    \I__10323\ : ClkMux
    port map (
            O => \N__42032\,
            I => \N__41659\
        );

    \I__10322\ : ClkMux
    port map (
            O => \N__42031\,
            I => \N__41659\
        );

    \I__10321\ : ClkMux
    port map (
            O => \N__42030\,
            I => \N__41659\
        );

    \I__10320\ : ClkMux
    port map (
            O => \N__42029\,
            I => \N__41659\
        );

    \I__10319\ : ClkMux
    port map (
            O => \N__42028\,
            I => \N__41659\
        );

    \I__10318\ : ClkMux
    port map (
            O => \N__42027\,
            I => \N__41659\
        );

    \I__10317\ : ClkMux
    port map (
            O => \N__42026\,
            I => \N__41659\
        );

    \I__10316\ : ClkMux
    port map (
            O => \N__42025\,
            I => \N__41659\
        );

    \I__10315\ : ClkMux
    port map (
            O => \N__42024\,
            I => \N__41659\
        );

    \I__10314\ : ClkMux
    port map (
            O => \N__42023\,
            I => \N__41659\
        );

    \I__10313\ : ClkMux
    port map (
            O => \N__42022\,
            I => \N__41659\
        );

    \I__10312\ : ClkMux
    port map (
            O => \N__42021\,
            I => \N__41659\
        );

    \I__10311\ : ClkMux
    port map (
            O => \N__42020\,
            I => \N__41659\
        );

    \I__10310\ : ClkMux
    port map (
            O => \N__42019\,
            I => \N__41659\
        );

    \I__10309\ : ClkMux
    port map (
            O => \N__42018\,
            I => \N__41659\
        );

    \I__10308\ : ClkMux
    port map (
            O => \N__42017\,
            I => \N__41659\
        );

    \I__10307\ : ClkMux
    port map (
            O => \N__42016\,
            I => \N__41659\
        );

    \I__10306\ : ClkMux
    port map (
            O => \N__42015\,
            I => \N__41659\
        );

    \I__10305\ : ClkMux
    port map (
            O => \N__42014\,
            I => \N__41659\
        );

    \I__10304\ : ClkMux
    port map (
            O => \N__42013\,
            I => \N__41659\
        );

    \I__10303\ : ClkMux
    port map (
            O => \N__42012\,
            I => \N__41659\
        );

    \I__10302\ : ClkMux
    port map (
            O => \N__42011\,
            I => \N__41659\
        );

    \I__10301\ : ClkMux
    port map (
            O => \N__42010\,
            I => \N__41659\
        );

    \I__10300\ : ClkMux
    port map (
            O => \N__42009\,
            I => \N__41659\
        );

    \I__10299\ : ClkMux
    port map (
            O => \N__42008\,
            I => \N__41659\
        );

    \I__10298\ : ClkMux
    port map (
            O => \N__42007\,
            I => \N__41659\
        );

    \I__10297\ : ClkMux
    port map (
            O => \N__42006\,
            I => \N__41659\
        );

    \I__10296\ : ClkMux
    port map (
            O => \N__42005\,
            I => \N__41659\
        );

    \I__10295\ : ClkMux
    port map (
            O => \N__42004\,
            I => \N__41659\
        );

    \I__10294\ : ClkMux
    port map (
            O => \N__42003\,
            I => \N__41659\
        );

    \I__10293\ : ClkMux
    port map (
            O => \N__42002\,
            I => \N__41659\
        );

    \I__10292\ : ClkMux
    port map (
            O => \N__42001\,
            I => \N__41659\
        );

    \I__10291\ : ClkMux
    port map (
            O => \N__42000\,
            I => \N__41659\
        );

    \I__10290\ : ClkMux
    port map (
            O => \N__41999\,
            I => \N__41659\
        );

    \I__10289\ : ClkMux
    port map (
            O => \N__41998\,
            I => \N__41659\
        );

    \I__10288\ : ClkMux
    port map (
            O => \N__41997\,
            I => \N__41659\
        );

    \I__10287\ : ClkMux
    port map (
            O => \N__41996\,
            I => \N__41659\
        );

    \I__10286\ : ClkMux
    port map (
            O => \N__41995\,
            I => \N__41659\
        );

    \I__10285\ : ClkMux
    port map (
            O => \N__41994\,
            I => \N__41659\
        );

    \I__10284\ : ClkMux
    port map (
            O => \N__41993\,
            I => \N__41659\
        );

    \I__10283\ : ClkMux
    port map (
            O => \N__41992\,
            I => \N__41659\
        );

    \I__10282\ : ClkMux
    port map (
            O => \N__41991\,
            I => \N__41659\
        );

    \I__10281\ : ClkMux
    port map (
            O => \N__41990\,
            I => \N__41659\
        );

    \I__10280\ : ClkMux
    port map (
            O => \N__41989\,
            I => \N__41659\
        );

    \I__10279\ : ClkMux
    port map (
            O => \N__41988\,
            I => \N__41659\
        );

    \I__10278\ : ClkMux
    port map (
            O => \N__41987\,
            I => \N__41659\
        );

    \I__10277\ : ClkMux
    port map (
            O => \N__41986\,
            I => \N__41659\
        );

    \I__10276\ : ClkMux
    port map (
            O => \N__41985\,
            I => \N__41659\
        );

    \I__10275\ : ClkMux
    port map (
            O => \N__41984\,
            I => \N__41659\
        );

    \I__10274\ : GlobalMux
    port map (
            O => \N__41659\,
            I => \N__41656\
        );

    \I__10273\ : gio2CtrlBuf
    port map (
            O => \N__41656\,
            I => clk_0_c_g
        );

    \I__10272\ : SRMux
    port map (
            O => \N__41653\,
            I => \N__41608\
        );

    \I__10271\ : SRMux
    port map (
            O => \N__41652\,
            I => \N__41608\
        );

    \I__10270\ : SRMux
    port map (
            O => \N__41651\,
            I => \N__41608\
        );

    \I__10269\ : SRMux
    port map (
            O => \N__41650\,
            I => \N__41608\
        );

    \I__10268\ : SRMux
    port map (
            O => \N__41649\,
            I => \N__41608\
        );

    \I__10267\ : SRMux
    port map (
            O => \N__41648\,
            I => \N__41608\
        );

    \I__10266\ : SRMux
    port map (
            O => \N__41647\,
            I => \N__41608\
        );

    \I__10265\ : SRMux
    port map (
            O => \N__41646\,
            I => \N__41608\
        );

    \I__10264\ : SRMux
    port map (
            O => \N__41645\,
            I => \N__41608\
        );

    \I__10263\ : SRMux
    port map (
            O => \N__41644\,
            I => \N__41608\
        );

    \I__10262\ : SRMux
    port map (
            O => \N__41643\,
            I => \N__41608\
        );

    \I__10261\ : SRMux
    port map (
            O => \N__41642\,
            I => \N__41608\
        );

    \I__10260\ : SRMux
    port map (
            O => \N__41641\,
            I => \N__41608\
        );

    \I__10259\ : SRMux
    port map (
            O => \N__41640\,
            I => \N__41608\
        );

    \I__10258\ : SRMux
    port map (
            O => \N__41639\,
            I => \N__41608\
        );

    \I__10257\ : GlobalMux
    port map (
            O => \N__41608\,
            I => \N__41605\
        );

    \I__10256\ : gio2CtrlBuf
    port map (
            O => \N__41605\,
            I => \N_620_g\
        );

    \I__10255\ : InMux
    port map (
            O => \N__41602\,
            I => \N__41598\
        );

    \I__10254\ : InMux
    port map (
            O => \N__41601\,
            I => \N__41595\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__41598\,
            I => \N__41592\
        );

    \I__10252\ : LocalMux
    port map (
            O => \N__41595\,
            I => \N__41589\
        );

    \I__10251\ : Span4Mux_v
    port map (
            O => \N__41592\,
            I => \N__41586\
        );

    \I__10250\ : Span12Mux_s9_h
    port map (
            O => \N__41589\,
            I => \N__41581\
        );

    \I__10249\ : Sp12to4
    port map (
            O => \N__41586\,
            I => \N__41581\
        );

    \I__10248\ : Span12Mux_v
    port map (
            O => \N__41581\,
            I => \N__41578\
        );

    \I__10247\ : Odrv12
    port map (
            O => \N__41578\,
            I => \M_this_map_ram_read_data_6\
        );

    \I__10246\ : IoInMux
    port map (
            O => \N__41575\,
            I => \N__41572\
        );

    \I__10245\ : LocalMux
    port map (
            O => \N__41572\,
            I => \N__41569\
        );

    \I__10244\ : Span4Mux_s3_h
    port map (
            O => \N__41569\,
            I => \N__41566\
        );

    \I__10243\ : Span4Mux_v
    port map (
            O => \N__41566\,
            I => \N__41563\
        );

    \I__10242\ : Odrv4
    port map (
            O => \N__41563\,
            I => \N_734_0\
        );

    \I__10241\ : CascadeMux
    port map (
            O => \N__41560\,
            I => \N__41557\
        );

    \I__10240\ : CascadeBuf
    port map (
            O => \N__41557\,
            I => \N__41554\
        );

    \I__10239\ : CascadeMux
    port map (
            O => \N__41554\,
            I => \N__41551\
        );

    \I__10238\ : InMux
    port map (
            O => \N__41551\,
            I => \N__41546\
        );

    \I__10237\ : CascadeMux
    port map (
            O => \N__41550\,
            I => \N__41543\
        );

    \I__10236\ : InMux
    port map (
            O => \N__41549\,
            I => \N__41539\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__41546\,
            I => \N__41536\
        );

    \I__10234\ : InMux
    port map (
            O => \N__41543\,
            I => \N__41533\
        );

    \I__10233\ : InMux
    port map (
            O => \N__41542\,
            I => \N__41530\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__41539\,
            I => \N__41527\
        );

    \I__10231\ : Span4Mux_v
    port map (
            O => \N__41536\,
            I => \N__41524\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__41533\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__10229\ : LocalMux
    port map (
            O => \N__41530\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__10228\ : Odrv4
    port map (
            O => \N__41527\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__10227\ : Odrv4
    port map (
            O => \N__41524\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__10226\ : InMux
    port map (
            O => \N__41515\,
            I => \N__41506\
        );

    \I__10225\ : InMux
    port map (
            O => \N__41514\,
            I => \N__41503\
        );

    \I__10224\ : InMux
    port map (
            O => \N__41513\,
            I => \N__41500\
        );

    \I__10223\ : InMux
    port map (
            O => \N__41512\,
            I => \N__41497\
        );

    \I__10222\ : InMux
    port map (
            O => \N__41511\,
            I => \N__41494\
        );

    \I__10221\ : InMux
    port map (
            O => \N__41510\,
            I => \N__41491\
        );

    \I__10220\ : InMux
    port map (
            O => \N__41509\,
            I => \N__41488\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__41506\,
            I => \N__41485\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__41503\,
            I => \N__41482\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__41500\,
            I => \N__41475\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__41497\,
            I => \N__41475\
        );

    \I__10215\ : LocalMux
    port map (
            O => \N__41494\,
            I => \N__41475\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__41491\,
            I => \N__41471\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__41488\,
            I => \N__41467\
        );

    \I__10212\ : Span4Mux_h
    port map (
            O => \N__41485\,
            I => \N__41461\
        );

    \I__10211\ : Span4Mux_v
    port map (
            O => \N__41482\,
            I => \N__41461\
        );

    \I__10210\ : Span4Mux_v
    port map (
            O => \N__41475\,
            I => \N__41458\
        );

    \I__10209\ : InMux
    port map (
            O => \N__41474\,
            I => \N__41455\
        );

    \I__10208\ : Span4Mux_h
    port map (
            O => \N__41471\,
            I => \N__41451\
        );

    \I__10207\ : InMux
    port map (
            O => \N__41470\,
            I => \N__41448\
        );

    \I__10206\ : Span4Mux_h
    port map (
            O => \N__41467\,
            I => \N__41445\
        );

    \I__10205\ : InMux
    port map (
            O => \N__41466\,
            I => \N__41442\
        );

    \I__10204\ : Span4Mux_v
    port map (
            O => \N__41461\,
            I => \N__41437\
        );

    \I__10203\ : Span4Mux_h
    port map (
            O => \N__41458\,
            I => \N__41437\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__41455\,
            I => \N__41434\
        );

    \I__10201\ : InMux
    port map (
            O => \N__41454\,
            I => \N__41431\
        );

    \I__10200\ : Span4Mux_v
    port map (
            O => \N__41451\,
            I => \N__41426\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__41448\,
            I => \N__41426\
        );

    \I__10198\ : Span4Mux_v
    port map (
            O => \N__41445\,
            I => \N__41421\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__41442\,
            I => \N__41421\
        );

    \I__10196\ : Sp12to4
    port map (
            O => \N__41437\,
            I => \N__41418\
        );

    \I__10195\ : Span12Mux_v
    port map (
            O => \N__41434\,
            I => \N__41413\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__41431\,
            I => \N__41413\
        );

    \I__10193\ : Span4Mux_h
    port map (
            O => \N__41426\,
            I => \N__41410\
        );

    \I__10192\ : Span4Mux_v
    port map (
            O => \N__41421\,
            I => \N__41407\
        );

    \I__10191\ : Span12Mux_h
    port map (
            O => \N__41418\,
            I => \N__41404\
        );

    \I__10190\ : Span12Mux_h
    port map (
            O => \N__41413\,
            I => \N__41401\
        );

    \I__10189\ : Span4Mux_v
    port map (
            O => \N__41410\,
            I => \N__41398\
        );

    \I__10188\ : Span4Mux_h
    port map (
            O => \N__41407\,
            I => \N__41395\
        );

    \I__10187\ : Odrv12
    port map (
            O => \N__41404\,
            I => port_data_in_3
        );

    \I__10186\ : Odrv12
    port map (
            O => \N__41401\,
            I => port_data_in_3
        );

    \I__10185\ : Odrv4
    port map (
            O => \N__41398\,
            I => port_data_in_3
        );

    \I__10184\ : Odrv4
    port map (
            O => \N__41395\,
            I => port_data_in_3
        );

    \I__10183\ : CascadeMux
    port map (
            O => \N__41386\,
            I => \N_1078_cascade_\
        );

    \I__10182\ : InMux
    port map (
            O => \N__41383\,
            I => \N__41380\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__41380\,
            I => \N__41377\
        );

    \I__10180\ : Odrv4
    port map (
            O => \N__41377\,
            I => \M_this_map_address_qc_0_1\
        );

    \I__10179\ : InMux
    port map (
            O => \N__41374\,
            I => \N__41371\
        );

    \I__10178\ : LocalMux
    port map (
            O => \N__41371\,
            I => \N__41368\
        );

    \I__10177\ : Span4Mux_v
    port map (
            O => \N__41368\,
            I => \N__41365\
        );

    \I__10176\ : Span4Mux_v
    port map (
            O => \N__41365\,
            I => \N__41361\
        );

    \I__10175\ : InMux
    port map (
            O => \N__41364\,
            I => \N__41358\
        );

    \I__10174\ : Sp12to4
    port map (
            O => \N__41361\,
            I => \N__41355\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__41358\,
            I => \M_this_map_ram_read_data_2\
        );

    \I__10172\ : Odrv12
    port map (
            O => \N__41355\,
            I => \M_this_map_ram_read_data_2\
        );

    \I__10171\ : IoInMux
    port map (
            O => \N__41350\,
            I => \N__41347\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__41347\,
            I => \N__41344\
        );

    \I__10169\ : Odrv4
    port map (
            O => \N__41344\,
            I => \N_726_0\
        );

    \I__10168\ : InMux
    port map (
            O => \N__41341\,
            I => \N__41338\
        );

    \I__10167\ : LocalMux
    port map (
            O => \N__41338\,
            I => \un1_M_this_ext_address_q_cry_7_c_RNIQ14FZ0\
        );

    \I__10166\ : IoInMux
    port map (
            O => \N__41335\,
            I => \N__41332\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__41332\,
            I => \N__41329\
        );

    \I__10164\ : Span4Mux_s2_v
    port map (
            O => \N__41329\,
            I => \N__41326\
        );

    \I__10163\ : Sp12to4
    port map (
            O => \N__41326\,
            I => \N__41323\
        );

    \I__10162\ : Span12Mux_h
    port map (
            O => \N__41323\,
            I => \N__41319\
        );

    \I__10161\ : InMux
    port map (
            O => \N__41322\,
            I => \N__41316\
        );

    \I__10160\ : Odrv12
    port map (
            O => \N__41319\,
            I => \M_this_ext_address_qZ0Z_8\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__41316\,
            I => \M_this_ext_address_qZ0Z_8\
        );

    \I__10158\ : InMux
    port map (
            O => \N__41311\,
            I => \N__41308\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__41308\,
            I => \un1_M_this_ext_address_q_cry_0_THRU_CO\
        );

    \I__10156\ : IoInMux
    port map (
            O => \N__41305\,
            I => \N__41302\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__41302\,
            I => \N__41299\
        );

    \I__10154\ : Span4Mux_s2_v
    port map (
            O => \N__41299\,
            I => \N__41296\
        );

    \I__10153\ : Span4Mux_v
    port map (
            O => \N__41296\,
            I => \N__41292\
        );

    \I__10152\ : CascadeMux
    port map (
            O => \N__41295\,
            I => \N__41289\
        );

    \I__10151\ : Span4Mux_v
    port map (
            O => \N__41292\,
            I => \N__41285\
        );

    \I__10150\ : InMux
    port map (
            O => \N__41289\,
            I => \N__41282\
        );

    \I__10149\ : InMux
    port map (
            O => \N__41288\,
            I => \N__41279\
        );

    \I__10148\ : Odrv4
    port map (
            O => \N__41285\,
            I => \M_this_ext_address_qZ0Z_1\
        );

    \I__10147\ : LocalMux
    port map (
            O => \N__41282\,
            I => \M_this_ext_address_qZ0Z_1\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__41279\,
            I => \M_this_ext_address_qZ0Z_1\
        );

    \I__10145\ : InMux
    port map (
            O => \N__41272\,
            I => \N__41269\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__41269\,
            I => \un1_M_this_ext_address_q_cry_2_THRU_CO\
        );

    \I__10143\ : IoInMux
    port map (
            O => \N__41266\,
            I => \N__41263\
        );

    \I__10142\ : LocalMux
    port map (
            O => \N__41263\,
            I => \N__41260\
        );

    \I__10141\ : IoSpan4Mux
    port map (
            O => \N__41260\,
            I => \N__41257\
        );

    \I__10140\ : Span4Mux_s3_h
    port map (
            O => \N__41257\,
            I => \N__41253\
        );

    \I__10139\ : CascadeMux
    port map (
            O => \N__41256\,
            I => \N__41250\
        );

    \I__10138\ : Span4Mux_v
    port map (
            O => \N__41253\,
            I => \N__41246\
        );

    \I__10137\ : InMux
    port map (
            O => \N__41250\,
            I => \N__41243\
        );

    \I__10136\ : InMux
    port map (
            O => \N__41249\,
            I => \N__41240\
        );

    \I__10135\ : Odrv4
    port map (
            O => \N__41246\,
            I => \M_this_ext_address_qZ0Z_3\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__41243\,
            I => \M_this_ext_address_qZ0Z_3\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__41240\,
            I => \M_this_ext_address_qZ0Z_3\
        );

    \I__10132\ : InMux
    port map (
            O => \N__41233\,
            I => \N__41230\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__41230\,
            I => \un1_M_this_ext_address_q_cry_3_THRU_CO\
        );

    \I__10130\ : IoInMux
    port map (
            O => \N__41227\,
            I => \N__41224\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__41224\,
            I => \N__41221\
        );

    \I__10128\ : IoSpan4Mux
    port map (
            O => \N__41221\,
            I => \N__41218\
        );

    \I__10127\ : Span4Mux_s0_h
    port map (
            O => \N__41218\,
            I => \N__41215\
        );

    \I__10126\ : Span4Mux_h
    port map (
            O => \N__41215\,
            I => \N__41210\
        );

    \I__10125\ : InMux
    port map (
            O => \N__41214\,
            I => \N__41207\
        );

    \I__10124\ : InMux
    port map (
            O => \N__41213\,
            I => \N__41204\
        );

    \I__10123\ : Odrv4
    port map (
            O => \N__41210\,
            I => \M_this_ext_address_qZ0Z_4\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__41207\,
            I => \M_this_ext_address_qZ0Z_4\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__41204\,
            I => \M_this_ext_address_qZ0Z_4\
        );

    \I__10120\ : InMux
    port map (
            O => \N__41197\,
            I => \N__41194\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__41194\,
            I => \un1_M_this_ext_address_q_cry_4_THRU_CO\
        );

    \I__10118\ : IoInMux
    port map (
            O => \N__41191\,
            I => \N__41188\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__41188\,
            I => \N__41185\
        );

    \I__10116\ : IoSpan4Mux
    port map (
            O => \N__41185\,
            I => \N__41181\
        );

    \I__10115\ : CascadeMux
    port map (
            O => \N__41184\,
            I => \N__41178\
        );

    \I__10114\ : Span4Mux_s2_h
    port map (
            O => \N__41181\,
            I => \N__41174\
        );

    \I__10113\ : InMux
    port map (
            O => \N__41178\,
            I => \N__41171\
        );

    \I__10112\ : InMux
    port map (
            O => \N__41177\,
            I => \N__41168\
        );

    \I__10111\ : Odrv4
    port map (
            O => \N__41174\,
            I => \M_this_ext_address_qZ0Z_5\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__41171\,
            I => \M_this_ext_address_qZ0Z_5\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__41168\,
            I => \M_this_ext_address_qZ0Z_5\
        );

    \I__10108\ : CascadeMux
    port map (
            O => \N__41161\,
            I => \N__41157\
        );

    \I__10107\ : CascadeMux
    port map (
            O => \N__41160\,
            I => \N__41154\
        );

    \I__10106\ : InMux
    port map (
            O => \N__41157\,
            I => \N__41146\
        );

    \I__10105\ : InMux
    port map (
            O => \N__41154\,
            I => \N__41146\
        );

    \I__10104\ : CascadeMux
    port map (
            O => \N__41153\,
            I => \N__41142\
        );

    \I__10103\ : InMux
    port map (
            O => \N__41152\,
            I => \N__41137\
        );

    \I__10102\ : InMux
    port map (
            O => \N__41151\,
            I => \N__41137\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__41146\,
            I => \N__41126\
        );

    \I__10100\ : InMux
    port map (
            O => \N__41145\,
            I => \N__41123\
        );

    \I__10099\ : InMux
    port map (
            O => \N__41142\,
            I => \N__41120\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__41137\,
            I => \N__41117\
        );

    \I__10097\ : InMux
    port map (
            O => \N__41136\,
            I => \N__41104\
        );

    \I__10096\ : InMux
    port map (
            O => \N__41135\,
            I => \N__41104\
        );

    \I__10095\ : InMux
    port map (
            O => \N__41134\,
            I => \N__41104\
        );

    \I__10094\ : InMux
    port map (
            O => \N__41133\,
            I => \N__41104\
        );

    \I__10093\ : InMux
    port map (
            O => \N__41132\,
            I => \N__41104\
        );

    \I__10092\ : InMux
    port map (
            O => \N__41131\,
            I => \N__41104\
        );

    \I__10091\ : CascadeMux
    port map (
            O => \N__41130\,
            I => \N__41101\
        );

    \I__10090\ : CascadeMux
    port map (
            O => \N__41129\,
            I => \N__41098\
        );

    \I__10089\ : Span4Mux_h
    port map (
            O => \N__41126\,
            I => \N__41092\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__41123\,
            I => \N__41085\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__41120\,
            I => \N__41085\
        );

    \I__10086\ : Span4Mux_h
    port map (
            O => \N__41117\,
            I => \N__41085\
        );

    \I__10085\ : LocalMux
    port map (
            O => \N__41104\,
            I => \N__41082\
        );

    \I__10084\ : InMux
    port map (
            O => \N__41101\,
            I => \N__41079\
        );

    \I__10083\ : InMux
    port map (
            O => \N__41098\,
            I => \N__41076\
        );

    \I__10082\ : InMux
    port map (
            O => \N__41097\,
            I => \N__41069\
        );

    \I__10081\ : InMux
    port map (
            O => \N__41096\,
            I => \N__41069\
        );

    \I__10080\ : InMux
    port map (
            O => \N__41095\,
            I => \N__41069\
        );

    \I__10079\ : Span4Mux_v
    port map (
            O => \N__41092\,
            I => \N__41062\
        );

    \I__10078\ : Span4Mux_v
    port map (
            O => \N__41085\,
            I => \N__41062\
        );

    \I__10077\ : Span4Mux_h
    port map (
            O => \N__41082\,
            I => \N__41062\
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__41079\,
            I => \N__41053\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__41076\,
            I => \N__41053\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__41069\,
            I => \N__41053\
        );

    \I__10073\ : Span4Mux_h
    port map (
            O => \N__41062\,
            I => \N__41050\
        );

    \I__10072\ : InMux
    port map (
            O => \N__41061\,
            I => \N__41045\
        );

    \I__10071\ : InMux
    port map (
            O => \N__41060\,
            I => \N__41045\
        );

    \I__10070\ : Odrv12
    port map (
            O => \N__41053\,
            I => \N_773_0\
        );

    \I__10069\ : Odrv4
    port map (
            O => \N__41050\,
            I => \N_773_0\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__41045\,
            I => \N_773_0\
        );

    \I__10067\ : InMux
    port map (
            O => \N__41038\,
            I => \un1_M_this_ext_address_q_cry_14\
        );

    \I__10066\ : InMux
    port map (
            O => \N__41035\,
            I => \N__41032\
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__41032\,
            I => \N__41029\
        );

    \I__10064\ : Odrv12
    port map (
            O => \N__41029\,
            I => \un1_M_this_ext_address_q_cry_14_c_RNIMSSAZ0\
        );

    \I__10063\ : InMux
    port map (
            O => \N__41026\,
            I => \N__41023\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__41023\,
            I => \un1_M_this_ext_address_q_cry_9_c_RNI55NHZ0\
        );

    \I__10061\ : IoInMux
    port map (
            O => \N__41020\,
            I => \N__41017\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__41017\,
            I => \N__41014\
        );

    \I__10059\ : Span4Mux_s1_v
    port map (
            O => \N__41014\,
            I => \N__41011\
        );

    \I__10058\ : Span4Mux_v
    port map (
            O => \N__41011\,
            I => \N__41008\
        );

    \I__10057\ : Span4Mux_v
    port map (
            O => \N__41008\,
            I => \N__41005\
        );

    \I__10056\ : Span4Mux_h
    port map (
            O => \N__41005\,
            I => \N__41001\
        );

    \I__10055\ : InMux
    port map (
            O => \N__41004\,
            I => \N__40998\
        );

    \I__10054\ : Odrv4
    port map (
            O => \N__41001\,
            I => \M_this_ext_address_qZ0Z_10\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__40998\,
            I => \M_this_ext_address_qZ0Z_10\
        );

    \I__10052\ : InMux
    port map (
            O => \N__40993\,
            I => \N__40990\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__40990\,
            I => \N__40987\
        );

    \I__10050\ : Odrv4
    port map (
            O => \N__40987\,
            I => \un1_M_this_ext_address_q_cry_6_THRU_CO\
        );

    \I__10049\ : IoInMux
    port map (
            O => \N__40984\,
            I => \N__40981\
        );

    \I__10048\ : LocalMux
    port map (
            O => \N__40981\,
            I => \N__40978\
        );

    \I__10047\ : Span4Mux_s2_h
    port map (
            O => \N__40978\,
            I => \N__40975\
        );

    \I__10046\ : Span4Mux_h
    port map (
            O => \N__40975\,
            I => \N__40972\
        );

    \I__10045\ : Sp12to4
    port map (
            O => \N__40972\,
            I => \N__40968\
        );

    \I__10044\ : InMux
    port map (
            O => \N__40971\,
            I => \N__40964\
        );

    \I__10043\ : Span12Mux_s11_v
    port map (
            O => \N__40968\,
            I => \N__40961\
        );

    \I__10042\ : InMux
    port map (
            O => \N__40967\,
            I => \N__40958\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__40964\,
            I => \N__40955\
        );

    \I__10040\ : Odrv12
    port map (
            O => \N__40961\,
            I => \M_this_ext_address_qZ0Z_7\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__40958\,
            I => \M_this_ext_address_qZ0Z_7\
        );

    \I__10038\ : Odrv4
    port map (
            O => \N__40955\,
            I => \M_this_ext_address_qZ0Z_7\
        );

    \I__10037\ : InMux
    port map (
            O => \N__40948\,
            I => \N__40945\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__40945\,
            I => \un1_M_this_ext_address_q_cry_10_c_RNIEGOAZ0\
        );

    \I__10035\ : IoInMux
    port map (
            O => \N__40942\,
            I => \N__40939\
        );

    \I__10034\ : LocalMux
    port map (
            O => \N__40939\,
            I => \N__40936\
        );

    \I__10033\ : Span4Mux_s2_v
    port map (
            O => \N__40936\,
            I => \N__40933\
        );

    \I__10032\ : Span4Mux_h
    port map (
            O => \N__40933\,
            I => \N__40930\
        );

    \I__10031\ : Span4Mux_v
    port map (
            O => \N__40930\,
            I => \N__40926\
        );

    \I__10030\ : InMux
    port map (
            O => \N__40929\,
            I => \N__40923\
        );

    \I__10029\ : Odrv4
    port map (
            O => \N__40926\,
            I => \M_this_ext_address_qZ0Z_11\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__40923\,
            I => \M_this_ext_address_qZ0Z_11\
        );

    \I__10027\ : InMux
    port map (
            O => \N__40918\,
            I => \N__40915\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__40915\,
            I => \un1_M_this_ext_address_q_cry_11_c_RNIGJPAZ0\
        );

    \I__10025\ : IoInMux
    port map (
            O => \N__40912\,
            I => \N__40909\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__40909\,
            I => \N__40906\
        );

    \I__10023\ : Span4Mux_s1_h
    port map (
            O => \N__40906\,
            I => \N__40903\
        );

    \I__10022\ : Span4Mux_h
    port map (
            O => \N__40903\,
            I => \N__40899\
        );

    \I__10021\ : InMux
    port map (
            O => \N__40902\,
            I => \N__40896\
        );

    \I__10020\ : Odrv4
    port map (
            O => \N__40899\,
            I => \M_this_ext_address_qZ0Z_12\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__40896\,
            I => \M_this_ext_address_qZ0Z_12\
        );

    \I__10018\ : InMux
    port map (
            O => \N__40891\,
            I => \N__40885\
        );

    \I__10017\ : InMux
    port map (
            O => \N__40890\,
            I => \N__40885\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__40885\,
            I => \N__40882\
        );

    \I__10015\ : Span4Mux_v
    port map (
            O => \N__40882\,
            I => \N__40877\
        );

    \I__10014\ : InMux
    port map (
            O => \N__40881\,
            I => \N__40874\
        );

    \I__10013\ : InMux
    port map (
            O => \N__40880\,
            I => \N__40871\
        );

    \I__10012\ : Span4Mux_v
    port map (
            O => \N__40877\,
            I => \N__40866\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__40874\,
            I => \N__40866\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__40871\,
            I => \N__40863\
        );

    \I__10009\ : Span4Mux_h
    port map (
            O => \N__40866\,
            I => \N__40858\
        );

    \I__10008\ : Span4Mux_h
    port map (
            O => \N__40863\,
            I => \N__40855\
        );

    \I__10007\ : InMux
    port map (
            O => \N__40862\,
            I => \N__40852\
        );

    \I__10006\ : InMux
    port map (
            O => \N__40861\,
            I => \N__40849\
        );

    \I__10005\ : Odrv4
    port map (
            O => \N__40858\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__10004\ : Odrv4
    port map (
            O => \N__40855\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__40852\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__40849\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__10001\ : InMux
    port map (
            O => \N__40840\,
            I => \N__40836\
        );

    \I__10000\ : InMux
    port map (
            O => \N__40839\,
            I => \N__40833\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__40836\,
            I => \N__40830\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__40833\,
            I => \M_this_ctrl_flags_qZ0Z_4\
        );

    \I__9997\ : Odrv4
    port map (
            O => \N__40830\,
            I => \M_this_ctrl_flags_qZ0Z_4\
        );

    \I__9996\ : CascadeMux
    port map (
            O => \N__40825\,
            I => \N__40822\
        );

    \I__9995\ : CascadeBuf
    port map (
            O => \N__40822\,
            I => \N__40819\
        );

    \I__9994\ : CascadeMux
    port map (
            O => \N__40819\,
            I => \N__40816\
        );

    \I__9993\ : InMux
    port map (
            O => \N__40816\,
            I => \N__40813\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__40813\,
            I => \N__40809\
        );

    \I__9991\ : InMux
    port map (
            O => \N__40812\,
            I => \N__40805\
        );

    \I__9990\ : Span4Mux_s3_v
    port map (
            O => \N__40809\,
            I => \N__40802\
        );

    \I__9989\ : InMux
    port map (
            O => \N__40808\,
            I => \N__40799\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__40805\,
            I => \N__40796\
        );

    \I__9987\ : Span4Mux_v
    port map (
            O => \N__40802\,
            I => \N__40793\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__40799\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__9985\ : Odrv4
    port map (
            O => \N__40796\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__9984\ : Odrv4
    port map (
            O => \N__40793\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__9983\ : InMux
    port map (
            O => \N__40786\,
            I => \N__40779\
        );

    \I__9982\ : InMux
    port map (
            O => \N__40785\,
            I => \N__40776\
        );

    \I__9981\ : InMux
    port map (
            O => \N__40784\,
            I => \N__40773\
        );

    \I__9980\ : InMux
    port map (
            O => \N__40783\,
            I => \N__40770\
        );

    \I__9979\ : InMux
    port map (
            O => \N__40782\,
            I => \N__40767\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__40779\,
            I => \N__40764\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__40776\,
            I => \N__40760\
        );

    \I__9976\ : LocalMux
    port map (
            O => \N__40773\,
            I => \N__40757\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__40770\,
            I => \N__40752\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__40767\,
            I => \N__40752\
        );

    \I__9973\ : Span4Mux_v
    port map (
            O => \N__40764\,
            I => \N__40748\
        );

    \I__9972\ : InMux
    port map (
            O => \N__40763\,
            I => \N__40744\
        );

    \I__9971\ : Span4Mux_h
    port map (
            O => \N__40760\,
            I => \N__40739\
        );

    \I__9970\ : Span4Mux_v
    port map (
            O => \N__40757\,
            I => \N__40739\
        );

    \I__9969\ : Span4Mux_v
    port map (
            O => \N__40752\,
            I => \N__40736\
        );

    \I__9968\ : InMux
    port map (
            O => \N__40751\,
            I => \N__40733\
        );

    \I__9967\ : Span4Mux_v
    port map (
            O => \N__40748\,
            I => \N__40730\
        );

    \I__9966\ : InMux
    port map (
            O => \N__40747\,
            I => \N__40727\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__40744\,
            I => \N__40723\
        );

    \I__9964\ : Span4Mux_v
    port map (
            O => \N__40739\,
            I => \N__40718\
        );

    \I__9963\ : Span4Mux_h
    port map (
            O => \N__40736\,
            I => \N__40718\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__40733\,
            I => \N__40715\
        );

    \I__9961\ : Span4Mux_h
    port map (
            O => \N__40730\,
            I => \N__40710\
        );

    \I__9960\ : LocalMux
    port map (
            O => \N__40727\,
            I => \N__40710\
        );

    \I__9959\ : CascadeMux
    port map (
            O => \N__40726\,
            I => \N__40706\
        );

    \I__9958\ : Span4Mux_v
    port map (
            O => \N__40723\,
            I => \N__40702\
        );

    \I__9957\ : Span4Mux_h
    port map (
            O => \N__40718\,
            I => \N__40697\
        );

    \I__9956\ : Span4Mux_v
    port map (
            O => \N__40715\,
            I => \N__40697\
        );

    \I__9955\ : Span4Mux_h
    port map (
            O => \N__40710\,
            I => \N__40694\
        );

    \I__9954\ : InMux
    port map (
            O => \N__40709\,
            I => \N__40689\
        );

    \I__9953\ : InMux
    port map (
            O => \N__40706\,
            I => \N__40689\
        );

    \I__9952\ : InMux
    port map (
            O => \N__40705\,
            I => \N__40686\
        );

    \I__9951\ : Sp12to4
    port map (
            O => \N__40702\,
            I => \N__40680\
        );

    \I__9950\ : Sp12to4
    port map (
            O => \N__40697\,
            I => \N__40680\
        );

    \I__9949\ : Span4Mux_v
    port map (
            O => \N__40694\,
            I => \N__40677\
        );

    \I__9948\ : LocalMux
    port map (
            O => \N__40689\,
            I => \N__40672\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__40686\,
            I => \N__40672\
        );

    \I__9946\ : InMux
    port map (
            O => \N__40685\,
            I => \N__40669\
        );

    \I__9945\ : Span12Mux_h
    port map (
            O => \N__40680\,
            I => \N__40662\
        );

    \I__9944\ : Sp12to4
    port map (
            O => \N__40677\,
            I => \N__40662\
        );

    \I__9943\ : Span12Mux_v
    port map (
            O => \N__40672\,
            I => \N__40662\
        );

    \I__9942\ : LocalMux
    port map (
            O => \N__40669\,
            I => \N__40659\
        );

    \I__9941\ : Odrv12
    port map (
            O => \N__40662\,
            I => port_data_in_4
        );

    \I__9940\ : Odrv12
    port map (
            O => \N__40659\,
            I => port_data_in_4
        );

    \I__9939\ : CascadeMux
    port map (
            O => \N__40654\,
            I => \N_1081_cascade_\
        );

    \I__9938\ : InMux
    port map (
            O => \N__40651\,
            I => \N__40648\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__40648\,
            I => \N__40645\
        );

    \I__9936\ : Odrv4
    port map (
            O => \N__40645\,
            I => \M_this_map_address_qc_1_1\
        );

    \I__9935\ : InMux
    port map (
            O => \N__40642\,
            I => \un1_M_this_ext_address_q_cry_6\
        );

    \I__9934\ : InMux
    port map (
            O => \N__40639\,
            I => \bfn_26_22_0_\
        );

    \I__9933\ : IoInMux
    port map (
            O => \N__40636\,
            I => \N__40633\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__40633\,
            I => \N__40630\
        );

    \I__9931\ : IoSpan4Mux
    port map (
            O => \N__40630\,
            I => \N__40627\
        );

    \I__9930\ : Span4Mux_s2_v
    port map (
            O => \N__40627\,
            I => \N__40623\
        );

    \I__9929\ : InMux
    port map (
            O => \N__40626\,
            I => \N__40620\
        );

    \I__9928\ : Span4Mux_v
    port map (
            O => \N__40623\,
            I => \N__40617\
        );

    \I__9927\ : LocalMux
    port map (
            O => \N__40620\,
            I => \N__40614\
        );

    \I__9926\ : Span4Mux_v
    port map (
            O => \N__40617\,
            I => \N__40609\
        );

    \I__9925\ : Span4Mux_h
    port map (
            O => \N__40614\,
            I => \N__40609\
        );

    \I__9924\ : Odrv4
    port map (
            O => \N__40609\,
            I => \M_this_ext_address_qZ0Z_9\
        );

    \I__9923\ : InMux
    port map (
            O => \N__40606\,
            I => \N__40603\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__40603\,
            I => \N__40600\
        );

    \I__9921\ : Span4Mux_h
    port map (
            O => \N__40600\,
            I => \N__40597\
        );

    \I__9920\ : Odrv4
    port map (
            O => \N__40597\,
            I => \un1_M_this_ext_address_q_cry_8_c_RNIS45FZ0\
        );

    \I__9919\ : InMux
    port map (
            O => \N__40594\,
            I => \un1_M_this_ext_address_q_cry_8\
        );

    \I__9918\ : InMux
    port map (
            O => \N__40591\,
            I => \un1_M_this_ext_address_q_cry_9\
        );

    \I__9917\ : InMux
    port map (
            O => \N__40588\,
            I => \un1_M_this_ext_address_q_cry_10\
        );

    \I__9916\ : InMux
    port map (
            O => \N__40585\,
            I => \un1_M_this_ext_address_q_cry_11\
        );

    \I__9915\ : IoInMux
    port map (
            O => \N__40582\,
            I => \N__40579\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__40579\,
            I => \N__40576\
        );

    \I__9913\ : IoSpan4Mux
    port map (
            O => \N__40576\,
            I => \N__40573\
        );

    \I__9912\ : Span4Mux_s2_h
    port map (
            O => \N__40573\,
            I => \N__40569\
        );

    \I__9911\ : InMux
    port map (
            O => \N__40572\,
            I => \N__40566\
        );

    \I__9910\ : Span4Mux_h
    port map (
            O => \N__40569\,
            I => \N__40561\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__40566\,
            I => \N__40561\
        );

    \I__9908\ : Span4Mux_v
    port map (
            O => \N__40561\,
            I => \N__40558\
        );

    \I__9907\ : Odrv4
    port map (
            O => \N__40558\,
            I => \M_this_ext_address_qZ0Z_13\
        );

    \I__9906\ : InMux
    port map (
            O => \N__40555\,
            I => \N__40552\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__40552\,
            I => \N__40549\
        );

    \I__9904\ : Odrv12
    port map (
            O => \N__40549\,
            I => \un1_M_this_ext_address_q_cry_12_c_RNIIMQAZ0\
        );

    \I__9903\ : InMux
    port map (
            O => \N__40546\,
            I => \un1_M_this_ext_address_q_cry_12\
        );

    \I__9902\ : IoInMux
    port map (
            O => \N__40543\,
            I => \N__40540\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__40540\,
            I => \N__40537\
        );

    \I__9900\ : Span4Mux_s2_h
    port map (
            O => \N__40537\,
            I => \N__40533\
        );

    \I__9899\ : InMux
    port map (
            O => \N__40536\,
            I => \N__40530\
        );

    \I__9898\ : Span4Mux_h
    port map (
            O => \N__40533\,
            I => \N__40527\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__40530\,
            I => \N__40524\
        );

    \I__9896\ : Odrv4
    port map (
            O => \N__40527\,
            I => \M_this_ext_address_qZ0Z_14\
        );

    \I__9895\ : Odrv12
    port map (
            O => \N__40524\,
            I => \M_this_ext_address_qZ0Z_14\
        );

    \I__9894\ : InMux
    port map (
            O => \N__40519\,
            I => \N__40516\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__40516\,
            I => \N__40513\
        );

    \I__9892\ : Odrv12
    port map (
            O => \N__40513\,
            I => \un1_M_this_ext_address_q_cry_13_c_RNIKPRAZ0\
        );

    \I__9891\ : InMux
    port map (
            O => \N__40510\,
            I => \un1_M_this_ext_address_q_cry_13\
        );

    \I__9890\ : IoInMux
    port map (
            O => \N__40507\,
            I => \N__40504\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__40504\,
            I => \N__40500\
        );

    \I__9888\ : InMux
    port map (
            O => \N__40503\,
            I => \N__40497\
        );

    \I__9887\ : Span12Mux_s1_h
    port map (
            O => \N__40500\,
            I => \N__40494\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__40497\,
            I => \N__40491\
        );

    \I__9885\ : Span12Mux_v
    port map (
            O => \N__40494\,
            I => \N__40488\
        );

    \I__9884\ : Span4Mux_v
    port map (
            O => \N__40491\,
            I => \N__40485\
        );

    \I__9883\ : Odrv12
    port map (
            O => \N__40488\,
            I => \M_this_ext_address_qZ0Z_15\
        );

    \I__9882\ : Odrv4
    port map (
            O => \N__40485\,
            I => \M_this_ext_address_qZ0Z_15\
        );

    \I__9881\ : CascadeMux
    port map (
            O => \N__40480\,
            I => \N__40476\
        );

    \I__9880\ : InMux
    port map (
            O => \N__40479\,
            I => \N__40473\
        );

    \I__9879\ : InMux
    port map (
            O => \N__40476\,
            I => \N__40470\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__40473\,
            I => \N__40467\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__40470\,
            I => \N__40464\
        );

    \I__9876\ : Span4Mux_v
    port map (
            O => \N__40467\,
            I => \N__40459\
        );

    \I__9875\ : Span4Mux_v
    port map (
            O => \N__40464\,
            I => \N__40459\
        );

    \I__9874\ : Span4Mux_h
    port map (
            O => \N__40459\,
            I => \N__40455\
        );

    \I__9873\ : InMux
    port map (
            O => \N__40458\,
            I => \N__40452\
        );

    \I__9872\ : Span4Mux_h
    port map (
            O => \N__40455\,
            I => \N__40449\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__40452\,
            I => \M_this_ctrl_flags_qZ0Z_6\
        );

    \I__9870\ : Odrv4
    port map (
            O => \N__40449\,
            I => \M_this_ctrl_flags_qZ0Z_6\
        );

    \I__9869\ : InMux
    port map (
            O => \N__40444\,
            I => \N__40440\
        );

    \I__9868\ : InMux
    port map (
            O => \N__40443\,
            I => \N__40437\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__40440\,
            I => \N__40430\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__40437\,
            I => \N__40430\
        );

    \I__9865\ : CascadeMux
    port map (
            O => \N__40436\,
            I => \N__40427\
        );

    \I__9864\ : InMux
    port map (
            O => \N__40435\,
            I => \N__40424\
        );

    \I__9863\ : Span4Mux_v
    port map (
            O => \N__40430\,
            I => \N__40421\
        );

    \I__9862\ : InMux
    port map (
            O => \N__40427\,
            I => \N__40416\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__40424\,
            I => \N__40412\
        );

    \I__9860\ : Span4Mux_h
    port map (
            O => \N__40421\,
            I => \N__40408\
        );

    \I__9859\ : InMux
    port map (
            O => \N__40420\,
            I => \N__40405\
        );

    \I__9858\ : CascadeMux
    port map (
            O => \N__40419\,
            I => \N__40401\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__40416\,
            I => \N__40398\
        );

    \I__9856\ : InMux
    port map (
            O => \N__40415\,
            I => \N__40394\
        );

    \I__9855\ : Span4Mux_v
    port map (
            O => \N__40412\,
            I => \N__40391\
        );

    \I__9854\ : InMux
    port map (
            O => \N__40411\,
            I => \N__40388\
        );

    \I__9853\ : Span4Mux_v
    port map (
            O => \N__40408\,
            I => \N__40383\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__40405\,
            I => \N__40383\
        );

    \I__9851\ : InMux
    port map (
            O => \N__40404\,
            I => \N__40378\
        );

    \I__9850\ : InMux
    port map (
            O => \N__40401\,
            I => \N__40378\
        );

    \I__9849\ : Span4Mux_v
    port map (
            O => \N__40398\,
            I => \N__40375\
        );

    \I__9848\ : InMux
    port map (
            O => \N__40397\,
            I => \N__40372\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__40394\,
            I => \N__40369\
        );

    \I__9846\ : Span4Mux_h
    port map (
            O => \N__40391\,
            I => \N__40364\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__40388\,
            I => \N__40364\
        );

    \I__9844\ : Span4Mux_v
    port map (
            O => \N__40383\,
            I => \N__40361\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__40378\,
            I => \N__40358\
        );

    \I__9842\ : Span4Mux_h
    port map (
            O => \N__40375\,
            I => \N__40355\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__40372\,
            I => \N__40352\
        );

    \I__9840\ : Span12Mux_h
    port map (
            O => \N__40369\,
            I => \N__40347\
        );

    \I__9839\ : Sp12to4
    port map (
            O => \N__40364\,
            I => \N__40347\
        );

    \I__9838\ : Span4Mux_v
    port map (
            O => \N__40361\,
            I => \N__40344\
        );

    \I__9837\ : Span4Mux_v
    port map (
            O => \N__40358\,
            I => \N__40341\
        );

    \I__9836\ : Sp12to4
    port map (
            O => \N__40355\,
            I => \N__40336\
        );

    \I__9835\ : Span12Mux_s9_v
    port map (
            O => \N__40352\,
            I => \N__40336\
        );

    \I__9834\ : Span12Mux_v
    port map (
            O => \N__40347\,
            I => \N__40331\
        );

    \I__9833\ : Sp12to4
    port map (
            O => \N__40344\,
            I => \N__40331\
        );

    \I__9832\ : Span4Mux_h
    port map (
            O => \N__40341\,
            I => \N__40328\
        );

    \I__9831\ : Span12Mux_v
    port map (
            O => \N__40336\,
            I => \N__40325\
        );

    \I__9830\ : Span12Mux_h
    port map (
            O => \N__40331\,
            I => \N__40322\
        );

    \I__9829\ : Span4Mux_v
    port map (
            O => \N__40328\,
            I => \N__40319\
        );

    \I__9828\ : Odrv12
    port map (
            O => \N__40325\,
            I => port_data_in_6
        );

    \I__9827\ : Odrv12
    port map (
            O => \N__40322\,
            I => port_data_in_6
        );

    \I__9826\ : Odrv4
    port map (
            O => \N__40319\,
            I => port_data_in_6
        );

    \I__9825\ : InMux
    port map (
            O => \N__40312\,
            I => \N__40308\
        );

    \I__9824\ : InMux
    port map (
            O => \N__40311\,
            I => \N__40305\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__40308\,
            I => \N__40300\
        );

    \I__9822\ : LocalMux
    port map (
            O => \N__40305\,
            I => \N__40300\
        );

    \I__9821\ : Span4Mux_h
    port map (
            O => \N__40300\,
            I => \N__40297\
        );

    \I__9820\ : Span4Mux_h
    port map (
            O => \N__40297\,
            I => \N__40294\
        );

    \I__9819\ : Odrv4
    port map (
            O => \N__40294\,
            I => \N_247\
        );

    \I__9818\ : IoInMux
    port map (
            O => \N__40291\,
            I => \N__40288\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__40288\,
            I => \N__40285\
        );

    \I__9816\ : IoSpan4Mux
    port map (
            O => \N__40285\,
            I => \N__40282\
        );

    \I__9815\ : Span4Mux_s3_v
    port map (
            O => \N__40282\,
            I => \N__40277\
        );

    \I__9814\ : CascadeMux
    port map (
            O => \N__40281\,
            I => \N__40274\
        );

    \I__9813\ : CascadeMux
    port map (
            O => \N__40280\,
            I => \N__40271\
        );

    \I__9812\ : Sp12to4
    port map (
            O => \N__40277\,
            I => \N__40268\
        );

    \I__9811\ : InMux
    port map (
            O => \N__40274\,
            I => \N__40265\
        );

    \I__9810\ : InMux
    port map (
            O => \N__40271\,
            I => \N__40262\
        );

    \I__9809\ : Span12Mux_s11_v
    port map (
            O => \N__40268\,
            I => \N__40259\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__40265\,
            I => \N__40254\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__40262\,
            I => \N__40254\
        );

    \I__9806\ : Odrv12
    port map (
            O => \N__40259\,
            I => \M_this_ext_address_qZ0Z_0\
        );

    \I__9805\ : Odrv4
    port map (
            O => \N__40254\,
            I => \M_this_ext_address_qZ0Z_0\
        );

    \I__9804\ : InMux
    port map (
            O => \N__40249\,
            I => \un1_M_this_ext_address_q_cry_0\
        );

    \I__9803\ : IoInMux
    port map (
            O => \N__40246\,
            I => \N__40243\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__40243\,
            I => \N__40240\
        );

    \I__9801\ : IoSpan4Mux
    port map (
            O => \N__40240\,
            I => \N__40237\
        );

    \I__9800\ : Span4Mux_s3_v
    port map (
            O => \N__40237\,
            I => \N__40233\
        );

    \I__9799\ : CascadeMux
    port map (
            O => \N__40236\,
            I => \N__40229\
        );

    \I__9798\ : Span4Mux_v
    port map (
            O => \N__40233\,
            I => \N__40226\
        );

    \I__9797\ : InMux
    port map (
            O => \N__40232\,
            I => \N__40223\
        );

    \I__9796\ : InMux
    port map (
            O => \N__40229\,
            I => \N__40220\
        );

    \I__9795\ : Span4Mux_v
    port map (
            O => \N__40226\,
            I => \N__40215\
        );

    \I__9794\ : LocalMux
    port map (
            O => \N__40223\,
            I => \N__40215\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__40220\,
            I => \M_this_ext_address_qZ0Z_2\
        );

    \I__9792\ : Odrv4
    port map (
            O => \N__40215\,
            I => \M_this_ext_address_qZ0Z_2\
        );

    \I__9791\ : InMux
    port map (
            O => \N__40210\,
            I => \N__40207\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__40207\,
            I => \N__40204\
        );

    \I__9789\ : Odrv4
    port map (
            O => \N__40204\,
            I => \un1_M_this_ext_address_q_cry_1_THRU_CO\
        );

    \I__9788\ : InMux
    port map (
            O => \N__40201\,
            I => \un1_M_this_ext_address_q_cry_1\
        );

    \I__9787\ : InMux
    port map (
            O => \N__40198\,
            I => \un1_M_this_ext_address_q_cry_2\
        );

    \I__9786\ : InMux
    port map (
            O => \N__40195\,
            I => \un1_M_this_ext_address_q_cry_3\
        );

    \I__9785\ : InMux
    port map (
            O => \N__40192\,
            I => \un1_M_this_ext_address_q_cry_4\
        );

    \I__9784\ : InMux
    port map (
            O => \N__40189\,
            I => \un1_M_this_ext_address_q_cry_5\
        );

    \I__9783\ : InMux
    port map (
            O => \N__40186\,
            I => \N__40183\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__40183\,
            I => \N_919_0\
        );

    \I__9781\ : InMux
    port map (
            O => \N__40180\,
            I => \N__40177\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__40177\,
            I => \N__40174\
        );

    \I__9779\ : Odrv4
    port map (
            O => \N__40174\,
            I => \N_923_0\
        );

    \I__9778\ : InMux
    port map (
            O => \N__40171\,
            I => \N__40168\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__40168\,
            I => \N_920_0\
        );

    \I__9776\ : InMux
    port map (
            O => \N__40165\,
            I => \N__40162\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__40162\,
            I => \N__40159\
        );

    \I__9774\ : Odrv4
    port map (
            O => \N__40159\,
            I => \N_922_0\
        );

    \I__9773\ : CEMux
    port map (
            O => \N__40156\,
            I => \N__40146\
        );

    \I__9772\ : InMux
    port map (
            O => \N__40155\,
            I => \N__40141\
        );

    \I__9771\ : InMux
    port map (
            O => \N__40154\,
            I => \N__40141\
        );

    \I__9770\ : InMux
    port map (
            O => \N__40153\,
            I => \N__40136\
        );

    \I__9769\ : InMux
    port map (
            O => \N__40152\,
            I => \N__40136\
        );

    \I__9768\ : InMux
    port map (
            O => \N__40151\,
            I => \N__40133\
        );

    \I__9767\ : InMux
    port map (
            O => \N__40150\,
            I => \N__40130\
        );

    \I__9766\ : CEMux
    port map (
            O => \N__40149\,
            I => \N__40126\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__40146\,
            I => \N__40123\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__40141\,
            I => \N__40113\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__40136\,
            I => \N__40113\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__40133\,
            I => \N__40113\
        );

    \I__9761\ : LocalMux
    port map (
            O => \N__40130\,
            I => \N__40113\
        );

    \I__9760\ : InMux
    port map (
            O => \N__40129\,
            I => \N__40110\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__40126\,
            I => \N__40107\
        );

    \I__9758\ : Span4Mux_s2_v
    port map (
            O => \N__40123\,
            I => \N__40104\
        );

    \I__9757\ : InMux
    port map (
            O => \N__40122\,
            I => \N__40101\
        );

    \I__9756\ : Span4Mux_v
    port map (
            O => \N__40113\,
            I => \N__40096\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__40110\,
            I => \N__40096\
        );

    \I__9754\ : Span4Mux_h
    port map (
            O => \N__40107\,
            I => \N__40093\
        );

    \I__9753\ : Span4Mux_h
    port map (
            O => \N__40104\,
            I => \N__40088\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__40101\,
            I => \N__40088\
        );

    \I__9751\ : Span4Mux_v
    port map (
            O => \N__40096\,
            I => \N__40085\
        );

    \I__9750\ : Span4Mux_v
    port map (
            O => \N__40093\,
            I => \N__40080\
        );

    \I__9749\ : Span4Mux_v
    port map (
            O => \N__40088\,
            I => \N__40080\
        );

    \I__9748\ : Odrv4
    port map (
            O => \N__40085\,
            I => \N_296_0\
        );

    \I__9747\ : Odrv4
    port map (
            O => \N__40080\,
            I => \N_296_0\
        );

    \I__9746\ : InMux
    port map (
            O => \N__40075\,
            I => \N__40072\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__40072\,
            I => \N_924_0\
        );

    \I__9744\ : InMux
    port map (
            O => \N__40069\,
            I => \N__40065\
        );

    \I__9743\ : InMux
    port map (
            O => \N__40068\,
            I => \N__40062\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__40065\,
            I => \N__40053\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__40062\,
            I => \N__40053\
        );

    \I__9740\ : InMux
    port map (
            O => \N__40061\,
            I => \N__40049\
        );

    \I__9739\ : InMux
    port map (
            O => \N__40060\,
            I => \N__40046\
        );

    \I__9738\ : InMux
    port map (
            O => \N__40059\,
            I => \N__40043\
        );

    \I__9737\ : InMux
    port map (
            O => \N__40058\,
            I => \N__40040\
        );

    \I__9736\ : Span4Mux_v
    port map (
            O => \N__40053\,
            I => \N__40036\
        );

    \I__9735\ : CascadeMux
    port map (
            O => \N__40052\,
            I => \N__40033\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__40049\,
            I => \N__40029\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__40046\,
            I => \N__40022\
        );

    \I__9732\ : LocalMux
    port map (
            O => \N__40043\,
            I => \N__40022\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__40040\,
            I => \N__40022\
        );

    \I__9730\ : InMux
    port map (
            O => \N__40039\,
            I => \N__40019\
        );

    \I__9729\ : Span4Mux_h
    port map (
            O => \N__40036\,
            I => \N__40016\
        );

    \I__9728\ : InMux
    port map (
            O => \N__40033\,
            I => \N__40013\
        );

    \I__9727\ : CascadeMux
    port map (
            O => \N__40032\,
            I => \N__40009\
        );

    \I__9726\ : Span4Mux_v
    port map (
            O => \N__40029\,
            I => \N__40006\
        );

    \I__9725\ : Span4Mux_v
    port map (
            O => \N__40022\,
            I => \N__40003\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__40019\,
            I => \N__40000\
        );

    \I__9723\ : Span4Mux_h
    port map (
            O => \N__40016\,
            I => \N__39995\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__40013\,
            I => \N__39995\
        );

    \I__9721\ : InMux
    port map (
            O => \N__40012\,
            I => \N__39990\
        );

    \I__9720\ : InMux
    port map (
            O => \N__40009\,
            I => \N__39990\
        );

    \I__9719\ : Span4Mux_v
    port map (
            O => \N__40006\,
            I => \N__39987\
        );

    \I__9718\ : Span4Mux_v
    port map (
            O => \N__40003\,
            I => \N__39982\
        );

    \I__9717\ : Span4Mux_v
    port map (
            O => \N__40000\,
            I => \N__39982\
        );

    \I__9716\ : Span4Mux_v
    port map (
            O => \N__39995\,
            I => \N__39979\
        );

    \I__9715\ : LocalMux
    port map (
            O => \N__39990\,
            I => \N__39976\
        );

    \I__9714\ : Span4Mux_v
    port map (
            O => \N__39987\,
            I => \N__39973\
        );

    \I__9713\ : Sp12to4
    port map (
            O => \N__39982\,
            I => \N__39970\
        );

    \I__9712\ : Span4Mux_h
    port map (
            O => \N__39979\,
            I => \N__39965\
        );

    \I__9711\ : Span4Mux_v
    port map (
            O => \N__39976\,
            I => \N__39965\
        );

    \I__9710\ : Sp12to4
    port map (
            O => \N__39973\,
            I => \N__39960\
        );

    \I__9709\ : Span12Mux_h
    port map (
            O => \N__39970\,
            I => \N__39960\
        );

    \I__9708\ : Span4Mux_h
    port map (
            O => \N__39965\,
            I => \N__39957\
        );

    \I__9707\ : Odrv12
    port map (
            O => \N__39960\,
            I => port_data_in_5
        );

    \I__9706\ : Odrv4
    port map (
            O => \N__39957\,
            I => port_data_in_5
        );

    \I__9705\ : CascadeMux
    port map (
            O => \N__39952\,
            I => \N__39949\
        );

    \I__9704\ : InMux
    port map (
            O => \N__39949\,
            I => \N__39946\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__39946\,
            I => \N__39942\
        );

    \I__9702\ : InMux
    port map (
            O => \N__39945\,
            I => \N__39939\
        );

    \I__9701\ : Span12Mux_h
    port map (
            O => \N__39942\,
            I => \N__39936\
        );

    \I__9700\ : LocalMux
    port map (
            O => \N__39939\,
            I => \M_this_ctrl_flags_qZ0Z_5\
        );

    \I__9699\ : Odrv12
    port map (
            O => \N__39936\,
            I => \M_this_ctrl_flags_qZ0Z_5\
        );

    \I__9698\ : InMux
    port map (
            O => \N__39931\,
            I => \N__39928\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__39928\,
            I => \N__39923\
        );

    \I__9696\ : InMux
    port map (
            O => \N__39927\,
            I => \N__39920\
        );

    \I__9695\ : InMux
    port map (
            O => \N__39926\,
            I => \N__39917\
        );

    \I__9694\ : Span4Mux_h
    port map (
            O => \N__39923\,
            I => \N__39910\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__39920\,
            I => \N__39910\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__39917\,
            I => \N__39910\
        );

    \I__9691\ : Span4Mux_v
    port map (
            O => \N__39910\,
            I => \N__39907\
        );

    \I__9690\ : Span4Mux_h
    port map (
            O => \N__39907\,
            I => \N__39902\
        );

    \I__9689\ : InMux
    port map (
            O => \N__39906\,
            I => \N__39899\
        );

    \I__9688\ : InMux
    port map (
            O => \N__39905\,
            I => \N__39894\
        );

    \I__9687\ : Span4Mux_v
    port map (
            O => \N__39902\,
            I => \N__39889\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__39899\,
            I => \N__39889\
        );

    \I__9685\ : CascadeMux
    port map (
            O => \N__39898\,
            I => \N__39886\
        );

    \I__9684\ : CascadeMux
    port map (
            O => \N__39897\,
            I => \N__39883\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__39894\,
            I => \N__39880\
        );

    \I__9682\ : Span4Mux_h
    port map (
            O => \N__39889\,
            I => \N__39877\
        );

    \I__9681\ : InMux
    port map (
            O => \N__39886\,
            I => \N__39874\
        );

    \I__9680\ : InMux
    port map (
            O => \N__39883\,
            I => \N__39871\
        );

    \I__9679\ : Span4Mux_h
    port map (
            O => \N__39880\,
            I => \N__39867\
        );

    \I__9678\ : Span4Mux_h
    port map (
            O => \N__39877\,
            I => \N__39860\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__39874\,
            I => \N__39860\
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__39871\,
            I => \N__39860\
        );

    \I__9675\ : InMux
    port map (
            O => \N__39870\,
            I => \N__39857\
        );

    \I__9674\ : Span4Mux_v
    port map (
            O => \N__39867\,
            I => \N__39853\
        );

    \I__9673\ : Span4Mux_v
    port map (
            O => \N__39860\,
            I => \N__39850\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__39857\,
            I => \N__39847\
        );

    \I__9671\ : InMux
    port map (
            O => \N__39856\,
            I => \N__39844\
        );

    \I__9670\ : Span4Mux_v
    port map (
            O => \N__39853\,
            I => \N__39839\
        );

    \I__9669\ : Span4Mux_h
    port map (
            O => \N__39850\,
            I => \N__39839\
        );

    \I__9668\ : Span12Mux_s10_v
    port map (
            O => \N__39847\,
            I => \N__39835\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__39844\,
            I => \N__39832\
        );

    \I__9666\ : Sp12to4
    port map (
            O => \N__39839\,
            I => \N__39829\
        );

    \I__9665\ : InMux
    port map (
            O => \N__39838\,
            I => \N__39826\
        );

    \I__9664\ : Span12Mux_v
    port map (
            O => \N__39835\,
            I => \N__39823\
        );

    \I__9663\ : Span12Mux_h
    port map (
            O => \N__39832\,
            I => \N__39816\
        );

    \I__9662\ : Span12Mux_s6_h
    port map (
            O => \N__39829\,
            I => \N__39816\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__39826\,
            I => \N__39816\
        );

    \I__9660\ : Span12Mux_h
    port map (
            O => \N__39823\,
            I => \N__39813\
        );

    \I__9659\ : Span12Mux_v
    port map (
            O => \N__39816\,
            I => \N__39810\
        );

    \I__9658\ : Odrv12
    port map (
            O => \N__39813\,
            I => port_data_in_7
        );

    \I__9657\ : Odrv12
    port map (
            O => \N__39810\,
            I => port_data_in_7
        );

    \I__9656\ : InMux
    port map (
            O => \N__39805\,
            I => \un1_M_this_map_address_q_cry_5\
        );

    \I__9655\ : InMux
    port map (
            O => \N__39802\,
            I => \un1_M_this_map_address_q_cry_6\
        );

    \I__9654\ : InMux
    port map (
            O => \N__39799\,
            I => \bfn_24_24_0_\
        );

    \I__9653\ : InMux
    port map (
            O => \N__39796\,
            I => \un1_M_this_map_address_q_cry_8\
        );

    \I__9652\ : InMux
    port map (
            O => \N__39793\,
            I => \N__39790\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__39790\,
            I => \N__39787\
        );

    \I__9650\ : Odrv4
    port map (
            O => \N__39787\,
            I => \un1_M_this_map_address_q_cry_5_THRU_CO\
        );

    \I__9649\ : InMux
    port map (
            O => \N__39784\,
            I => \N__39778\
        );

    \I__9648\ : InMux
    port map (
            O => \N__39783\,
            I => \N__39774\
        );

    \I__9647\ : InMux
    port map (
            O => \N__39782\,
            I => \N__39771\
        );

    \I__9646\ : InMux
    port map (
            O => \N__39781\,
            I => \N__39768\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__39778\,
            I => \N__39765\
        );

    \I__9644\ : InMux
    port map (
            O => \N__39777\,
            I => \N__39762\
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__39774\,
            I => \N__39757\
        );

    \I__9642\ : LocalMux
    port map (
            O => \N__39771\,
            I => \N__39754\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__39768\,
            I => \N__39750\
        );

    \I__9640\ : Span4Mux_v
    port map (
            O => \N__39765\,
            I => \N__39745\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__39762\,
            I => \N__39745\
        );

    \I__9638\ : InMux
    port map (
            O => \N__39761\,
            I => \N__39742\
        );

    \I__9637\ : InMux
    port map (
            O => \N__39760\,
            I => \N__39739\
        );

    \I__9636\ : Span4Mux_h
    port map (
            O => \N__39757\,
            I => \N__39736\
        );

    \I__9635\ : Span4Mux_h
    port map (
            O => \N__39754\,
            I => \N__39733\
        );

    \I__9634\ : InMux
    port map (
            O => \N__39753\,
            I => \N__39730\
        );

    \I__9633\ : Span4Mux_v
    port map (
            O => \N__39750\,
            I => \N__39725\
        );

    \I__9632\ : Span4Mux_v
    port map (
            O => \N__39745\,
            I => \N__39720\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__39742\,
            I => \N__39720\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__39739\,
            I => \N__39717\
        );

    \I__9629\ : Span4Mux_h
    port map (
            O => \N__39736\,
            I => \N__39710\
        );

    \I__9628\ : Span4Mux_v
    port map (
            O => \N__39733\,
            I => \N__39710\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__39730\,
            I => \N__39710\
        );

    \I__9626\ : InMux
    port map (
            O => \N__39729\,
            I => \N__39707\
        );

    \I__9625\ : InMux
    port map (
            O => \N__39728\,
            I => \N__39704\
        );

    \I__9624\ : Span4Mux_v
    port map (
            O => \N__39725\,
            I => \N__39701\
        );

    \I__9623\ : Span4Mux_v
    port map (
            O => \N__39720\,
            I => \N__39698\
        );

    \I__9622\ : Span4Mux_v
    port map (
            O => \N__39717\,
            I => \N__39695\
        );

    \I__9621\ : Span4Mux_h
    port map (
            O => \N__39710\,
            I => \N__39690\
        );

    \I__9620\ : LocalMux
    port map (
            O => \N__39707\,
            I => \N__39690\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__39704\,
            I => \N__39687\
        );

    \I__9618\ : Sp12to4
    port map (
            O => \N__39701\,
            I => \N__39681\
        );

    \I__9617\ : Sp12to4
    port map (
            O => \N__39698\,
            I => \N__39681\
        );

    \I__9616\ : Span4Mux_v
    port map (
            O => \N__39695\,
            I => \N__39678\
        );

    \I__9615\ : Span4Mux_v
    port map (
            O => \N__39690\,
            I => \N__39673\
        );

    \I__9614\ : Span4Mux_h
    port map (
            O => \N__39687\,
            I => \N__39673\
        );

    \I__9613\ : InMux
    port map (
            O => \N__39686\,
            I => \N__39670\
        );

    \I__9612\ : Span12Mux_h
    port map (
            O => \N__39681\,
            I => \N__39667\
        );

    \I__9611\ : IoSpan4Mux
    port map (
            O => \N__39678\,
            I => \N__39664\
        );

    \I__9610\ : Span4Mux_v
    port map (
            O => \N__39673\,
            I => \N__39661\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__39670\,
            I => \N__39658\
        );

    \I__9608\ : Odrv12
    port map (
            O => \N__39667\,
            I => port_data_in_1
        );

    \I__9607\ : Odrv4
    port map (
            O => \N__39664\,
            I => port_data_in_1
        );

    \I__9606\ : Odrv4
    port map (
            O => \N__39661\,
            I => port_data_in_1
        );

    \I__9605\ : Odrv12
    port map (
            O => \N__39658\,
            I => port_data_in_1
        );

    \I__9604\ : CascadeMux
    port map (
            O => \N__39649\,
            I => \M_this_map_address_qc_8_1_cascade_\
        );

    \I__9603\ : CascadeMux
    port map (
            O => \N__39646\,
            I => \N__39643\
        );

    \I__9602\ : CascadeBuf
    port map (
            O => \N__39643\,
            I => \N__39640\
        );

    \I__9601\ : CascadeMux
    port map (
            O => \N__39640\,
            I => \N__39637\
        );

    \I__9600\ : InMux
    port map (
            O => \N__39637\,
            I => \N__39634\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__39634\,
            I => \N__39629\
        );

    \I__9598\ : CascadeMux
    port map (
            O => \N__39633\,
            I => \N__39626\
        );

    \I__9597\ : InMux
    port map (
            O => \N__39632\,
            I => \N__39623\
        );

    \I__9596\ : Span4Mux_s1_v
    port map (
            O => \N__39629\,
            I => \N__39620\
        );

    \I__9595\ : InMux
    port map (
            O => \N__39626\,
            I => \N__39617\
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__39623\,
            I => \N__39614\
        );

    \I__9593\ : Span4Mux_v
    port map (
            O => \N__39620\,
            I => \N__39611\
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__39617\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__9591\ : Odrv4
    port map (
            O => \N__39614\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__39611\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__9589\ : InMux
    port map (
            O => \N__39604\,
            I => \N__39601\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__39601\,
            I => \un1_M_this_map_address_q_cry_7_THRU_CO\
        );

    \I__9587\ : InMux
    port map (
            O => \N__39598\,
            I => \N__39595\
        );

    \I__9586\ : LocalMux
    port map (
            O => \N__39595\,
            I => \N__39592\
        );

    \I__9585\ : Odrv4
    port map (
            O => \N__39592\,
            I => \un1_M_this_map_address_q_axb_0\
        );

    \I__9584\ : InMux
    port map (
            O => \N__39589\,
            I => \N__39586\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__39586\,
            I => \M_this_map_address_qc_2_0\
        );

    \I__9582\ : CascadeMux
    port map (
            O => \N__39583\,
            I => \N__39580\
        );

    \I__9581\ : InMux
    port map (
            O => \N__39580\,
            I => \N__39577\
        );

    \I__9580\ : LocalMux
    port map (
            O => \N__39577\,
            I => \N_1097\
        );

    \I__9579\ : CascadeMux
    port map (
            O => \N__39574\,
            I => \N__39571\
        );

    \I__9578\ : CascadeBuf
    port map (
            O => \N__39571\,
            I => \N__39568\
        );

    \I__9577\ : CascadeMux
    port map (
            O => \N__39568\,
            I => \N__39565\
        );

    \I__9576\ : InMux
    port map (
            O => \N__39565\,
            I => \N__39559\
        );

    \I__9575\ : CascadeMux
    port map (
            O => \N__39564\,
            I => \N__39556\
        );

    \I__9574\ : InMux
    port map (
            O => \N__39563\,
            I => \N__39551\
        );

    \I__9573\ : InMux
    port map (
            O => \N__39562\,
            I => \N__39551\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__39559\,
            I => \N__39548\
        );

    \I__9571\ : InMux
    port map (
            O => \N__39556\,
            I => \N__39544\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__39551\,
            I => \N__39541\
        );

    \I__9569\ : Span4Mux_s1_v
    port map (
            O => \N__39548\,
            I => \N__39538\
        );

    \I__9568\ : InMux
    port map (
            O => \N__39547\,
            I => \N__39535\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__39544\,
            I => \N__39532\
        );

    \I__9566\ : Span4Mux_h
    port map (
            O => \N__39541\,
            I => \N__39527\
        );

    \I__9565\ : Span4Mux_v
    port map (
            O => \N__39538\,
            I => \N__39527\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__39535\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__9563\ : Odrv4
    port map (
            O => \N__39532\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__9562\ : Odrv4
    port map (
            O => \N__39527\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__9561\ : InMux
    port map (
            O => \N__39520\,
            I => \N__39517\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__39517\,
            I => \N__39514\
        );

    \I__9559\ : Span4Mux_s2_v
    port map (
            O => \N__39514\,
            I => \N__39511\
        );

    \I__9558\ : Odrv4
    port map (
            O => \N__39511\,
            I => \N_921_0\
        );

    \I__9557\ : InMux
    port map (
            O => \N__39508\,
            I => \N__39502\
        );

    \I__9556\ : CascadeMux
    port map (
            O => \N__39507\,
            I => \N__39499\
        );

    \I__9555\ : InMux
    port map (
            O => \N__39506\,
            I => \N__39496\
        );

    \I__9554\ : InMux
    port map (
            O => \N__39505\,
            I => \N__39493\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__39502\,
            I => \N__39489\
        );

    \I__9552\ : InMux
    port map (
            O => \N__39499\,
            I => \N__39486\
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__39496\,
            I => \N__39482\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__39493\,
            I => \N__39479\
        );

    \I__9549\ : InMux
    port map (
            O => \N__39492\,
            I => \N__39476\
        );

    \I__9548\ : Span4Mux_h
    port map (
            O => \N__39489\,
            I => \N__39473\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__39486\,
            I => \N__39470\
        );

    \I__9546\ : InMux
    port map (
            O => \N__39485\,
            I => \N__39467\
        );

    \I__9545\ : Span4Mux_v
    port map (
            O => \N__39482\,
            I => \N__39462\
        );

    \I__9544\ : Span4Mux_v
    port map (
            O => \N__39479\,
            I => \N__39462\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__39476\,
            I => \N__39456\
        );

    \I__9542\ : Span4Mux_v
    port map (
            O => \N__39473\,
            I => \N__39449\
        );

    \I__9541\ : Span4Mux_h
    port map (
            O => \N__39470\,
            I => \N__39449\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__39467\,
            I => \N__39449\
        );

    \I__9539\ : Sp12to4
    port map (
            O => \N__39462\,
            I => \N__39446\
        );

    \I__9538\ : InMux
    port map (
            O => \N__39461\,
            I => \N__39443\
        );

    \I__9537\ : InMux
    port map (
            O => \N__39460\,
            I => \N__39440\
        );

    \I__9536\ : InMux
    port map (
            O => \N__39459\,
            I => \N__39437\
        );

    \I__9535\ : Span4Mux_h
    port map (
            O => \N__39456\,
            I => \N__39434\
        );

    \I__9534\ : Span4Mux_h
    port map (
            O => \N__39449\,
            I => \N__39431\
        );

    \I__9533\ : Span12Mux_h
    port map (
            O => \N__39446\,
            I => \N__39422\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__39443\,
            I => \N__39422\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__39440\,
            I => \N__39422\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__39437\,
            I => \N__39422\
        );

    \I__9529\ : Odrv4
    port map (
            O => \N__39434\,
            I => \N_842_0\
        );

    \I__9528\ : Odrv4
    port map (
            O => \N__39431\,
            I => \N_842_0\
        );

    \I__9527\ : Odrv12
    port map (
            O => \N__39422\,
            I => \N_842_0\
        );

    \I__9526\ : InMux
    port map (
            O => \N__39415\,
            I => \N__39412\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__39412\,
            I => \N__39409\
        );

    \I__9524\ : Odrv12
    port map (
            O => \N__39409\,
            I => \M_this_status_flags_qZ0Z_7\
        );

    \I__9523\ : InMux
    port map (
            O => \N__39406\,
            I => \N__39403\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__39403\,
            I => \N__39400\
        );

    \I__9521\ : Span4Mux_h
    port map (
            O => \N__39400\,
            I => \N__39397\
        );

    \I__9520\ : Odrv4
    port map (
            O => \N__39397\,
            I => \M_this_map_address_qc_3_1\
        );

    \I__9519\ : InMux
    port map (
            O => \N__39394\,
            I => \N__39391\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__39391\,
            I => \un1_M_this_map_address_q_cry_0_c_RNOZ0\
        );

    \I__9517\ : CascadeMux
    port map (
            O => \N__39388\,
            I => \N__39385\
        );

    \I__9516\ : CascadeBuf
    port map (
            O => \N__39385\,
            I => \N__39382\
        );

    \I__9515\ : CascadeMux
    port map (
            O => \N__39382\,
            I => \N__39378\
        );

    \I__9514\ : InMux
    port map (
            O => \N__39381\,
            I => \N__39374\
        );

    \I__9513\ : InMux
    port map (
            O => \N__39378\,
            I => \N__39371\
        );

    \I__9512\ : CascadeMux
    port map (
            O => \N__39377\,
            I => \N__39368\
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__39374\,
            I => \N__39365\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__39371\,
            I => \N__39361\
        );

    \I__9509\ : InMux
    port map (
            O => \N__39368\,
            I => \N__39358\
        );

    \I__9508\ : Span4Mux_h
    port map (
            O => \N__39365\,
            I => \N__39355\
        );

    \I__9507\ : InMux
    port map (
            O => \N__39364\,
            I => \N__39352\
        );

    \I__9506\ : Span12Mux_s10_v
    port map (
            O => \N__39361\,
            I => \N__39349\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__39358\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__9504\ : Odrv4
    port map (
            O => \N__39355\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__39352\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__9502\ : Odrv12
    port map (
            O => \N__39349\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__9501\ : InMux
    port map (
            O => \N__39340\,
            I => \N__39337\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__39337\,
            I => \un1_M_this_map_address_q_cry_0_THRU_CO\
        );

    \I__9499\ : InMux
    port map (
            O => \N__39334\,
            I => \un1_M_this_map_address_q_cry_0\
        );

    \I__9498\ : CascadeMux
    port map (
            O => \N__39331\,
            I => \N__39328\
        );

    \I__9497\ : CascadeBuf
    port map (
            O => \N__39328\,
            I => \N__39325\
        );

    \I__9496\ : CascadeMux
    port map (
            O => \N__39325\,
            I => \N__39322\
        );

    \I__9495\ : InMux
    port map (
            O => \N__39322\,
            I => \N__39319\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__39319\,
            I => \N__39314\
        );

    \I__9493\ : InMux
    port map (
            O => \N__39318\,
            I => \N__39311\
        );

    \I__9492\ : InMux
    port map (
            O => \N__39317\,
            I => \N__39308\
        );

    \I__9491\ : Span12Mux_s9_h
    port map (
            O => \N__39314\,
            I => \N__39305\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__39311\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__39308\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__9488\ : Odrv12
    port map (
            O => \N__39305\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__9487\ : InMux
    port map (
            O => \N__39298\,
            I => \N__39295\
        );

    \I__9486\ : LocalMux
    port map (
            O => \N__39295\,
            I => \M_this_map_address_q_RNO_1Z0Z_2\
        );

    \I__9485\ : InMux
    port map (
            O => \N__39292\,
            I => \un1_M_this_map_address_q_cry_1\
        );

    \I__9484\ : CascadeMux
    port map (
            O => \N__39289\,
            I => \N__39286\
        );

    \I__9483\ : CascadeBuf
    port map (
            O => \N__39286\,
            I => \N__39283\
        );

    \I__9482\ : CascadeMux
    port map (
            O => \N__39283\,
            I => \N__39280\
        );

    \I__9481\ : InMux
    port map (
            O => \N__39280\,
            I => \N__39277\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__39277\,
            I => \N__39274\
        );

    \I__9479\ : Span4Mux_v
    port map (
            O => \N__39274\,
            I => \N__39269\
        );

    \I__9478\ : InMux
    port map (
            O => \N__39273\,
            I => \N__39266\
        );

    \I__9477\ : InMux
    port map (
            O => \N__39272\,
            I => \N__39263\
        );

    \I__9476\ : Span4Mux_v
    port map (
            O => \N__39269\,
            I => \N__39260\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__39266\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__39263\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__9473\ : Odrv4
    port map (
            O => \N__39260\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__9472\ : InMux
    port map (
            O => \N__39253\,
            I => \N__39250\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__39250\,
            I => \M_this_map_address_q_RNO_1Z0Z_3\
        );

    \I__9470\ : InMux
    port map (
            O => \N__39247\,
            I => \un1_M_this_map_address_q_cry_2\
        );

    \I__9469\ : CascadeMux
    port map (
            O => \N__39244\,
            I => \N__39241\
        );

    \I__9468\ : CascadeBuf
    port map (
            O => \N__39241\,
            I => \N__39238\
        );

    \I__9467\ : CascadeMux
    port map (
            O => \N__39238\,
            I => \N__39235\
        );

    \I__9466\ : InMux
    port map (
            O => \N__39235\,
            I => \N__39232\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__39232\,
            I => \N__39229\
        );

    \I__9464\ : Span4Mux_v
    port map (
            O => \N__39229\,
            I => \N__39224\
        );

    \I__9463\ : InMux
    port map (
            O => \N__39228\,
            I => \N__39221\
        );

    \I__9462\ : InMux
    port map (
            O => \N__39227\,
            I => \N__39218\
        );

    \I__9461\ : Span4Mux_v
    port map (
            O => \N__39224\,
            I => \N__39215\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__39221\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__39218\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__9458\ : Odrv4
    port map (
            O => \N__39215\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__9457\ : InMux
    port map (
            O => \N__39208\,
            I => \N__39205\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__39205\,
            I => \M_this_map_address_q_RNO_1Z0Z_4\
        );

    \I__9455\ : InMux
    port map (
            O => \N__39202\,
            I => \un1_M_this_map_address_q_cry_3\
        );

    \I__9454\ : InMux
    port map (
            O => \N__39199\,
            I => \N__39195\
        );

    \I__9453\ : InMux
    port map (
            O => \N__39198\,
            I => \N__39192\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__39195\,
            I => \un1_M_this_state_q_7_i_0_a3_0_0\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__39192\,
            I => \un1_M_this_state_q_7_i_0_a3_0_0\
        );

    \I__9450\ : InMux
    port map (
            O => \N__39187\,
            I => \un1_M_this_map_address_q_cry_4\
        );

    \I__9449\ : CEMux
    port map (
            O => \N__39184\,
            I => \N__39181\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__39181\,
            I => \N__39177\
        );

    \I__9447\ : CEMux
    port map (
            O => \N__39180\,
            I => \N__39174\
        );

    \I__9446\ : Span4Mux_h
    port map (
            O => \N__39177\,
            I => \N__39169\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__39174\,
            I => \N__39169\
        );

    \I__9444\ : Span4Mux_v
    port map (
            O => \N__39169\,
            I => \N__39166\
        );

    \I__9443\ : Odrv4
    port map (
            O => \N__39166\,
            I => \this_spr_ram.mem_WE_10\
        );

    \I__9442\ : InMux
    port map (
            O => \N__39163\,
            I => \N__39160\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__39160\,
            I => \N__39157\
        );

    \I__9440\ : Odrv4
    port map (
            O => \N__39157\,
            I => \this_spr_ram.mem_out_bus4_0\
        );

    \I__9439\ : InMux
    port map (
            O => \N__39154\,
            I => \N__39151\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__39151\,
            I => \N__39148\
        );

    \I__9437\ : Sp12to4
    port map (
            O => \N__39148\,
            I => \N__39145\
        );

    \I__9436\ : Span12Mux_v
    port map (
            O => \N__39145\,
            I => \N__39142\
        );

    \I__9435\ : Odrv12
    port map (
            O => \N__39142\,
            I => \this_spr_ram.mem_out_bus0_0\
        );

    \I__9434\ : InMux
    port map (
            O => \N__39139\,
            I => \N__39136\
        );

    \I__9433\ : LocalMux
    port map (
            O => \N__39136\,
            I => \this_spr_ram.mem_mem_0_0_RNIK6VFZ0\
        );

    \I__9432\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39130\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__39130\,
            I => \N__39127\
        );

    \I__9430\ : Span4Mux_v
    port map (
            O => \N__39127\,
            I => \N__39124\
        );

    \I__9429\ : Odrv4
    port map (
            O => \N__39124\,
            I => \this_spr_ram.mem_out_bus2_1\
        );

    \I__9428\ : InMux
    port map (
            O => \N__39121\,
            I => \N__39118\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__39118\,
            I => \N__39114\
        );

    \I__9426\ : InMux
    port map (
            O => \N__39117\,
            I => \N__39101\
        );

    \I__9425\ : Span4Mux_v
    port map (
            O => \N__39114\,
            I => \N__39094\
        );

    \I__9424\ : InMux
    port map (
            O => \N__39113\,
            I => \N__39081\
        );

    \I__9423\ : InMux
    port map (
            O => \N__39112\,
            I => \N__39081\
        );

    \I__9422\ : InMux
    port map (
            O => \N__39111\,
            I => \N__39081\
        );

    \I__9421\ : InMux
    port map (
            O => \N__39110\,
            I => \N__39081\
        );

    \I__9420\ : InMux
    port map (
            O => \N__39109\,
            I => \N__39081\
        );

    \I__9419\ : InMux
    port map (
            O => \N__39108\,
            I => \N__39081\
        );

    \I__9418\ : InMux
    port map (
            O => \N__39107\,
            I => \N__39076\
        );

    \I__9417\ : InMux
    port map (
            O => \N__39106\,
            I => \N__39076\
        );

    \I__9416\ : InMux
    port map (
            O => \N__39105\,
            I => \N__39073\
        );

    \I__9415\ : InMux
    port map (
            O => \N__39104\,
            I => \N__39070\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__39101\,
            I => \N__39067\
        );

    \I__9413\ : InMux
    port map (
            O => \N__39100\,
            I => \N__39062\
        );

    \I__9412\ : InMux
    port map (
            O => \N__39099\,
            I => \N__39062\
        );

    \I__9411\ : InMux
    port map (
            O => \N__39098\,
            I => \N__39059\
        );

    \I__9410\ : InMux
    port map (
            O => \N__39097\,
            I => \N__39056\
        );

    \I__9409\ : Span4Mux_v
    port map (
            O => \N__39094\,
            I => \N__39051\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__39081\,
            I => \N__39051\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__39076\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9406\ : LocalMux
    port map (
            O => \N__39073\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__39070\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9404\ : Odrv4
    port map (
            O => \N__39067\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__39062\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__39059\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__39056\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9400\ : Odrv4
    port map (
            O => \N__39051\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9399\ : InMux
    port map (
            O => \N__39034\,
            I => \N__39031\
        );

    \I__9398\ : LocalMux
    port map (
            O => \N__39031\,
            I => \N__39028\
        );

    \I__9397\ : Span4Mux_v
    port map (
            O => \N__39028\,
            I => \N__39025\
        );

    \I__9396\ : Span4Mux_v
    port map (
            O => \N__39025\,
            I => \N__39022\
        );

    \I__9395\ : Odrv4
    port map (
            O => \N__39022\,
            I => \this_spr_ram.mem_out_bus6_1\
        );

    \I__9394\ : InMux
    port map (
            O => \N__39019\,
            I => \N__39016\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__39016\,
            I => \N__39013\
        );

    \I__9392\ : Odrv4
    port map (
            O => \N__39013\,
            I => \this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0\
        );

    \I__9391\ : InMux
    port map (
            O => \N__39010\,
            I => \N__39007\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__39007\,
            I => \N__39003\
        );

    \I__9389\ : InMux
    port map (
            O => \N__39006\,
            I => \N__39000\
        );

    \I__9388\ : Span4Mux_v
    port map (
            O => \N__39003\,
            I => \N__38995\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__39000\,
            I => \N__38995\
        );

    \I__9386\ : Span4Mux_h
    port map (
            O => \N__38995\,
            I => \N__38992\
        );

    \I__9385\ : Sp12to4
    port map (
            O => \N__38992\,
            I => \N__38989\
        );

    \I__9384\ : Span12Mux_v
    port map (
            O => \N__38989\,
            I => \N__38986\
        );

    \I__9383\ : Odrv12
    port map (
            O => \N__38986\,
            I => \M_this_map_ram_read_data_7\
        );

    \I__9382\ : IoInMux
    port map (
            O => \N__38983\,
            I => \N__38980\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__38980\,
            I => \N__38977\
        );

    \I__9380\ : IoSpan4Mux
    port map (
            O => \N__38977\,
            I => \N__38974\
        );

    \I__9379\ : IoSpan4Mux
    port map (
            O => \N__38974\,
            I => \N__38971\
        );

    \I__9378\ : Span4Mux_s3_h
    port map (
            O => \N__38971\,
            I => \N__38968\
        );

    \I__9377\ : Span4Mux_h
    port map (
            O => \N__38968\,
            I => \N__38965\
        );

    \I__9376\ : Odrv4
    port map (
            O => \N__38965\,
            I => \IO_port_data_write_i_m2_i_m2_7\
        );

    \I__9375\ : CEMux
    port map (
            O => \N__38962\,
            I => \N__38958\
        );

    \I__9374\ : CEMux
    port map (
            O => \N__38961\,
            I => \N__38955\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__38958\,
            I => \N__38950\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__38955\,
            I => \N__38950\
        );

    \I__9371\ : Span4Mux_v
    port map (
            O => \N__38950\,
            I => \N__38947\
        );

    \I__9370\ : Odrv4
    port map (
            O => \N__38947\,
            I => \this_spr_ram.mem_WE_6\
        );

    \I__9369\ : CEMux
    port map (
            O => \N__38944\,
            I => \N__38940\
        );

    \I__9368\ : CEMux
    port map (
            O => \N__38943\,
            I => \N__38937\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__38940\,
            I => \N__38932\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__38937\,
            I => \N__38932\
        );

    \I__9365\ : Span4Mux_v
    port map (
            O => \N__38932\,
            I => \N__38929\
        );

    \I__9364\ : Odrv4
    port map (
            O => \N__38929\,
            I => \this_spr_ram.mem_WE_4\
        );

    \I__9363\ : InMux
    port map (
            O => \N__38926\,
            I => \N__38914\
        );

    \I__9362\ : InMux
    port map (
            O => \N__38925\,
            I => \N__38914\
        );

    \I__9361\ : InMux
    port map (
            O => \N__38924\,
            I => \N__38914\
        );

    \I__9360\ : InMux
    port map (
            O => \N__38923\,
            I => \N__38911\
        );

    \I__9359\ : InMux
    port map (
            O => \N__38922\,
            I => \N__38908\
        );

    \I__9358\ : InMux
    port map (
            O => \N__38921\,
            I => \N__38905\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__38914\,
            I => \N__38895\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__38911\,
            I => \N__38895\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__38908\,
            I => \N__38895\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__38905\,
            I => \N__38892\
        );

    \I__9353\ : InMux
    port map (
            O => \N__38904\,
            I => \N__38887\
        );

    \I__9352\ : InMux
    port map (
            O => \N__38903\,
            I => \N__38887\
        );

    \I__9351\ : InMux
    port map (
            O => \N__38902\,
            I => \N__38884\
        );

    \I__9350\ : Span4Mux_v
    port map (
            O => \N__38895\,
            I => \N__38881\
        );

    \I__9349\ : Span4Mux_h
    port map (
            O => \N__38892\,
            I => \N__38878\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__38887\,
            I => \N__38875\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__38884\,
            I => \M_this_spr_address_qZ0Z_12\
        );

    \I__9346\ : Odrv4
    port map (
            O => \N__38881\,
            I => \M_this_spr_address_qZ0Z_12\
        );

    \I__9345\ : Odrv4
    port map (
            O => \N__38878\,
            I => \M_this_spr_address_qZ0Z_12\
        );

    \I__9344\ : Odrv12
    port map (
            O => \N__38875\,
            I => \M_this_spr_address_qZ0Z_12\
        );

    \I__9343\ : CascadeMux
    port map (
            O => \N__38866\,
            I => \N__38862\
        );

    \I__9342\ : InMux
    port map (
            O => \N__38865\,
            I => \N__38855\
        );

    \I__9341\ : InMux
    port map (
            O => \N__38862\,
            I => \N__38848\
        );

    \I__9340\ : InMux
    port map (
            O => \N__38861\,
            I => \N__38848\
        );

    \I__9339\ : InMux
    port map (
            O => \N__38860\,
            I => \N__38848\
        );

    \I__9338\ : InMux
    port map (
            O => \N__38859\,
            I => \N__38843\
        );

    \I__9337\ : CascadeMux
    port map (
            O => \N__38858\,
            I => \N__38840\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__38855\,
            I => \N__38836\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__38848\,
            I => \N__38833\
        );

    \I__9334\ : InMux
    port map (
            O => \N__38847\,
            I => \N__38830\
        );

    \I__9333\ : InMux
    port map (
            O => \N__38846\,
            I => \N__38827\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__38843\,
            I => \N__38824\
        );

    \I__9331\ : InMux
    port map (
            O => \N__38840\,
            I => \N__38819\
        );

    \I__9330\ : InMux
    port map (
            O => \N__38839\,
            I => \N__38819\
        );

    \I__9329\ : Span4Mux_v
    port map (
            O => \N__38836\,
            I => \N__38814\
        );

    \I__9328\ : Span4Mux_v
    port map (
            O => \N__38833\,
            I => \N__38814\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__38830\,
            I => \N__38811\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__38827\,
            I => \N__38802\
        );

    \I__9325\ : Span4Mux_v
    port map (
            O => \N__38824\,
            I => \N__38802\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__38819\,
            I => \N__38802\
        );

    \I__9323\ : Span4Mux_h
    port map (
            O => \N__38814\,
            I => \N__38802\
        );

    \I__9322\ : Odrv4
    port map (
            O => \N__38811\,
            I => \M_this_spr_address_qZ0Z_11\
        );

    \I__9321\ : Odrv4
    port map (
            O => \N__38802\,
            I => \M_this_spr_address_qZ0Z_11\
        );

    \I__9320\ : CascadeMux
    port map (
            O => \N__38797\,
            I => \N__38790\
        );

    \I__9319\ : CascadeMux
    port map (
            O => \N__38796\,
            I => \N__38786\
        );

    \I__9318\ : CascadeMux
    port map (
            O => \N__38795\,
            I => \N__38783\
        );

    \I__9317\ : CascadeMux
    port map (
            O => \N__38794\,
            I => \N__38780\
        );

    \I__9316\ : CascadeMux
    port map (
            O => \N__38793\,
            I => \N__38777\
        );

    \I__9315\ : InMux
    port map (
            O => \N__38790\,
            I => \N__38769\
        );

    \I__9314\ : InMux
    port map (
            O => \N__38789\,
            I => \N__38769\
        );

    \I__9313\ : InMux
    port map (
            O => \N__38786\,
            I => \N__38769\
        );

    \I__9312\ : InMux
    port map (
            O => \N__38783\,
            I => \N__38766\
        );

    \I__9311\ : InMux
    port map (
            O => \N__38780\,
            I => \N__38763\
        );

    \I__9310\ : InMux
    port map (
            O => \N__38777\,
            I => \N__38760\
        );

    \I__9309\ : CascadeMux
    port map (
            O => \N__38776\,
            I => \N__38756\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__38769\,
            I => \N__38748\
        );

    \I__9307\ : LocalMux
    port map (
            O => \N__38766\,
            I => \N__38748\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__38763\,
            I => \N__38748\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__38760\,
            I => \N__38745\
        );

    \I__9304\ : InMux
    port map (
            O => \N__38759\,
            I => \N__38740\
        );

    \I__9303\ : InMux
    port map (
            O => \N__38756\,
            I => \N__38740\
        );

    \I__9302\ : InMux
    port map (
            O => \N__38755\,
            I => \N__38737\
        );

    \I__9301\ : Span4Mux_v
    port map (
            O => \N__38748\,
            I => \N__38734\
        );

    \I__9300\ : Span4Mux_h
    port map (
            O => \N__38745\,
            I => \N__38731\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__38740\,
            I => \N__38728\
        );

    \I__9298\ : LocalMux
    port map (
            O => \N__38737\,
            I => \M_this_spr_address_qZ0Z_13\
        );

    \I__9297\ : Odrv4
    port map (
            O => \N__38734\,
            I => \M_this_spr_address_qZ0Z_13\
        );

    \I__9296\ : Odrv4
    port map (
            O => \N__38731\,
            I => \M_this_spr_address_qZ0Z_13\
        );

    \I__9295\ : Odrv4
    port map (
            O => \N__38728\,
            I => \M_this_spr_address_qZ0Z_13\
        );

    \I__9294\ : InMux
    port map (
            O => \N__38719\,
            I => \N__38713\
        );

    \I__9293\ : InMux
    port map (
            O => \N__38718\,
            I => \N__38710\
        );

    \I__9292\ : InMux
    port map (
            O => \N__38717\,
            I => \N__38704\
        );

    \I__9291\ : InMux
    port map (
            O => \N__38716\,
            I => \N__38704\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__38713\,
            I => \N__38698\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__38710\,
            I => \N__38695\
        );

    \I__9288\ : InMux
    port map (
            O => \N__38709\,
            I => \N__38692\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__38704\,
            I => \N__38689\
        );

    \I__9286\ : InMux
    port map (
            O => \N__38703\,
            I => \N__38682\
        );

    \I__9285\ : InMux
    port map (
            O => \N__38702\,
            I => \N__38682\
        );

    \I__9284\ : InMux
    port map (
            O => \N__38701\,
            I => \N__38682\
        );

    \I__9283\ : Span4Mux_h
    port map (
            O => \N__38698\,
            I => \N__38679\
        );

    \I__9282\ : Span4Mux_h
    port map (
            O => \N__38695\,
            I => \N__38674\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__38692\,
            I => \N__38674\
        );

    \I__9280\ : Span4Mux_h
    port map (
            O => \N__38689\,
            I => \N__38671\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__38682\,
            I => \N__38668\
        );

    \I__9278\ : Span4Mux_v
    port map (
            O => \N__38679\,
            I => \N__38665\
        );

    \I__9277\ : Span4Mux_v
    port map (
            O => \N__38674\,
            I => \N__38662\
        );

    \I__9276\ : Span4Mux_v
    port map (
            O => \N__38671\,
            I => \N__38657\
        );

    \I__9275\ : Span4Mux_h
    port map (
            O => \N__38668\,
            I => \N__38657\
        );

    \I__9274\ : Odrv4
    port map (
            O => \N__38665\,
            I => \M_this_spr_ram_write_en_0_i_1_0_0\
        );

    \I__9273\ : Odrv4
    port map (
            O => \N__38662\,
            I => \M_this_spr_ram_write_en_0_i_1_0_0\
        );

    \I__9272\ : Odrv4
    port map (
            O => \N__38657\,
            I => \M_this_spr_ram_write_en_0_i_1_0_0\
        );

    \I__9271\ : CEMux
    port map (
            O => \N__38650\,
            I => \N__38647\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__38647\,
            I => \N__38643\
        );

    \I__9269\ : CEMux
    port map (
            O => \N__38646\,
            I => \N__38640\
        );

    \I__9268\ : Sp12to4
    port map (
            O => \N__38643\,
            I => \N__38637\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__38640\,
            I => \N__38634\
        );

    \I__9266\ : Span12Mux_v
    port map (
            O => \N__38637\,
            I => \N__38631\
        );

    \I__9265\ : Span4Mux_v
    port map (
            O => \N__38634\,
            I => \N__38628\
        );

    \I__9264\ : Span12Mux_h
    port map (
            O => \N__38631\,
            I => \N__38625\
        );

    \I__9263\ : Span4Mux_v
    port map (
            O => \N__38628\,
            I => \N__38622\
        );

    \I__9262\ : Odrv12
    port map (
            O => \N__38625\,
            I => \this_spr_ram.mem_WE_2\
        );

    \I__9261\ : Odrv4
    port map (
            O => \N__38622\,
            I => \this_spr_ram.mem_WE_2\
        );

    \I__9260\ : InMux
    port map (
            O => \N__38617\,
            I => \N__38614\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__38614\,
            I => \N_1066\
        );

    \I__9258\ : CascadeMux
    port map (
            O => \N__38611\,
            I => \M_this_map_address_qc_6_0_cascade_\
        );

    \I__9257\ : InMux
    port map (
            O => \N__38608\,
            I => \N__38602\
        );

    \I__9256\ : InMux
    port map (
            O => \N__38607\,
            I => \N__38599\
        );

    \I__9255\ : InMux
    port map (
            O => \N__38606\,
            I => \N__38592\
        );

    \I__9254\ : InMux
    port map (
            O => \N__38605\,
            I => \N__38589\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__38602\,
            I => \N__38581\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__38599\,
            I => \N__38581\
        );

    \I__9251\ : InMux
    port map (
            O => \N__38598\,
            I => \N__38578\
        );

    \I__9250\ : InMux
    port map (
            O => \N__38597\,
            I => \N__38571\
        );

    \I__9249\ : InMux
    port map (
            O => \N__38596\,
            I => \N__38571\
        );

    \I__9248\ : InMux
    port map (
            O => \N__38595\,
            I => \N__38571\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__38592\,
            I => \N__38566\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__38589\,
            I => \N__38566\
        );

    \I__9245\ : InMux
    port map (
            O => \N__38588\,
            I => \N__38563\
        );

    \I__9244\ : InMux
    port map (
            O => \N__38587\,
            I => \N__38560\
        );

    \I__9243\ : InMux
    port map (
            O => \N__38586\,
            I => \N__38557\
        );

    \I__9242\ : Span4Mux_v
    port map (
            O => \N__38581\,
            I => \N__38550\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__38578\,
            I => \N__38550\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__38571\,
            I => \N__38550\
        );

    \I__9239\ : Span4Mux_v
    port map (
            O => \N__38566\,
            I => \N__38545\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__38563\,
            I => \N__38545\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__38560\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__9236\ : LocalMux
    port map (
            O => \N__38557\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__9235\ : Odrv4
    port map (
            O => \N__38550\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__9234\ : Odrv4
    port map (
            O => \N__38545\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__9233\ : InMux
    port map (
            O => \N__38536\,
            I => \N__38527\
        );

    \I__9232\ : InMux
    port map (
            O => \N__38535\,
            I => \N__38527\
        );

    \I__9231\ : InMux
    port map (
            O => \N__38534\,
            I => \N__38524\
        );

    \I__9230\ : InMux
    port map (
            O => \N__38533\,
            I => \N__38519\
        );

    \I__9229\ : InMux
    port map (
            O => \N__38532\,
            I => \N__38519\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__38527\,
            I => \N__38514\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__38524\,
            I => \N__38514\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__38519\,
            I => \N__38511\
        );

    \I__9225\ : Span4Mux_h
    port map (
            O => \N__38514\,
            I => \N__38508\
        );

    \I__9224\ : Odrv12
    port map (
            O => \N__38511\,
            I => \N_794_0\
        );

    \I__9223\ : Odrv4
    port map (
            O => \N__38508\,
            I => \N_794_0\
        );

    \I__9222\ : InMux
    port map (
            O => \N__38503\,
            I => \N__38500\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__38500\,
            I => \N__38497\
        );

    \I__9220\ : Odrv4
    port map (
            O => \N__38497\,
            I => \M_this_map_address_qc_4_0\
        );

    \I__9219\ : InMux
    port map (
            O => \N__38494\,
            I => \N__38491\
        );

    \I__9218\ : LocalMux
    port map (
            O => \N__38491\,
            I => \N__38488\
        );

    \I__9217\ : Span4Mux_h
    port map (
            O => \N__38488\,
            I => \N__38485\
        );

    \I__9216\ : Odrv4
    port map (
            O => \N__38485\,
            I => \N_918_0\
        );

    \I__9215\ : InMux
    port map (
            O => \N__38482\,
            I => \N__38479\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__38479\,
            I => \N__38475\
        );

    \I__9213\ : InMux
    port map (
            O => \N__38478\,
            I => \N__38472\
        );

    \I__9212\ : Span12Mux_v
    port map (
            O => \N__38475\,
            I => \N__38469\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__38472\,
            I => \N__38466\
        );

    \I__9210\ : Odrv12
    port map (
            O => \N__38469\,
            I => m5_i_a2_i_o3_i_a3
        );

    \I__9209\ : Odrv12
    port map (
            O => \N__38466\,
            I => m5_i_a2_i_o3_i_a3
        );

    \I__9208\ : IoInMux
    port map (
            O => \N__38461\,
            I => \N__38458\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__38458\,
            I => \N__38454\
        );

    \I__9206\ : IoInMux
    port map (
            O => \N__38457\,
            I => \N__38451\
        );

    \I__9205\ : IoSpan4Mux
    port map (
            O => \N__38454\,
            I => \N__38446\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__38451\,
            I => \N__38446\
        );

    \I__9203\ : IoSpan4Mux
    port map (
            O => \N__38446\,
            I => \N__38442\
        );

    \I__9202\ : IoInMux
    port map (
            O => \N__38445\,
            I => \N__38439\
        );

    \I__9201\ : IoSpan4Mux
    port map (
            O => \N__38442\,
            I => \N__38432\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__38439\,
            I => \N__38432\
        );

    \I__9199\ : IoInMux
    port map (
            O => \N__38438\,
            I => \N__38428\
        );

    \I__9198\ : IoInMux
    port map (
            O => \N__38437\,
            I => \N__38425\
        );

    \I__9197\ : IoSpan4Mux
    port map (
            O => \N__38432\,
            I => \N__38422\
        );

    \I__9196\ : IoInMux
    port map (
            O => \N__38431\,
            I => \N__38419\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__38428\,
            I => \N__38414\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__38425\,
            I => \N__38414\
        );

    \I__9193\ : IoSpan4Mux
    port map (
            O => \N__38422\,
            I => \N__38408\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__38419\,
            I => \N__38408\
        );

    \I__9191\ : IoSpan4Mux
    port map (
            O => \N__38414\,
            I => \N__38405\
        );

    \I__9190\ : IoInMux
    port map (
            O => \N__38413\,
            I => \N__38402\
        );

    \I__9189\ : IoSpan4Mux
    port map (
            O => \N__38408\,
            I => \N__38398\
        );

    \I__9188\ : IoSpan4Mux
    port map (
            O => \N__38405\,
            I => \N__38395\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__38402\,
            I => \N__38392\
        );

    \I__9186\ : IoInMux
    port map (
            O => \N__38401\,
            I => \N__38389\
        );

    \I__9185\ : Span4Mux_s1_h
    port map (
            O => \N__38398\,
            I => \N__38386\
        );

    \I__9184\ : IoSpan4Mux
    port map (
            O => \N__38395\,
            I => \N__38383\
        );

    \I__9183\ : IoSpan4Mux
    port map (
            O => \N__38392\,
            I => \N__38380\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__38389\,
            I => \N__38377\
        );

    \I__9181\ : Span4Mux_h
    port map (
            O => \N__38386\,
            I => \N__38368\
        );

    \I__9180\ : Span4Mux_s2_v
    port map (
            O => \N__38383\,
            I => \N__38368\
        );

    \I__9179\ : Span4Mux_s2_v
    port map (
            O => \N__38380\,
            I => \N__38368\
        );

    \I__9178\ : Span4Mux_s2_v
    port map (
            O => \N__38377\,
            I => \N__38368\
        );

    \I__9177\ : Odrv4
    port map (
            O => \N__38368\,
            I => \N_1048_i_0\
        );

    \I__9176\ : CEMux
    port map (
            O => \N__38365\,
            I => \N__38361\
        );

    \I__9175\ : CEMux
    port map (
            O => \N__38364\,
            I => \N__38358\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__38361\,
            I => \N__38353\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__38358\,
            I => \N__38353\
        );

    \I__9172\ : Span4Mux_v
    port map (
            O => \N__38353\,
            I => \N__38350\
        );

    \I__9171\ : Odrv4
    port map (
            O => \N__38350\,
            I => \this_spr_ram.mem_WE_12\
        );

    \I__9170\ : CEMux
    port map (
            O => \N__38347\,
            I => \N__38343\
        );

    \I__9169\ : CEMux
    port map (
            O => \N__38346\,
            I => \N__38340\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__38343\,
            I => \N__38337\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__38340\,
            I => \N__38334\
        );

    \I__9166\ : Span4Mux_v
    port map (
            O => \N__38337\,
            I => \N__38331\
        );

    \I__9165\ : Span4Mux_h
    port map (
            O => \N__38334\,
            I => \N__38328\
        );

    \I__9164\ : Odrv4
    port map (
            O => \N__38331\,
            I => \this_spr_ram.mem_WE_8\
        );

    \I__9163\ : Odrv4
    port map (
            O => \N__38328\,
            I => \this_spr_ram.mem_WE_8\
        );

    \I__9162\ : CEMux
    port map (
            O => \N__38323\,
            I => \N__38319\
        );

    \I__9161\ : CEMux
    port map (
            O => \N__38322\,
            I => \N__38316\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__38319\,
            I => \N__38313\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__38316\,
            I => \N__38310\
        );

    \I__9158\ : Span4Mux_h
    port map (
            O => \N__38313\,
            I => \N__38307\
        );

    \I__9157\ : Span4Mux_h
    port map (
            O => \N__38310\,
            I => \N__38304\
        );

    \I__9156\ : Span4Mux_v
    port map (
            O => \N__38307\,
            I => \N__38301\
        );

    \I__9155\ : Span4Mux_v
    port map (
            O => \N__38304\,
            I => \N__38298\
        );

    \I__9154\ : Span4Mux_v
    port map (
            O => \N__38301\,
            I => \N__38295\
        );

    \I__9153\ : Span4Mux_v
    port map (
            O => \N__38298\,
            I => \N__38292\
        );

    \I__9152\ : Odrv4
    port map (
            O => \N__38295\,
            I => \this_spr_ram.mem_WE_14\
        );

    \I__9151\ : Odrv4
    port map (
            O => \N__38292\,
            I => \this_spr_ram.mem_WE_14\
        );

    \I__9150\ : InMux
    port map (
            O => \N__38287\,
            I => \N__38282\
        );

    \I__9149\ : InMux
    port map (
            O => \N__38286\,
            I => \N__38277\
        );

    \I__9148\ : InMux
    port map (
            O => \N__38285\,
            I => \N__38277\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__38282\,
            I => \N__38270\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__38277\,
            I => \N__38270\
        );

    \I__9145\ : InMux
    port map (
            O => \N__38276\,
            I => \N__38265\
        );

    \I__9144\ : InMux
    port map (
            O => \N__38275\,
            I => \N__38265\
        );

    \I__9143\ : Odrv4
    port map (
            O => \N__38270\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__38265\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__9141\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38257\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__38257\,
            I => \this_ppu_un1_M_this_state_q_7_i_0_0_0\
        );

    \I__9139\ : CascadeMux
    port map (
            O => \N__38254\,
            I => \un1_M_this_state_q_7_i_0_a3_0_0_cascade_\
        );

    \I__9138\ : InMux
    port map (
            O => \N__38251\,
            I => \N__38248\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__38248\,
            I => \N__38245\
        );

    \I__9136\ : Span4Mux_h
    port map (
            O => \N__38245\,
            I => \N__38242\
        );

    \I__9135\ : Span4Mux_h
    port map (
            O => \N__38242\,
            I => \N__38239\
        );

    \I__9134\ : Span4Mux_h
    port map (
            O => \N__38239\,
            I => \N__38236\
        );

    \I__9133\ : Odrv4
    port map (
            O => \N__38236\,
            I => \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0\
        );

    \I__9132\ : InMux
    port map (
            O => \N__38233\,
            I => \N__38230\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__38230\,
            I => \N__38227\
        );

    \I__9130\ : Span4Mux_v
    port map (
            O => \N__38227\,
            I => \N__38223\
        );

    \I__9129\ : InMux
    port map (
            O => \N__38226\,
            I => \N__38220\
        );

    \I__9128\ : Sp12to4
    port map (
            O => \N__38223\,
            I => \N__38217\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__38220\,
            I => \N__38214\
        );

    \I__9126\ : Span12Mux_h
    port map (
            O => \N__38217\,
            I => \N__38209\
        );

    \I__9125\ : Span12Mux_v
    port map (
            O => \N__38214\,
            I => \N__38209\
        );

    \I__9124\ : Odrv12
    port map (
            O => \N__38209\,
            I => \M_this_map_ram_read_data_0\
        );

    \I__9123\ : InMux
    port map (
            O => \N__38206\,
            I => \N__38199\
        );

    \I__9122\ : InMux
    port map (
            O => \N__38205\,
            I => \N__38199\
        );

    \I__9121\ : InMux
    port map (
            O => \N__38204\,
            I => \N__38195\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__38199\,
            I => \N__38192\
        );

    \I__9119\ : InMux
    port map (
            O => \N__38198\,
            I => \N__38189\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__38195\,
            I => \N__38184\
        );

    \I__9117\ : Span4Mux_v
    port map (
            O => \N__38192\,
            I => \N__38179\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__38189\,
            I => \N__38179\
        );

    \I__9115\ : InMux
    port map (
            O => \N__38188\,
            I => \N__38169\
        );

    \I__9114\ : InMux
    port map (
            O => \N__38187\,
            I => \N__38169\
        );

    \I__9113\ : Span4Mux_v
    port map (
            O => \N__38184\,
            I => \N__38164\
        );

    \I__9112\ : Span4Mux_v
    port map (
            O => \N__38179\,
            I => \N__38164\
        );

    \I__9111\ : InMux
    port map (
            O => \N__38178\,
            I => \N__38152\
        );

    \I__9110\ : InMux
    port map (
            O => \N__38177\,
            I => \N__38152\
        );

    \I__9109\ : InMux
    port map (
            O => \N__38176\,
            I => \N__38152\
        );

    \I__9108\ : InMux
    port map (
            O => \N__38175\,
            I => \N__38152\
        );

    \I__9107\ : InMux
    port map (
            O => \N__38174\,
            I => \N__38152\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__38169\,
            I => \N__38147\
        );

    \I__9105\ : Span4Mux_h
    port map (
            O => \N__38164\,
            I => \N__38144\
        );

    \I__9104\ : InMux
    port map (
            O => \N__38163\,
            I => \N__38141\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__38152\,
            I => \N__38138\
        );

    \I__9102\ : InMux
    port map (
            O => \N__38151\,
            I => \N__38135\
        );

    \I__9101\ : InMux
    port map (
            O => \N__38150\,
            I => \N__38132\
        );

    \I__9100\ : Span4Mux_h
    port map (
            O => \N__38147\,
            I => \N__38129\
        );

    \I__9099\ : Span4Mux_h
    port map (
            O => \N__38144\,
            I => \N__38126\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__38141\,
            I => \N__38121\
        );

    \I__9097\ : Span4Mux_v
    port map (
            O => \N__38138\,
            I => \N__38121\
        );

    \I__9096\ : LocalMux
    port map (
            O => \N__38135\,
            I => \N__38114\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__38132\,
            I => \N__38114\
        );

    \I__9094\ : Span4Mux_h
    port map (
            O => \N__38129\,
            I => \N__38114\
        );

    \I__9093\ : Odrv4
    port map (
            O => \N__38126\,
            I => \this_ppu.N_785_0\
        );

    \I__9092\ : Odrv4
    port map (
            O => \N__38121\,
            I => \this_ppu.N_785_0\
        );

    \I__9091\ : Odrv4
    port map (
            O => \N__38114\,
            I => \this_ppu.N_785_0\
        );

    \I__9090\ : CascadeMux
    port map (
            O => \N__38107\,
            I => \N__38101\
        );

    \I__9089\ : CascadeMux
    port map (
            O => \N__38106\,
            I => \N__38098\
        );

    \I__9088\ : CascadeMux
    port map (
            O => \N__38105\,
            I => \N__38094\
        );

    \I__9087\ : CascadeMux
    port map (
            O => \N__38104\,
            I => \N__38091\
        );

    \I__9086\ : InMux
    port map (
            O => \N__38101\,
            I => \N__38087\
        );

    \I__9085\ : InMux
    port map (
            O => \N__38098\,
            I => \N__38084\
        );

    \I__9084\ : CascadeMux
    port map (
            O => \N__38097\,
            I => \N__38081\
        );

    \I__9083\ : InMux
    port map (
            O => \N__38094\,
            I => \N__38076\
        );

    \I__9082\ : InMux
    port map (
            O => \N__38091\,
            I => \N__38073\
        );

    \I__9081\ : CascadeMux
    port map (
            O => \N__38090\,
            I => \N__38070\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__38087\,
            I => \N__38063\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__38084\,
            I => \N__38063\
        );

    \I__9078\ : InMux
    port map (
            O => \N__38081\,
            I => \N__38060\
        );

    \I__9077\ : CascadeMux
    port map (
            O => \N__38080\,
            I => \N__38057\
        );

    \I__9076\ : CascadeMux
    port map (
            O => \N__38079\,
            I => \N__38054\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__38076\,
            I => \N__38050\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__38073\,
            I => \N__38047\
        );

    \I__9073\ : InMux
    port map (
            O => \N__38070\,
            I => \N__38044\
        );

    \I__9072\ : CascadeMux
    port map (
            O => \N__38069\,
            I => \N__38041\
        );

    \I__9071\ : CascadeMux
    port map (
            O => \N__38068\,
            I => \N__38034\
        );

    \I__9070\ : Span4Mux_v
    port map (
            O => \N__38063\,
            I => \N__38029\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__38060\,
            I => \N__38029\
        );

    \I__9068\ : InMux
    port map (
            O => \N__38057\,
            I => \N__38026\
        );

    \I__9067\ : InMux
    port map (
            O => \N__38054\,
            I => \N__38023\
        );

    \I__9066\ : CascadeMux
    port map (
            O => \N__38053\,
            I => \N__38020\
        );

    \I__9065\ : Span4Mux_v
    port map (
            O => \N__38050\,
            I => \N__38013\
        );

    \I__9064\ : Span4Mux_h
    port map (
            O => \N__38047\,
            I => \N__38013\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__38044\,
            I => \N__38013\
        );

    \I__9062\ : InMux
    port map (
            O => \N__38041\,
            I => \N__38010\
        );

    \I__9061\ : CascadeMux
    port map (
            O => \N__38040\,
            I => \N__38007\
        );

    \I__9060\ : CascadeMux
    port map (
            O => \N__38039\,
            I => \N__38004\
        );

    \I__9059\ : CascadeMux
    port map (
            O => \N__38038\,
            I => \N__38001\
        );

    \I__9058\ : CascadeMux
    port map (
            O => \N__38037\,
            I => \N__37998\
        );

    \I__9057\ : InMux
    port map (
            O => \N__38034\,
            I => \N__37994\
        );

    \I__9056\ : Span4Mux_h
    port map (
            O => \N__38029\,
            I => \N__37991\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__38026\,
            I => \N__37986\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__38023\,
            I => \N__37986\
        );

    \I__9053\ : InMux
    port map (
            O => \N__38020\,
            I => \N__37983\
        );

    \I__9052\ : Span4Mux_v
    port map (
            O => \N__38013\,
            I => \N__37978\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__38010\,
            I => \N__37978\
        );

    \I__9050\ : InMux
    port map (
            O => \N__38007\,
            I => \N__37975\
        );

    \I__9049\ : InMux
    port map (
            O => \N__38004\,
            I => \N__37972\
        );

    \I__9048\ : InMux
    port map (
            O => \N__38001\,
            I => \N__37969\
        );

    \I__9047\ : InMux
    port map (
            O => \N__37998\,
            I => \N__37966\
        );

    \I__9046\ : CascadeMux
    port map (
            O => \N__37997\,
            I => \N__37963\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__37994\,
            I => \N__37960\
        );

    \I__9044\ : Span4Mux_v
    port map (
            O => \N__37991\,
            I => \N__37957\
        );

    \I__9043\ : Span12Mux_s10_v
    port map (
            O => \N__37986\,
            I => \N__37946\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__37983\,
            I => \N__37946\
        );

    \I__9041\ : Sp12to4
    port map (
            O => \N__37978\,
            I => \N__37946\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__37975\,
            I => \N__37946\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__37972\,
            I => \N__37946\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__37969\,
            I => \N__37943\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__37966\,
            I => \N__37940\
        );

    \I__9036\ : InMux
    port map (
            O => \N__37963\,
            I => \N__37937\
        );

    \I__9035\ : Span4Mux_v
    port map (
            O => \N__37960\,
            I => \N__37934\
        );

    \I__9034\ : Sp12to4
    port map (
            O => \N__37957\,
            I => \N__37929\
        );

    \I__9033\ : Span12Mux_v
    port map (
            O => \N__37946\,
            I => \N__37929\
        );

    \I__9032\ : Span4Mux_h
    port map (
            O => \N__37943\,
            I => \N__37924\
        );

    \I__9031\ : Span4Mux_h
    port map (
            O => \N__37940\,
            I => \N__37924\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__37937\,
            I => \N__37921\
        );

    \I__9029\ : Odrv4
    port map (
            O => \N__37934\,
            I => \read_data_RNI4PFJ1_0\
        );

    \I__9028\ : Odrv12
    port map (
            O => \N__37929\,
            I => \read_data_RNI4PFJ1_0\
        );

    \I__9027\ : Odrv4
    port map (
            O => \N__37924\,
            I => \read_data_RNI4PFJ1_0\
        );

    \I__9026\ : Odrv12
    port map (
            O => \N__37921\,
            I => \read_data_RNI4PFJ1_0\
        );

    \I__9025\ : CascadeMux
    port map (
            O => \N__37912\,
            I => \N__37909\
        );

    \I__9024\ : InMux
    port map (
            O => \N__37909\,
            I => \N__37906\
        );

    \I__9023\ : LocalMux
    port map (
            O => \N__37906\,
            I => \N__37903\
        );

    \I__9022\ : Odrv4
    port map (
            O => \N__37903\,
            I => \N_1058\
        );

    \I__9021\ : CascadeMux
    port map (
            O => \N__37900\,
            I => \N_1062_cascade_\
        );

    \I__9020\ : InMux
    port map (
            O => \N__37897\,
            I => \N__37894\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__37894\,
            I => \M_this_map_address_qc_5_0\
        );

    \I__9018\ : InMux
    port map (
            O => \N__37891\,
            I => \N__37888\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__37888\,
            I => \N__37885\
        );

    \I__9016\ : Sp12to4
    port map (
            O => \N__37885\,
            I => \N__37882\
        );

    \I__9015\ : Span12Mux_v
    port map (
            O => \N__37882\,
            I => \N__37879\
        );

    \I__9014\ : Span12Mux_h
    port map (
            O => \N__37879\,
            I => \N__37876\
        );

    \I__9013\ : Odrv12
    port map (
            O => \N__37876\,
            I => \this_spr_ram.mem_out_bus7_2\
        );

    \I__9012\ : InMux
    port map (
            O => \N__37873\,
            I => \N__37870\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__37870\,
            I => \N__37867\
        );

    \I__9010\ : Span4Mux_v
    port map (
            O => \N__37867\,
            I => \N__37864\
        );

    \I__9009\ : Odrv4
    port map (
            O => \N__37864\,
            I => \this_spr_ram.mem_out_bus3_2\
        );

    \I__9008\ : InMux
    port map (
            O => \N__37861\,
            I => \N__37858\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__37858\,
            I => \N__37855\
        );

    \I__9006\ : Span4Mux_h
    port map (
            O => \N__37855\,
            I => \N__37852\
        );

    \I__9005\ : Odrv4
    port map (
            O => \N__37852\,
            I => \this_spr_ram.mem_mem_3_1_RNISI5GZ0\
        );

    \I__9004\ : CascadeMux
    port map (
            O => \N__37849\,
            I => \N__37846\
        );

    \I__9003\ : InMux
    port map (
            O => \N__37846\,
            I => \N__37843\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__37843\,
            I => \N__37840\
        );

    \I__9001\ : Span12Mux_h
    port map (
            O => \N__37840\,
            I => \N__37837\
        );

    \I__9000\ : Span12Mux_v
    port map (
            O => \N__37837\,
            I => \N__37834\
        );

    \I__8999\ : Odrv12
    port map (
            O => \N__37834\,
            I => \this_spr_ram.mem_out_bus7_3\
        );

    \I__8998\ : InMux
    port map (
            O => \N__37831\,
            I => \N__37828\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__37828\,
            I => \N__37825\
        );

    \I__8996\ : Span4Mux_h
    port map (
            O => \N__37825\,
            I => \N__37822\
        );

    \I__8995\ : Odrv4
    port map (
            O => \N__37822\,
            I => \this_spr_ram.mem_out_bus3_3\
        );

    \I__8994\ : InMux
    port map (
            O => \N__37819\,
            I => \N__37816\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__37816\,
            I => \this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0\
        );

    \I__8992\ : InMux
    port map (
            O => \N__37813\,
            I => \N__37810\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__37810\,
            I => \N__37807\
        );

    \I__8990\ : Span4Mux_v
    port map (
            O => \N__37807\,
            I => \N__37804\
        );

    \I__8989\ : Sp12to4
    port map (
            O => \N__37804\,
            I => \N__37801\
        );

    \I__8988\ : Span12Mux_h
    port map (
            O => \N__37801\,
            I => \N__37797\
        );

    \I__8987\ : InMux
    port map (
            O => \N__37800\,
            I => \N__37794\
        );

    \I__8986\ : Odrv12
    port map (
            O => \N__37797\,
            I => \M_this_ctrl_flags_qZ0Z_7\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__37794\,
            I => \M_this_ctrl_flags_qZ0Z_7\
        );

    \I__8984\ : InMux
    port map (
            O => \N__37789\,
            I => \N__37786\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__37786\,
            I => \N__37782\
        );

    \I__8982\ : InMux
    port map (
            O => \N__37785\,
            I => \N__37778\
        );

    \I__8981\ : Span4Mux_v
    port map (
            O => \N__37782\,
            I => \N__37775\
        );

    \I__8980\ : InMux
    port map (
            O => \N__37781\,
            I => \N__37772\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__37778\,
            I => \N__37769\
        );

    \I__8978\ : Odrv4
    port map (
            O => \N__37775\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__37772\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__8976\ : Odrv4
    port map (
            O => \N__37769\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__8975\ : IoInMux
    port map (
            O => \N__37762\,
            I => \N__37759\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__37759\,
            I => \N__37756\
        );

    \I__8973\ : Span4Mux_s2_h
    port map (
            O => \N__37756\,
            I => \N__37752\
        );

    \I__8972\ : InMux
    port map (
            O => \N__37755\,
            I => \N__37749\
        );

    \I__8971\ : Sp12to4
    port map (
            O => \N__37752\,
            I => \N__37744\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__37749\,
            I => \N__37741\
        );

    \I__8969\ : InMux
    port map (
            O => \N__37748\,
            I => \N__37737\
        );

    \I__8968\ : InMux
    port map (
            O => \N__37747\,
            I => \N__37731\
        );

    \I__8967\ : Span12Mux_s10_v
    port map (
            O => \N__37744\,
            I => \N__37727\
        );

    \I__8966\ : Span4Mux_v
    port map (
            O => \N__37741\,
            I => \N__37724\
        );

    \I__8965\ : InMux
    port map (
            O => \N__37740\,
            I => \N__37721\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__37737\,
            I => \N__37718\
        );

    \I__8963\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37715\
        );

    \I__8962\ : InMux
    port map (
            O => \N__37735\,
            I => \N__37712\
        );

    \I__8961\ : InMux
    port map (
            O => \N__37734\,
            I => \N__37709\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__37731\,
            I => \N__37706\
        );

    \I__8959\ : InMux
    port map (
            O => \N__37730\,
            I => \N__37703\
        );

    \I__8958\ : Span12Mux_h
    port map (
            O => \N__37727\,
            I => \N__37700\
        );

    \I__8957\ : Sp12to4
    port map (
            O => \N__37724\,
            I => \N__37697\
        );

    \I__8956\ : LocalMux
    port map (
            O => \N__37721\,
            I => \N__37693\
        );

    \I__8955\ : Span4Mux_v
    port map (
            O => \N__37718\,
            I => \N__37688\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__37715\,
            I => \N__37688\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__37712\,
            I => \N__37685\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__37709\,
            I => \N__37682\
        );

    \I__8951\ : Span4Mux_v
    port map (
            O => \N__37706\,
            I => \N__37677\
        );

    \I__8950\ : LocalMux
    port map (
            O => \N__37703\,
            I => \N__37677\
        );

    \I__8949\ : Span12Mux_v
    port map (
            O => \N__37700\,
            I => \N__37674\
        );

    \I__8948\ : Span12Mux_s6_h
    port map (
            O => \N__37697\,
            I => \N__37671\
        );

    \I__8947\ : InMux
    port map (
            O => \N__37696\,
            I => \N__37668\
        );

    \I__8946\ : Span4Mux_v
    port map (
            O => \N__37693\,
            I => \N__37665\
        );

    \I__8945\ : Span4Mux_h
    port map (
            O => \N__37688\,
            I => \N__37662\
        );

    \I__8944\ : Span12Mux_h
    port map (
            O => \N__37685\,
            I => \N__37657\
        );

    \I__8943\ : Span12Mux_h
    port map (
            O => \N__37682\,
            I => \N__37657\
        );

    \I__8942\ : Span4Mux_h
    port map (
            O => \N__37677\,
            I => \N__37654\
        );

    \I__8941\ : Odrv12
    port map (
            O => \N__37674\,
            I => \N_38_i_0\
        );

    \I__8940\ : Odrv12
    port map (
            O => \N__37671\,
            I => \N_38_i_0\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__37668\,
            I => \N_38_i_0\
        );

    \I__8938\ : Odrv4
    port map (
            O => \N__37665\,
            I => \N_38_i_0\
        );

    \I__8937\ : Odrv4
    port map (
            O => \N__37662\,
            I => \N_38_i_0\
        );

    \I__8936\ : Odrv12
    port map (
            O => \N__37657\,
            I => \N_38_i_0\
        );

    \I__8935\ : Odrv4
    port map (
            O => \N__37654\,
            I => \N_38_i_0\
        );

    \I__8934\ : IoInMux
    port map (
            O => \N__37639\,
            I => \N__37636\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__37636\,
            I => \N__37632\
        );

    \I__8932\ : IoInMux
    port map (
            O => \N__37635\,
            I => \N__37629\
        );

    \I__8931\ : IoSpan4Mux
    port map (
            O => \N__37632\,
            I => \N__37624\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__37629\,
            I => \N__37624\
        );

    \I__8929\ : IoSpan4Mux
    port map (
            O => \N__37624\,
            I => \N__37619\
        );

    \I__8928\ : IoInMux
    port map (
            O => \N__37623\,
            I => \N__37616\
        );

    \I__8927\ : IoInMux
    port map (
            O => \N__37622\,
            I => \N__37613\
        );

    \I__8926\ : IoSpan4Mux
    port map (
            O => \N__37619\,
            I => \N__37601\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__37616\,
            I => \N__37601\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__37613\,
            I => \N__37598\
        );

    \I__8923\ : IoInMux
    port map (
            O => \N__37612\,
            I => \N__37595\
        );

    \I__8922\ : IoInMux
    port map (
            O => \N__37611\,
            I => \N__37592\
        );

    \I__8921\ : IoInMux
    port map (
            O => \N__37610\,
            I => \N__37589\
        );

    \I__8920\ : IoInMux
    port map (
            O => \N__37609\,
            I => \N__37586\
        );

    \I__8919\ : IoInMux
    port map (
            O => \N__37608\,
            I => \N__37581\
        );

    \I__8918\ : IoInMux
    port map (
            O => \N__37607\,
            I => \N__37578\
        );

    \I__8917\ : IoInMux
    port map (
            O => \N__37606\,
            I => \N__37573\
        );

    \I__8916\ : IoSpan4Mux
    port map (
            O => \N__37601\,
            I => \N__37570\
        );

    \I__8915\ : IoSpan4Mux
    port map (
            O => \N__37598\,
            I => \N__37563\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__37595\,
            I => \N__37563\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__37592\,
            I => \N__37563\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__37589\,
            I => \N__37558\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__37586\,
            I => \N__37555\
        );

    \I__8910\ : IoInMux
    port map (
            O => \N__37585\,
            I => \N__37552\
        );

    \I__8909\ : IoInMux
    port map (
            O => \N__37584\,
            I => \N__37549\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__37581\,
            I => \N__37544\
        );

    \I__8907\ : LocalMux
    port map (
            O => \N__37578\,
            I => \N__37544\
        );

    \I__8906\ : IoInMux
    port map (
            O => \N__37577\,
            I => \N__37541\
        );

    \I__8905\ : IoInMux
    port map (
            O => \N__37576\,
            I => \N__37538\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__37573\,
            I => \N__37535\
        );

    \I__8903\ : IoSpan4Mux
    port map (
            O => \N__37570\,
            I => \N__37530\
        );

    \I__8902\ : IoSpan4Mux
    port map (
            O => \N__37563\,
            I => \N__37530\
        );

    \I__8901\ : IoInMux
    port map (
            O => \N__37562\,
            I => \N__37527\
        );

    \I__8900\ : IoInMux
    port map (
            O => \N__37561\,
            I => \N__37524\
        );

    \I__8899\ : IoSpan4Mux
    port map (
            O => \N__37558\,
            I => \N__37521\
        );

    \I__8898\ : IoSpan4Mux
    port map (
            O => \N__37555\,
            I => \N__37514\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__37552\,
            I => \N__37514\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__37549\,
            I => \N__37514\
        );

    \I__8895\ : IoSpan4Mux
    port map (
            O => \N__37544\,
            I => \N__37507\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__37541\,
            I => \N__37507\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__37538\,
            I => \N__37507\
        );

    \I__8892\ : Span4Mux_s1_h
    port map (
            O => \N__37535\,
            I => \N__37504\
        );

    \I__8891\ : Span4Mux_s1_h
    port map (
            O => \N__37530\,
            I => \N__37501\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__37527\,
            I => \N__37496\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__37524\,
            I => \N__37496\
        );

    \I__8888\ : Span4Mux_s3_h
    port map (
            O => \N__37521\,
            I => \N__37493\
        );

    \I__8887\ : IoSpan4Mux
    port map (
            O => \N__37514\,
            I => \N__37488\
        );

    \I__8886\ : IoSpan4Mux
    port map (
            O => \N__37507\,
            I => \N__37488\
        );

    \I__8885\ : Span4Mux_v
    port map (
            O => \N__37504\,
            I => \N__37481\
        );

    \I__8884\ : Span4Mux_v
    port map (
            O => \N__37501\,
            I => \N__37481\
        );

    \I__8883\ : Span4Mux_s1_h
    port map (
            O => \N__37496\,
            I => \N__37481\
        );

    \I__8882\ : Sp12to4
    port map (
            O => \N__37493\,
            I => \N__37478\
        );

    \I__8881\ : Span4Mux_s3_v
    port map (
            O => \N__37488\,
            I => \N__37475\
        );

    \I__8880\ : Span4Mux_h
    port map (
            O => \N__37481\,
            I => \N__37472\
        );

    \I__8879\ : Span12Mux_s11_h
    port map (
            O => \N__37478\,
            I => \N__37469\
        );

    \I__8878\ : Span4Mux_v
    port map (
            O => \N__37475\,
            I => \N__37464\
        );

    \I__8877\ : Span4Mux_h
    port map (
            O => \N__37472\,
            I => \N__37464\
        );

    \I__8876\ : Odrv12
    port map (
            O => \N__37469\,
            I => \N_38_i_0_i\
        );

    \I__8875\ : Odrv4
    port map (
            O => \N__37464\,
            I => \N_38_i_0_i\
        );

    \I__8874\ : InMux
    port map (
            O => \N__37459\,
            I => \N__37456\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__37456\,
            I => \N__37452\
        );

    \I__8872\ : InMux
    port map (
            O => \N__37455\,
            I => \N__37449\
        );

    \I__8871\ : Span4Mux_h
    port map (
            O => \N__37452\,
            I => \N__37446\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__37449\,
            I => \this_ppu.N_856_0\
        );

    \I__8869\ : Odrv4
    port map (
            O => \N__37446\,
            I => \this_ppu.N_856_0\
        );

    \I__8868\ : CascadeMux
    port map (
            O => \N__37441\,
            I => \this_ppu_un1_M_this_state_q_7_i_0_0_0_cascade_\
        );

    \I__8867\ : InMux
    port map (
            O => \N__37438\,
            I => \N__37434\
        );

    \I__8866\ : InMux
    port map (
            O => \N__37437\,
            I => \N__37431\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__37434\,
            I => \N__37428\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__37431\,
            I => \N__37423\
        );

    \I__8863\ : Span4Mux_h
    port map (
            O => \N__37428\,
            I => \N__37420\
        );

    \I__8862\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37417\
        );

    \I__8861\ : InMux
    port map (
            O => \N__37426\,
            I => \N__37414\
        );

    \I__8860\ : Odrv12
    port map (
            O => \N__37423\,
            I => \N_816_0\
        );

    \I__8859\ : Odrv4
    port map (
            O => \N__37420\,
            I => \N_816_0\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__37417\,
            I => \N_816_0\
        );

    \I__8857\ : LocalMux
    port map (
            O => \N__37414\,
            I => \N_816_0\
        );

    \I__8856\ : InMux
    port map (
            O => \N__37405\,
            I => \N__37402\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__37402\,
            I => \N_1416\
        );

    \I__8854\ : InMux
    port map (
            O => \N__37399\,
            I => \N__37396\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__37396\,
            I => \N__37391\
        );

    \I__8852\ : InMux
    port map (
            O => \N__37395\,
            I => \N__37388\
        );

    \I__8851\ : InMux
    port map (
            O => \N__37394\,
            I => \N__37383\
        );

    \I__8850\ : Span4Mux_v
    port map (
            O => \N__37391\,
            I => \N__37378\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__37388\,
            I => \N__37378\
        );

    \I__8848\ : InMux
    port map (
            O => \N__37387\,
            I => \N__37375\
        );

    \I__8847\ : InMux
    port map (
            O => \N__37386\,
            I => \N__37372\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__37383\,
            I => \N__37369\
        );

    \I__8845\ : Odrv4
    port map (
            O => \N__37378\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__37375\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__37372\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__8842\ : Odrv4
    port map (
            O => \N__37369\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__8841\ : IoInMux
    port map (
            O => \N__37360\,
            I => \N__37357\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__37357\,
            I => \N__37354\
        );

    \I__8839\ : Span12Mux_s9_h
    port map (
            O => \N__37354\,
            I => \N__37351\
        );

    \I__8838\ : Span12Mux_v
    port map (
            O => \N__37351\,
            I => \N__37348\
        );

    \I__8837\ : Odrv12
    port map (
            O => \N__37348\,
            I => led_c_6
        );

    \I__8836\ : CascadeMux
    port map (
            O => \N__37345\,
            I => \N__37340\
        );

    \I__8835\ : InMux
    port map (
            O => \N__37344\,
            I => \N__37337\
        );

    \I__8834\ : InMux
    port map (
            O => \N__37343\,
            I => \N__37334\
        );

    \I__8833\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37331\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__37337\,
            I => \N__37322\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__37334\,
            I => \N__37322\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__37331\,
            I => \N__37322\
        );

    \I__8829\ : InMux
    port map (
            O => \N__37330\,
            I => \N__37319\
        );

    \I__8828\ : InMux
    port map (
            O => \N__37329\,
            I => \N__37315\
        );

    \I__8827\ : Span4Mux_h
    port map (
            O => \N__37322\,
            I => \N__37312\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__37319\,
            I => \N__37309\
        );

    \I__8825\ : InMux
    port map (
            O => \N__37318\,
            I => \N__37306\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__37315\,
            I => \N__37303\
        );

    \I__8823\ : Span4Mux_h
    port map (
            O => \N__37312\,
            I => \N__37298\
        );

    \I__8822\ : Span4Mux_v
    port map (
            O => \N__37309\,
            I => \N__37298\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__37306\,
            I => \this_ppu.M_screen_y_qZ0Z_4\
        );

    \I__8820\ : Odrv4
    port map (
            O => \N__37303\,
            I => \this_ppu.M_screen_y_qZ0Z_4\
        );

    \I__8819\ : Odrv4
    port map (
            O => \N__37298\,
            I => \this_ppu.M_screen_y_qZ0Z_4\
        );

    \I__8818\ : InMux
    port map (
            O => \N__37291\,
            I => \N__37286\
        );

    \I__8817\ : InMux
    port map (
            O => \N__37290\,
            I => \N__37283\
        );

    \I__8816\ : InMux
    port map (
            O => \N__37289\,
            I => \N__37280\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__37286\,
            I => \N__37275\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__37283\,
            I => \N__37275\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__37280\,
            I => \N__37272\
        );

    \I__8812\ : Span12Mux_h
    port map (
            O => \N__37275\,
            I => \N__37269\
        );

    \I__8811\ : Odrv4
    port map (
            O => \N__37272\,
            I => \this_ppu.un3_M_screen_y_d_0_c4\
        );

    \I__8810\ : Odrv12
    port map (
            O => \N__37269\,
            I => \this_ppu.un3_M_screen_y_d_0_c4\
        );

    \I__8809\ : InMux
    port map (
            O => \N__37264\,
            I => \N__37261\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__37261\,
            I => \N__37256\
        );

    \I__8807\ : InMux
    port map (
            O => \N__37260\,
            I => \N__37245\
        );

    \I__8806\ : InMux
    port map (
            O => \N__37259\,
            I => \N__37245\
        );

    \I__8805\ : Span4Mux_h
    port map (
            O => \N__37256\,
            I => \N__37242\
        );

    \I__8804\ : CascadeMux
    port map (
            O => \N__37255\,
            I => \N__37239\
        );

    \I__8803\ : InMux
    port map (
            O => \N__37254\,
            I => \N__37222\
        );

    \I__8802\ : InMux
    port map (
            O => \N__37253\,
            I => \N__37222\
        );

    \I__8801\ : InMux
    port map (
            O => \N__37252\,
            I => \N__37222\
        );

    \I__8800\ : InMux
    port map (
            O => \N__37251\,
            I => \N__37222\
        );

    \I__8799\ : InMux
    port map (
            O => \N__37250\,
            I => \N__37222\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__37245\,
            I => \N__37219\
        );

    \I__8797\ : Span4Mux_h
    port map (
            O => \N__37242\,
            I => \N__37216\
        );

    \I__8796\ : InMux
    port map (
            O => \N__37239\,
            I => \N__37213\
        );

    \I__8795\ : InMux
    port map (
            O => \N__37238\,
            I => \N__37210\
        );

    \I__8794\ : InMux
    port map (
            O => \N__37237\,
            I => \N__37207\
        );

    \I__8793\ : InMux
    port map (
            O => \N__37236\,
            I => \N__37200\
        );

    \I__8792\ : InMux
    port map (
            O => \N__37235\,
            I => \N__37200\
        );

    \I__8791\ : InMux
    port map (
            O => \N__37234\,
            I => \N__37200\
        );

    \I__8790\ : InMux
    port map (
            O => \N__37233\,
            I => \N__37197\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__37222\,
            I => \N__37194\
        );

    \I__8788\ : Odrv4
    port map (
            O => \N__37219\,
            I => \N_861_0\
        );

    \I__8787\ : Odrv4
    port map (
            O => \N__37216\,
            I => \N_861_0\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__37213\,
            I => \N_861_0\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__37210\,
            I => \N_861_0\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__37207\,
            I => \N_861_0\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__37200\,
            I => \N_861_0\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__37197\,
            I => \N_861_0\
        );

    \I__8781\ : Odrv4
    port map (
            O => \N__37194\,
            I => \N_861_0\
        );

    \I__8780\ : CEMux
    port map (
            O => \N__37177\,
            I => \N__37173\
        );

    \I__8779\ : CEMux
    port map (
            O => \N__37176\,
            I => \N__37170\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__37173\,
            I => \N__37166\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__37170\,
            I => \N__37162\
        );

    \I__8776\ : CEMux
    port map (
            O => \N__37169\,
            I => \N__37159\
        );

    \I__8775\ : Span4Mux_v
    port map (
            O => \N__37166\,
            I => \N__37156\
        );

    \I__8774\ : CEMux
    port map (
            O => \N__37165\,
            I => \N__37153\
        );

    \I__8773\ : Span4Mux_h
    port map (
            O => \N__37162\,
            I => \N__37150\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__37159\,
            I => \N__37147\
        );

    \I__8771\ : Sp12to4
    port map (
            O => \N__37156\,
            I => \N__37142\
        );

    \I__8770\ : LocalMux
    port map (
            O => \N__37153\,
            I => \N__37142\
        );

    \I__8769\ : Odrv4
    port map (
            O => \N__37150\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_0\
        );

    \I__8768\ : Odrv4
    port map (
            O => \N__37147\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_0\
        );

    \I__8767\ : Odrv12
    port map (
            O => \N__37142\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_0\
        );

    \I__8766\ : InMux
    port map (
            O => \N__37135\,
            I => \N__37130\
        );

    \I__8765\ : CascadeMux
    port map (
            O => \N__37134\,
            I => \N__37127\
        );

    \I__8764\ : CascadeMux
    port map (
            O => \N__37133\,
            I => \N__37124\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__37130\,
            I => \N__37119\
        );

    \I__8762\ : InMux
    port map (
            O => \N__37127\,
            I => \N__37116\
        );

    \I__8761\ : InMux
    port map (
            O => \N__37124\,
            I => \N__37111\
        );

    \I__8760\ : InMux
    port map (
            O => \N__37123\,
            I => \N__37111\
        );

    \I__8759\ : InMux
    port map (
            O => \N__37122\,
            I => \N__37108\
        );

    \I__8758\ : Span12Mux_h
    port map (
            O => \N__37119\,
            I => \N__37105\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__37116\,
            I => \N__37100\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__37111\,
            I => \N__37100\
        );

    \I__8755\ : LocalMux
    port map (
            O => \N__37108\,
            I => \this_ppu.M_screen_y_qZ0Z_5\
        );

    \I__8754\ : Odrv12
    port map (
            O => \N__37105\,
            I => \this_ppu.M_screen_y_qZ0Z_5\
        );

    \I__8753\ : Odrv4
    port map (
            O => \N__37100\,
            I => \this_ppu.M_screen_y_qZ0Z_5\
        );

    \I__8752\ : CascadeMux
    port map (
            O => \N__37093\,
            I => \N__37090\
        );

    \I__8751\ : InMux
    port map (
            O => \N__37090\,
            I => \N__37087\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__37087\,
            I => \N__37083\
        );

    \I__8749\ : CascadeMux
    port map (
            O => \N__37086\,
            I => \N__37080\
        );

    \I__8748\ : Span4Mux_v
    port map (
            O => \N__37083\,
            I => \N__37077\
        );

    \I__8747\ : InMux
    port map (
            O => \N__37080\,
            I => \N__37074\
        );

    \I__8746\ : Span4Mux_h
    port map (
            O => \N__37077\,
            I => \N__37071\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__37074\,
            I => \N__37068\
        );

    \I__8744\ : Span4Mux_h
    port map (
            O => \N__37071\,
            I => \N__37063\
        );

    \I__8743\ : Span4Mux_h
    port map (
            O => \N__37068\,
            I => \N__37063\
        );

    \I__8742\ : Odrv4
    port map (
            O => \N__37063\,
            I => \M_this_scroll_qZ0Z_5\
        );

    \I__8741\ : InMux
    port map (
            O => \N__37060\,
            I => \N__37057\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__37057\,
            I => \N__37054\
        );

    \I__8739\ : Span4Mux_h
    port map (
            O => \N__37054\,
            I => \N__37051\
        );

    \I__8738\ : Span4Mux_h
    port map (
            O => \N__37051\,
            I => \N__37048\
        );

    \I__8737\ : Span4Mux_h
    port map (
            O => \N__37048\,
            I => \N__37045\
        );

    \I__8736\ : Odrv4
    port map (
            O => \N__37045\,
            I => \this_ppu.M_screen_y_q_esr_RNIJB7F7Z0Z_5\
        );

    \I__8735\ : CascadeMux
    port map (
            O => \N__37042\,
            I => \N__37039\
        );

    \I__8734\ : InMux
    port map (
            O => \N__37039\,
            I => \N__37034\
        );

    \I__8733\ : InMux
    port map (
            O => \N__37038\,
            I => \N__37031\
        );

    \I__8732\ : InMux
    port map (
            O => \N__37037\,
            I => \N__37028\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__37034\,
            I => \N__37020\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__37031\,
            I => \N__37020\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__37028\,
            I => \N__37020\
        );

    \I__8728\ : InMux
    port map (
            O => \N__37027\,
            I => \N__37017\
        );

    \I__8727\ : Span4Mux_v
    port map (
            O => \N__37020\,
            I => \N__37014\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__37017\,
            I => \this_spr_ram.mem_radregZ0Z_12\
        );

    \I__8725\ : Odrv4
    port map (
            O => \N__37014\,
            I => \this_spr_ram.mem_radregZ0Z_12\
        );

    \I__8724\ : InMux
    port map (
            O => \N__37009\,
            I => \N__37006\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__37006\,
            I => \this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0\
        );

    \I__8722\ : CascadeMux
    port map (
            O => \N__37003\,
            I => \N__36996\
        );

    \I__8721\ : InMux
    port map (
            O => \N__37002\,
            I => \N__36992\
        );

    \I__8720\ : InMux
    port map (
            O => \N__37001\,
            I => \N__36987\
        );

    \I__8719\ : InMux
    port map (
            O => \N__37000\,
            I => \N__36987\
        );

    \I__8718\ : InMux
    port map (
            O => \N__36999\,
            I => \N__36980\
        );

    \I__8717\ : InMux
    port map (
            O => \N__36996\,
            I => \N__36980\
        );

    \I__8716\ : InMux
    port map (
            O => \N__36995\,
            I => \N__36980\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__36992\,
            I => \N__36975\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__36987\,
            I => \N__36972\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__36980\,
            I => \N__36969\
        );

    \I__8712\ : InMux
    port map (
            O => \N__36979\,
            I => \N__36964\
        );

    \I__8711\ : InMux
    port map (
            O => \N__36978\,
            I => \N__36964\
        );

    \I__8710\ : Span4Mux_h
    port map (
            O => \N__36975\,
            I => \N__36961\
        );

    \I__8709\ : Odrv4
    port map (
            O => \N__36972\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__8708\ : Odrv4
    port map (
            O => \N__36969\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__36964\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__8706\ : Odrv4
    port map (
            O => \N__36961\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__8705\ : CascadeMux
    port map (
            O => \N__36952\,
            I => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\
        );

    \I__8704\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36946\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__36946\,
            I => \N__36942\
        );

    \I__8702\ : InMux
    port map (
            O => \N__36945\,
            I => \N__36939\
        );

    \I__8701\ : Odrv4
    port map (
            O => \N__36942\,
            I => \M_this_spr_ram_read_data_3\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__36939\,
            I => \M_this_spr_ram_read_data_3\
        );

    \I__8699\ : InMux
    port map (
            O => \N__36934\,
            I => \N__36931\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__36931\,
            I => \N__36928\
        );

    \I__8697\ : Span4Mux_h
    port map (
            O => \N__36928\,
            I => \N__36925\
        );

    \I__8696\ : Span4Mux_v
    port map (
            O => \N__36925\,
            I => \N__36922\
        );

    \I__8695\ : Odrv4
    port map (
            O => \N__36922\,
            I => \this_spr_ram.mem_out_bus5_3\
        );

    \I__8694\ : InMux
    port map (
            O => \N__36919\,
            I => \N__36916\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__36916\,
            I => \N__36913\
        );

    \I__8692\ : Span4Mux_h
    port map (
            O => \N__36913\,
            I => \N__36910\
        );

    \I__8691\ : Span4Mux_v
    port map (
            O => \N__36910\,
            I => \N__36907\
        );

    \I__8690\ : Span4Mux_v
    port map (
            O => \N__36907\,
            I => \N__36904\
        );

    \I__8689\ : Odrv4
    port map (
            O => \N__36904\,
            I => \this_spr_ram.mem_out_bus1_3\
        );

    \I__8688\ : InMux
    port map (
            O => \N__36901\,
            I => \N__36898\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__36898\,
            I => \this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0\
        );

    \I__8686\ : InMux
    port map (
            O => \N__36895\,
            I => \N__36892\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__36892\,
            I => \N__36889\
        );

    \I__8684\ : Span12Mux_h
    port map (
            O => \N__36889\,
            I => \N__36886\
        );

    \I__8683\ : Span12Mux_h
    port map (
            O => \N__36886\,
            I => \N__36883\
        );

    \I__8682\ : Odrv12
    port map (
            O => \N__36883\,
            I => \this_spr_ram.mem_out_bus6_3\
        );

    \I__8681\ : InMux
    port map (
            O => \N__36880\,
            I => \N__36877\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__36877\,
            I => \N__36874\
        );

    \I__8679\ : Span4Mux_h
    port map (
            O => \N__36874\,
            I => \N__36871\
        );

    \I__8678\ : Span4Mux_v
    port map (
            O => \N__36871\,
            I => \N__36868\
        );

    \I__8677\ : Odrv4
    port map (
            O => \N__36868\,
            I => \this_spr_ram.mem_out_bus2_3\
        );

    \I__8676\ : InMux
    port map (
            O => \N__36865\,
            I => \N__36862\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__36862\,
            I => \this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0\
        );

    \I__8674\ : InMux
    port map (
            O => \N__36859\,
            I => \N__36856\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__36856\,
            I => \N__36853\
        );

    \I__8672\ : Span4Mux_v
    port map (
            O => \N__36853\,
            I => \N__36850\
        );

    \I__8671\ : Span4Mux_h
    port map (
            O => \N__36850\,
            I => \N__36847\
        );

    \I__8670\ : Sp12to4
    port map (
            O => \N__36847\,
            I => \N__36844\
        );

    \I__8669\ : Span12Mux_h
    port map (
            O => \N__36844\,
            I => \N__36841\
        );

    \I__8668\ : Odrv12
    port map (
            O => \N__36841\,
            I => \this_spr_ram.mem_out_bus7_0\
        );

    \I__8667\ : InMux
    port map (
            O => \N__36838\,
            I => \N__36835\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__36835\,
            I => \N__36832\
        );

    \I__8665\ : Span4Mux_h
    port map (
            O => \N__36832\,
            I => \N__36829\
        );

    \I__8664\ : Odrv4
    port map (
            O => \N__36829\,
            I => \this_spr_ram.mem_out_bus3_0\
        );

    \I__8663\ : InMux
    port map (
            O => \N__36826\,
            I => \N__36823\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__36823\,
            I => \this_spr_ram.mem_mem_3_0_RNIQI5GZ0\
        );

    \I__8661\ : InMux
    port map (
            O => \N__36820\,
            I => \N__36817\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__36817\,
            I => \N__36814\
        );

    \I__8659\ : Sp12to4
    port map (
            O => \N__36814\,
            I => \N__36811\
        );

    \I__8658\ : Span12Mux_v
    port map (
            O => \N__36811\,
            I => \N__36808\
        );

    \I__8657\ : Span12Mux_h
    port map (
            O => \N__36808\,
            I => \N__36805\
        );

    \I__8656\ : Odrv12
    port map (
            O => \N__36805\,
            I => \this_spr_ram.mem_out_bus7_1\
        );

    \I__8655\ : InMux
    port map (
            O => \N__36802\,
            I => \N__36799\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__36799\,
            I => \N__36796\
        );

    \I__8653\ : Span4Mux_v
    port map (
            O => \N__36796\,
            I => \N__36793\
        );

    \I__8652\ : Odrv4
    port map (
            O => \N__36793\,
            I => \this_spr_ram.mem_out_bus3_1\
        );

    \I__8651\ : InMux
    port map (
            O => \N__36790\,
            I => \N__36787\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__36787\,
            I => \this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0\
        );

    \I__8649\ : InMux
    port map (
            O => \N__36784\,
            I => \N__36781\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__36781\,
            I => \N__36778\
        );

    \I__8647\ : Span4Mux_h
    port map (
            O => \N__36778\,
            I => \N__36775\
        );

    \I__8646\ : Sp12to4
    port map (
            O => \N__36775\,
            I => \N__36772\
        );

    \I__8645\ : Odrv12
    port map (
            O => \N__36772\,
            I => \this_spr_ram.mem_out_bus5_2\
        );

    \I__8644\ : InMux
    port map (
            O => \N__36769\,
            I => \N__36766\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__36766\,
            I => \N__36763\
        );

    \I__8642\ : Span4Mux_h
    port map (
            O => \N__36763\,
            I => \N__36760\
        );

    \I__8641\ : Span4Mux_v
    port map (
            O => \N__36760\,
            I => \N__36757\
        );

    \I__8640\ : Odrv4
    port map (
            O => \N__36757\,
            I => \this_spr_ram.mem_out_bus1_2\
        );

    \I__8639\ : InMux
    port map (
            O => \N__36754\,
            I => \N__36751\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__36751\,
            I => \this_spr_ram.mem_mem_1_1_RNIOA1GZ0\
        );

    \I__8637\ : InMux
    port map (
            O => \N__36748\,
            I => \N__36745\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__36745\,
            I => \N__36742\
        );

    \I__8635\ : Span4Mux_v
    port map (
            O => \N__36742\,
            I => \N__36739\
        );

    \I__8634\ : Span4Mux_v
    port map (
            O => \N__36739\,
            I => \N__36736\
        );

    \I__8633\ : Span4Mux_v
    port map (
            O => \N__36736\,
            I => \N__36733\
        );

    \I__8632\ : Odrv4
    port map (
            O => \N__36733\,
            I => \this_spr_ram.mem_out_bus6_0\
        );

    \I__8631\ : InMux
    port map (
            O => \N__36730\,
            I => \N__36727\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__36727\,
            I => \N__36724\
        );

    \I__8629\ : Span4Mux_v
    port map (
            O => \N__36724\,
            I => \N__36721\
        );

    \I__8628\ : Span4Mux_v
    port map (
            O => \N__36721\,
            I => \N__36718\
        );

    \I__8627\ : Odrv4
    port map (
            O => \N__36718\,
            I => \this_spr_ram.mem_out_bus2_0\
        );

    \I__8626\ : CascadeMux
    port map (
            O => \N__36715\,
            I => \this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_\
        );

    \I__8625\ : InMux
    port map (
            O => \N__36712\,
            I => \N__36709\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__36709\,
            I => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_0\
        );

    \I__8623\ : CEMux
    port map (
            O => \N__36706\,
            I => \N__36703\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__36703\,
            I => \N__36699\
        );

    \I__8621\ : CEMux
    port map (
            O => \N__36702\,
            I => \N__36696\
        );

    \I__8620\ : Span4Mux_s2_v
    port map (
            O => \N__36699\,
            I => \N__36691\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__36696\,
            I => \N__36691\
        );

    \I__8618\ : Span4Mux_h
    port map (
            O => \N__36691\,
            I => \N__36688\
        );

    \I__8617\ : Span4Mux_h
    port map (
            O => \N__36688\,
            I => \N__36685\
        );

    \I__8616\ : Sp12to4
    port map (
            O => \N__36685\,
            I => \N__36682\
        );

    \I__8615\ : Span12Mux_v
    port map (
            O => \N__36682\,
            I => \N__36679\
        );

    \I__8614\ : Odrv12
    port map (
            O => \N__36679\,
            I => \this_spr_ram.mem_WE_0\
        );

    \I__8613\ : InMux
    port map (
            O => \N__36676\,
            I => \N__36673\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__36673\,
            I => \N__36670\
        );

    \I__8611\ : Sp12to4
    port map (
            O => \N__36670\,
            I => \N__36667\
        );

    \I__8610\ : Span12Mux_h
    port map (
            O => \N__36667\,
            I => \N__36664\
        );

    \I__8609\ : Odrv12
    port map (
            O => \N__36664\,
            I => \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_7\
        );

    \I__8608\ : InMux
    port map (
            O => \N__36661\,
            I => \N__36658\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__36658\,
            I => \N__36655\
        );

    \I__8606\ : Span4Mux_v
    port map (
            O => \N__36655\,
            I => \N__36652\
        );

    \I__8605\ : Span4Mux_h
    port map (
            O => \N__36652\,
            I => \N__36649\
        );

    \I__8604\ : Sp12to4
    port map (
            O => \N__36649\,
            I => \N__36646\
        );

    \I__8603\ : Span12Mux_h
    port map (
            O => \N__36646\,
            I => \N__36643\
        );

    \I__8602\ : Odrv12
    port map (
            O => \N__36643\,
            I => \this_spr_ram.mem_out_bus6_2\
        );

    \I__8601\ : InMux
    port map (
            O => \N__36640\,
            I => \N__36637\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__36637\,
            I => \N__36634\
        );

    \I__8599\ : Span4Mux_h
    port map (
            O => \N__36634\,
            I => \N__36631\
        );

    \I__8598\ : Odrv4
    port map (
            O => \N__36631\,
            I => \this_spr_ram.mem_out_bus2_2\
        );

    \I__8597\ : InMux
    port map (
            O => \N__36628\,
            I => \N__36625\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__36625\,
            I => \this_spr_ram.mem_mem_2_1_RNIQE3GZ0\
        );

    \I__8595\ : InMux
    port map (
            O => \N__36622\,
            I => \N__36619\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__36619\,
            I => \N__36616\
        );

    \I__8593\ : Span4Mux_h
    port map (
            O => \N__36616\,
            I => \N__36613\
        );

    \I__8592\ : Odrv4
    port map (
            O => \N__36613\,
            I => \this_spr_ram.mem_out_bus4_3\
        );

    \I__8591\ : InMux
    port map (
            O => \N__36610\,
            I => \N__36607\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__36607\,
            I => \N__36604\
        );

    \I__8589\ : Span12Mux_h
    port map (
            O => \N__36604\,
            I => \N__36601\
        );

    \I__8588\ : Span12Mux_v
    port map (
            O => \N__36601\,
            I => \N__36598\
        );

    \I__8587\ : Odrv12
    port map (
            O => \N__36598\,
            I => \this_spr_ram.mem_out_bus0_3\
        );

    \I__8586\ : InMux
    port map (
            O => \N__36595\,
            I => \N__36591\
        );

    \I__8585\ : InMux
    port map (
            O => \N__36594\,
            I => \N__36588\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__36591\,
            I => \N__36585\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__36588\,
            I => \N__36582\
        );

    \I__8582\ : Span12Mux_h
    port map (
            O => \N__36585\,
            I => \N__36579\
        );

    \I__8581\ : Span4Mux_h
    port map (
            O => \N__36582\,
            I => \N__36576\
        );

    \I__8580\ : Odrv12
    port map (
            O => \N__36579\,
            I => \this_ppu.N_753_0\
        );

    \I__8579\ : Odrv4
    port map (
            O => \N__36576\,
            I => \this_ppu.N_753_0\
        );

    \I__8578\ : CascadeMux
    port map (
            O => \N__36571\,
            I => \N__36568\
        );

    \I__8577\ : InMux
    port map (
            O => \N__36568\,
            I => \N__36564\
        );

    \I__8576\ : CascadeMux
    port map (
            O => \N__36567\,
            I => \N__36561\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__36564\,
            I => \N__36557\
        );

    \I__8574\ : InMux
    port map (
            O => \N__36561\,
            I => \N__36554\
        );

    \I__8573\ : InMux
    port map (
            O => \N__36560\,
            I => \N__36551\
        );

    \I__8572\ : Span4Mux_v
    port map (
            O => \N__36557\,
            I => \N__36548\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__36554\,
            I => \N__36543\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__36551\,
            I => \N__36543\
        );

    \I__8569\ : Span4Mux_h
    port map (
            O => \N__36548\,
            I => \N__36538\
        );

    \I__8568\ : Span4Mux_v
    port map (
            O => \N__36543\,
            I => \N__36538\
        );

    \I__8567\ : Odrv4
    port map (
            O => \N__36538\,
            I => \this_ppu.M_screen_y_qZ0Z_6\
        );

    \I__8566\ : InMux
    port map (
            O => \N__36535\,
            I => \N__36528\
        );

    \I__8565\ : InMux
    port map (
            O => \N__36534\,
            I => \N__36525\
        );

    \I__8564\ : InMux
    port map (
            O => \N__36533\,
            I => \N__36522\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__36532\,
            I => \N__36519\
        );

    \I__8562\ : InMux
    port map (
            O => \N__36531\,
            I => \N__36515\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__36528\,
            I => \N__36506\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__36525\,
            I => \N__36506\
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__36522\,
            I => \N__36506\
        );

    \I__8558\ : InMux
    port map (
            O => \N__36519\,
            I => \N__36503\
        );

    \I__8557\ : InMux
    port map (
            O => \N__36518\,
            I => \N__36500\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__36515\,
            I => \N__36497\
        );

    \I__8555\ : InMux
    port map (
            O => \N__36514\,
            I => \N__36492\
        );

    \I__8554\ : InMux
    port map (
            O => \N__36513\,
            I => \N__36492\
        );

    \I__8553\ : Span4Mux_v
    port map (
            O => \N__36506\,
            I => \N__36485\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__36503\,
            I => \N__36485\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__36500\,
            I => \N__36485\
        );

    \I__8550\ : Span4Mux_h
    port map (
            O => \N__36497\,
            I => \N__36479\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__36492\,
            I => \N__36479\
        );

    \I__8548\ : Span4Mux_h
    port map (
            O => \N__36485\,
            I => \N__36473\
        );

    \I__8547\ : InMux
    port map (
            O => \N__36484\,
            I => \N__36470\
        );

    \I__8546\ : Span4Mux_v
    port map (
            O => \N__36479\,
            I => \N__36467\
        );

    \I__8545\ : InMux
    port map (
            O => \N__36478\,
            I => \N__36462\
        );

    \I__8544\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36462\
        );

    \I__8543\ : InMux
    port map (
            O => \N__36476\,
            I => \N__36459\
        );

    \I__8542\ : Span4Mux_h
    port map (
            O => \N__36473\,
            I => \N__36456\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__36470\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__8540\ : Odrv4
    port map (
            O => \N__36467\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__36462\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__36459\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__8537\ : Odrv4
    port map (
            O => \N__36456\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__8536\ : InMux
    port map (
            O => \N__36445\,
            I => \N__36439\
        );

    \I__8535\ : InMux
    port map (
            O => \N__36444\,
            I => \N__36434\
        );

    \I__8534\ : CascadeMux
    port map (
            O => \N__36443\,
            I => \N__36431\
        );

    \I__8533\ : CascadeMux
    port map (
            O => \N__36442\,
            I => \N__36427\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__36439\,
            I => \N__36424\
        );

    \I__8531\ : InMux
    port map (
            O => \N__36438\,
            I => \N__36421\
        );

    \I__8530\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36418\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__36434\,
            I => \N__36415\
        );

    \I__8528\ : InMux
    port map (
            O => \N__36431\,
            I => \N__36412\
        );

    \I__8527\ : InMux
    port map (
            O => \N__36430\,
            I => \N__36409\
        );

    \I__8526\ : InMux
    port map (
            O => \N__36427\,
            I => \N__36406\
        );

    \I__8525\ : Span4Mux_h
    port map (
            O => \N__36424\,
            I => \N__36403\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__36421\,
            I => \N__36398\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__36418\,
            I => \N__36398\
        );

    \I__8522\ : Span4Mux_v
    port map (
            O => \N__36415\,
            I => \N__36395\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__36412\,
            I => \N__36392\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__36409\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__36406\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8518\ : Odrv4
    port map (
            O => \N__36403\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8517\ : Odrv12
    port map (
            O => \N__36398\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8516\ : Odrv4
    port map (
            O => \N__36395\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8515\ : Odrv4
    port map (
            O => \N__36392\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8514\ : CascadeMux
    port map (
            O => \N__36379\,
            I => \N__36375\
        );

    \I__8513\ : InMux
    port map (
            O => \N__36378\,
            I => \N__36372\
        );

    \I__8512\ : InMux
    port map (
            O => \N__36375\,
            I => \N__36369\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__36372\,
            I => \N__36364\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__36369\,
            I => \N__36364\
        );

    \I__8509\ : Span12Mux_v
    port map (
            O => \N__36364\,
            I => \N__36361\
        );

    \I__8508\ : Odrv12
    port map (
            O => \N__36361\,
            I => \M_this_spr_ram_write_en_0_i_1_0\
        );

    \I__8507\ : CascadeMux
    port map (
            O => \N__36358\,
            I => \N__36355\
        );

    \I__8506\ : InMux
    port map (
            O => \N__36355\,
            I => \N__36351\
        );

    \I__8505\ : InMux
    port map (
            O => \N__36354\,
            I => \N__36347\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__36351\,
            I => \N__36344\
        );

    \I__8503\ : InMux
    port map (
            O => \N__36350\,
            I => \N__36340\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__36347\,
            I => \N__36337\
        );

    \I__8501\ : Span12Mux_h
    port map (
            O => \N__36344\,
            I => \N__36332\
        );

    \I__8500\ : InMux
    port map (
            O => \N__36343\,
            I => \N__36329\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__36340\,
            I => \N__36326\
        );

    \I__8498\ : Span4Mux_v
    port map (
            O => \N__36337\,
            I => \N__36323\
        );

    \I__8497\ : InMux
    port map (
            O => \N__36336\,
            I => \N__36318\
        );

    \I__8496\ : InMux
    port map (
            O => \N__36335\,
            I => \N__36318\
        );

    \I__8495\ : Odrv12
    port map (
            O => \N__36332\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__36329\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__8493\ : Odrv4
    port map (
            O => \N__36326\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__8492\ : Odrv4
    port map (
            O => \N__36323\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__36318\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__8490\ : InMux
    port map (
            O => \N__36307\,
            I => \N__36301\
        );

    \I__8489\ : InMux
    port map (
            O => \N__36306\,
            I => \N__36301\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__36301\,
            I => \N__36295\
        );

    \I__8487\ : InMux
    port map (
            O => \N__36300\,
            I => \N__36288\
        );

    \I__8486\ : InMux
    port map (
            O => \N__36299\,
            I => \N__36288\
        );

    \I__8485\ : InMux
    port map (
            O => \N__36298\,
            I => \N__36288\
        );

    \I__8484\ : Span4Mux_h
    port map (
            O => \N__36295\,
            I => \N__36282\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__36288\,
            I => \N__36282\
        );

    \I__8482\ : CascadeMux
    port map (
            O => \N__36287\,
            I => \N__36279\
        );

    \I__8481\ : Span4Mux_v
    port map (
            O => \N__36282\,
            I => \N__36276\
        );

    \I__8480\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36273\
        );

    \I__8479\ : Span4Mux_v
    port map (
            O => \N__36276\,
            I => \N__36269\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__36273\,
            I => \N__36266\
        );

    \I__8477\ : InMux
    port map (
            O => \N__36272\,
            I => \N__36263\
        );

    \I__8476\ : IoSpan4Mux
    port map (
            O => \N__36269\,
            I => \N__36260\
        );

    \I__8475\ : Span12Mux_h
    port map (
            O => \N__36266\,
            I => \N__36255\
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__36263\,
            I => \N__36255\
        );

    \I__8473\ : Odrv4
    port map (
            O => \N__36260\,
            I => port_address_in_2
        );

    \I__8472\ : Odrv12
    port map (
            O => \N__36255\,
            I => port_address_in_2
        );

    \I__8471\ : CascadeMux
    port map (
            O => \N__36250\,
            I => \N__36247\
        );

    \I__8470\ : InMux
    port map (
            O => \N__36247\,
            I => \N__36244\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__36244\,
            I => \N__36239\
        );

    \I__8468\ : InMux
    port map (
            O => \N__36243\,
            I => \N__36236\
        );

    \I__8467\ : InMux
    port map (
            O => \N__36242\,
            I => \N__36232\
        );

    \I__8466\ : Span4Mux_v
    port map (
            O => \N__36239\,
            I => \N__36227\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__36236\,
            I => \N__36227\
        );

    \I__8464\ : CascadeMux
    port map (
            O => \N__36235\,
            I => \N__36223\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__36232\,
            I => \N__36220\
        );

    \I__8462\ : Span4Mux_h
    port map (
            O => \N__36227\,
            I => \N__36217\
        );

    \I__8461\ : InMux
    port map (
            O => \N__36226\,
            I => \N__36214\
        );

    \I__8460\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36211\
        );

    \I__8459\ : Span4Mux_v
    port map (
            O => \N__36220\,
            I => \N__36207\
        );

    \I__8458\ : Span4Mux_h
    port map (
            O => \N__36217\,
            I => \N__36200\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__36214\,
            I => \N__36200\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__36211\,
            I => \N__36200\
        );

    \I__8455\ : CascadeMux
    port map (
            O => \N__36210\,
            I => \N__36197\
        );

    \I__8454\ : Span4Mux_h
    port map (
            O => \N__36207\,
            I => \N__36192\
        );

    \I__8453\ : Span4Mux_v
    port map (
            O => \N__36200\,
            I => \N__36189\
        );

    \I__8452\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36186\
        );

    \I__8451\ : InMux
    port map (
            O => \N__36196\,
            I => \N__36181\
        );

    \I__8450\ : InMux
    port map (
            O => \N__36195\,
            I => \N__36181\
        );

    \I__8449\ : Sp12to4
    port map (
            O => \N__36192\,
            I => \N__36178\
        );

    \I__8448\ : Span4Mux_h
    port map (
            O => \N__36189\,
            I => \N__36175\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__36186\,
            I => \N__36170\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__36181\,
            I => \N__36170\
        );

    \I__8445\ : Span12Mux_s6_h
    port map (
            O => \N__36178\,
            I => \N__36163\
        );

    \I__8444\ : Sp12to4
    port map (
            O => \N__36175\,
            I => \N__36163\
        );

    \I__8443\ : Span12Mux_h
    port map (
            O => \N__36170\,
            I => \N__36163\
        );

    \I__8442\ : Odrv12
    port map (
            O => \N__36163\,
            I => port_address_in_1
        );

    \I__8441\ : InMux
    port map (
            O => \N__36160\,
            I => \N__36157\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__36157\,
            I => \N__36149\
        );

    \I__8439\ : InMux
    port map (
            O => \N__36156\,
            I => \N__36146\
        );

    \I__8438\ : InMux
    port map (
            O => \N__36155\,
            I => \N__36141\
        );

    \I__8437\ : InMux
    port map (
            O => \N__36154\,
            I => \N__36141\
        );

    \I__8436\ : InMux
    port map (
            O => \N__36153\,
            I => \N__36138\
        );

    \I__8435\ : InMux
    port map (
            O => \N__36152\,
            I => \N__36135\
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__36149\,
            I => \M_this_substate_qZ0\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__36146\,
            I => \M_this_substate_qZ0\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__36141\,
            I => \M_this_substate_qZ0\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__36138\,
            I => \M_this_substate_qZ0\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__36135\,
            I => \M_this_substate_qZ0\
        );

    \I__8429\ : InMux
    port map (
            O => \N__36124\,
            I => \N__36121\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__36121\,
            I => \this_ppu_M_this_substate_d_0_sqmuxa_3_0_a3_0_a3_1\
        );

    \I__8427\ : CascadeMux
    port map (
            O => \N__36118\,
            I => \M_this_map_address_qc_3_0_cascade_\
        );

    \I__8426\ : InMux
    port map (
            O => \N__36115\,
            I => \N__36110\
        );

    \I__8425\ : CascadeMux
    port map (
            O => \N__36114\,
            I => \N__36107\
        );

    \I__8424\ : InMux
    port map (
            O => \N__36113\,
            I => \N__36104\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__36110\,
            I => \N__36101\
        );

    \I__8422\ : InMux
    port map (
            O => \N__36107\,
            I => \N__36096\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__36104\,
            I => \N__36091\
        );

    \I__8420\ : Span4Mux_h
    port map (
            O => \N__36101\,
            I => \N__36091\
        );

    \I__8419\ : InMux
    port map (
            O => \N__36100\,
            I => \N__36088\
        );

    \I__8418\ : InMux
    port map (
            O => \N__36099\,
            I => \N__36085\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__36096\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__8416\ : Odrv4
    port map (
            O => \N__36091\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__36088\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__36085\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__8413\ : InMux
    port map (
            O => \N__36076\,
            I => \N__36073\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__36073\,
            I => \N__36070\
        );

    \I__8411\ : Span4Mux_h
    port map (
            O => \N__36070\,
            I => \N__36067\
        );

    \I__8410\ : Odrv4
    port map (
            O => \N__36067\,
            I => \N_169_0\
        );

    \I__8409\ : IoInMux
    port map (
            O => \N__36064\,
            I => \N__36061\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__36061\,
            I => \N__36058\
        );

    \I__8407\ : IoSpan4Mux
    port map (
            O => \N__36058\,
            I => \N__36055\
        );

    \I__8406\ : IoSpan4Mux
    port map (
            O => \N__36055\,
            I => \N__36052\
        );

    \I__8405\ : Span4Mux_s1_h
    port map (
            O => \N__36052\,
            I => \N__36049\
        );

    \I__8404\ : Span4Mux_h
    port map (
            O => \N__36049\,
            I => \N__36046\
        );

    \I__8403\ : Odrv4
    port map (
            O => \N__36046\,
            I => \N_1048_i\
        );

    \I__8402\ : InMux
    port map (
            O => \N__36043\,
            I => \N__36040\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__36040\,
            I => \N__36037\
        );

    \I__8400\ : Span4Mux_h
    port map (
            O => \N__36037\,
            I => \N__36034\
        );

    \I__8399\ : Span4Mux_v
    port map (
            O => \N__36034\,
            I => \N__36031\
        );

    \I__8398\ : Odrv4
    port map (
            O => \N__36031\,
            I => \this_spr_ram.mem_out_bus5_1\
        );

    \I__8397\ : InMux
    port map (
            O => \N__36028\,
            I => \N__36025\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__36025\,
            I => \N__36022\
        );

    \I__8395\ : Span4Mux_v
    port map (
            O => \N__36022\,
            I => \N__36019\
        );

    \I__8394\ : Span4Mux_v
    port map (
            O => \N__36019\,
            I => \N__36016\
        );

    \I__8393\ : Odrv4
    port map (
            O => \N__36016\,
            I => \this_spr_ram.mem_out_bus1_1\
        );

    \I__8392\ : InMux
    port map (
            O => \N__36013\,
            I => \N__36010\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__36010\,
            I => \N__36007\
        );

    \I__8390\ : Span4Mux_v
    port map (
            O => \N__36007\,
            I => \N__36004\
        );

    \I__8389\ : Odrv4
    port map (
            O => \N__36004\,
            I => \this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0\
        );

    \I__8388\ : InMux
    port map (
            O => \N__36001\,
            I => \N__35995\
        );

    \I__8387\ : InMux
    port map (
            O => \N__36000\,
            I => \N__35995\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__35995\,
            I => \this_ppu.N_1257\
        );

    \I__8385\ : InMux
    port map (
            O => \N__35992\,
            I => \N__35989\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__35989\,
            I => \N__35985\
        );

    \I__8383\ : InMux
    port map (
            O => \N__35988\,
            I => \N__35982\
        );

    \I__8382\ : Span4Mux_v
    port map (
            O => \N__35985\,
            I => \N__35977\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__35982\,
            I => \N__35977\
        );

    \I__8380\ : Span4Mux_h
    port map (
            O => \N__35977\,
            I => \N__35973\
        );

    \I__8379\ : InMux
    port map (
            O => \N__35976\,
            I => \N__35970\
        );

    \I__8378\ : Odrv4
    port map (
            O => \N__35973\,
            I => \this_ppu.N_1322\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__35970\,
            I => \this_ppu.N_1322\
        );

    \I__8376\ : InMux
    port map (
            O => \N__35965\,
            I => \N__35961\
        );

    \I__8375\ : InMux
    port map (
            O => \N__35964\,
            I => \N__35957\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__35961\,
            I => \N__35954\
        );

    \I__8373\ : InMux
    port map (
            O => \N__35960\,
            I => \N__35951\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__35957\,
            I => \N__35946\
        );

    \I__8371\ : Span4Mux_h
    port map (
            O => \N__35954\,
            I => \N__35943\
        );

    \I__8370\ : LocalMux
    port map (
            O => \N__35951\,
            I => \N__35940\
        );

    \I__8369\ : InMux
    port map (
            O => \N__35950\,
            I => \N__35937\
        );

    \I__8368\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35933\
        );

    \I__8367\ : Span4Mux_v
    port map (
            O => \N__35946\,
            I => \N__35930\
        );

    \I__8366\ : Span4Mux_v
    port map (
            O => \N__35943\,
            I => \N__35925\
        );

    \I__8365\ : Span4Mux_h
    port map (
            O => \N__35940\,
            I => \N__35925\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__35937\,
            I => \N__35922\
        );

    \I__8363\ : InMux
    port map (
            O => \N__35936\,
            I => \N__35919\
        );

    \I__8362\ : LocalMux
    port map (
            O => \N__35933\,
            I => \N__35915\
        );

    \I__8361\ : Span4Mux_v
    port map (
            O => \N__35930\,
            I => \N__35911\
        );

    \I__8360\ : Span4Mux_v
    port map (
            O => \N__35925\,
            I => \N__35906\
        );

    \I__8359\ : Span4Mux_h
    port map (
            O => \N__35922\,
            I => \N__35906\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__35919\,
            I => \N__35903\
        );

    \I__8357\ : InMux
    port map (
            O => \N__35918\,
            I => \N__35900\
        );

    \I__8356\ : Span4Mux_h
    port map (
            O => \N__35915\,
            I => \N__35897\
        );

    \I__8355\ : InMux
    port map (
            O => \N__35914\,
            I => \N__35894\
        );

    \I__8354\ : Sp12to4
    port map (
            O => \N__35911\,
            I => \N__35891\
        );

    \I__8353\ : Span4Mux_v
    port map (
            O => \N__35906\,
            I => \N__35886\
        );

    \I__8352\ : Span4Mux_h
    port map (
            O => \N__35903\,
            I => \N__35886\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__35900\,
            I => \N__35883\
        );

    \I__8350\ : Span4Mux_v
    port map (
            O => \N__35897\,
            I => \N__35878\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__35894\,
            I => \N__35878\
        );

    \I__8348\ : Span12Mux_h
    port map (
            O => \N__35891\,
            I => \N__35875\
        );

    \I__8347\ : Span4Mux_v
    port map (
            O => \N__35886\,
            I => \N__35868\
        );

    \I__8346\ : Span4Mux_h
    port map (
            O => \N__35883\,
            I => \N__35868\
        );

    \I__8345\ : Span4Mux_h
    port map (
            O => \N__35878\,
            I => \N__35868\
        );

    \I__8344\ : Odrv12
    port map (
            O => \N__35875\,
            I => \M_this_spr_ram_write_data_1\
        );

    \I__8343\ : Odrv4
    port map (
            O => \N__35868\,
            I => \M_this_spr_ram_write_data_1\
        );

    \I__8342\ : IoInMux
    port map (
            O => \N__35863\,
            I => \N__35860\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__35860\,
            I => \N__35857\
        );

    \I__8340\ : Span4Mux_s3_h
    port map (
            O => \N__35857\,
            I => \N__35854\
        );

    \I__8339\ : Span4Mux_h
    port map (
            O => \N__35854\,
            I => \N__35851\
        );

    \I__8338\ : Span4Mux_h
    port map (
            O => \N__35851\,
            I => \N__35848\
        );

    \I__8337\ : Sp12to4
    port map (
            O => \N__35848\,
            I => \N__35842\
        );

    \I__8336\ : InMux
    port map (
            O => \N__35847\,
            I => \N__35834\
        );

    \I__8335\ : InMux
    port map (
            O => \N__35846\,
            I => \N__35834\
        );

    \I__8334\ : InMux
    port map (
            O => \N__35845\,
            I => \N__35831\
        );

    \I__8333\ : Span12Mux_v
    port map (
            O => \N__35842\,
            I => \N__35827\
        );

    \I__8332\ : InMux
    port map (
            O => \N__35841\,
            I => \N__35822\
        );

    \I__8331\ : InMux
    port map (
            O => \N__35840\,
            I => \N__35822\
        );

    \I__8330\ : InMux
    port map (
            O => \N__35839\,
            I => \N__35819\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__35834\,
            I => \N__35814\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__35831\,
            I => \N__35814\
        );

    \I__8327\ : InMux
    port map (
            O => \N__35830\,
            I => \N__35811\
        );

    \I__8326\ : Odrv12
    port map (
            O => \N__35827\,
            I => led_c_1
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__35822\,
            I => led_c_1
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__35819\,
            I => led_c_1
        );

    \I__8323\ : Odrv4
    port map (
            O => \N__35814\,
            I => led_c_1
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__35811\,
            I => led_c_1
        );

    \I__8321\ : CascadeMux
    port map (
            O => \N__35800\,
            I => \N_1416_cascade_\
        );

    \I__8320\ : CascadeMux
    port map (
            O => \N__35797\,
            I => \N__35794\
        );

    \I__8319\ : InMux
    port map (
            O => \N__35794\,
            I => \N__35788\
        );

    \I__8318\ : InMux
    port map (
            O => \N__35793\,
            I => \N__35788\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__35788\,
            I => \N_1151_3\
        );

    \I__8316\ : InMux
    port map (
            O => \N__35785\,
            I => \N__35778\
        );

    \I__8315\ : InMux
    port map (
            O => \N__35784\,
            I => \N__35774\
        );

    \I__8314\ : InMux
    port map (
            O => \N__35783\,
            I => \N__35770\
        );

    \I__8313\ : InMux
    port map (
            O => \N__35782\,
            I => \N__35767\
        );

    \I__8312\ : InMux
    port map (
            O => \N__35781\,
            I => \N__35764\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__35778\,
            I => \N__35760\
        );

    \I__8310\ : InMux
    port map (
            O => \N__35777\,
            I => \N__35757\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__35774\,
            I => \N__35754\
        );

    \I__8308\ : InMux
    port map (
            O => \N__35773\,
            I => \N__35751\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__35770\,
            I => \N__35748\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__35767\,
            I => \N__35743\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__35764\,
            I => \N__35743\
        );

    \I__8304\ : InMux
    port map (
            O => \N__35763\,
            I => \N__35740\
        );

    \I__8303\ : Span4Mux_h
    port map (
            O => \N__35760\,
            I => \N__35733\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__35757\,
            I => \N__35733\
        );

    \I__8301\ : Span4Mux_v
    port map (
            O => \N__35754\,
            I => \N__35733\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__35751\,
            I => \N__35726\
        );

    \I__8299\ : Span4Mux_v
    port map (
            O => \N__35748\,
            I => \N__35726\
        );

    \I__8298\ : Span4Mux_v
    port map (
            O => \N__35743\,
            I => \N__35726\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__35740\,
            I => \this_ppu.N_787_0\
        );

    \I__8296\ : Odrv4
    port map (
            O => \N__35733\,
            I => \this_ppu.N_787_0\
        );

    \I__8295\ : Odrv4
    port map (
            O => \N__35726\,
            I => \this_ppu.N_787_0\
        );

    \I__8294\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35716\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__35716\,
            I => \this_ppu.M_this_state_q_srsts_0_0_a2_1_sxZ0Z_0\
        );

    \I__8292\ : CascadeMux
    port map (
            O => \N__35713\,
            I => \N__35706\
        );

    \I__8291\ : InMux
    port map (
            O => \N__35712\,
            I => \N__35698\
        );

    \I__8290\ : InMux
    port map (
            O => \N__35711\,
            I => \N__35698\
        );

    \I__8289\ : InMux
    port map (
            O => \N__35710\,
            I => \N__35698\
        );

    \I__8288\ : InMux
    port map (
            O => \N__35709\,
            I => \N__35693\
        );

    \I__8287\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35693\
        );

    \I__8286\ : CascadeMux
    port map (
            O => \N__35705\,
            I => \N__35690\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__35698\,
            I => \N__35685\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__35693\,
            I => \N__35685\
        );

    \I__8283\ : InMux
    port map (
            O => \N__35690\,
            I => \N__35681\
        );

    \I__8282\ : Span4Mux_h
    port map (
            O => \N__35685\,
            I => \N__35678\
        );

    \I__8281\ : InMux
    port map (
            O => \N__35684\,
            I => \N__35675\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__35681\,
            I => \N__35672\
        );

    \I__8279\ : Odrv4
    port map (
            O => \N__35678\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__35675\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__8277\ : Odrv4
    port map (
            O => \N__35672\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__8276\ : InMux
    port map (
            O => \N__35665\,
            I => \N__35660\
        );

    \I__8275\ : InMux
    port map (
            O => \N__35664\,
            I => \N__35657\
        );

    \I__8274\ : InMux
    port map (
            O => \N__35663\,
            I => \N__35653\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__35660\,
            I => \N__35648\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__35657\,
            I => \N__35648\
        );

    \I__8271\ : InMux
    port map (
            O => \N__35656\,
            I => \N__35645\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__35653\,
            I => \N__35642\
        );

    \I__8269\ : Span4Mux_h
    port map (
            O => \N__35648\,
            I => \N__35637\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__35645\,
            I => \N__35637\
        );

    \I__8267\ : Span4Mux_h
    port map (
            O => \N__35642\,
            I => \N__35634\
        );

    \I__8266\ : Odrv4
    port map (
            O => \N__35637\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__8265\ : Odrv4
    port map (
            O => \N__35634\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__8264\ : CascadeMux
    port map (
            O => \N__35629\,
            I => \N__35626\
        );

    \I__8263\ : InMux
    port map (
            O => \N__35626\,
            I => \N__35623\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__35623\,
            I => \N__35620\
        );

    \I__8261\ : Odrv4
    port map (
            O => \N__35620\,
            I => \this_vga_signals.g2_1_0\
        );

    \I__8260\ : CascadeMux
    port map (
            O => \N__35617\,
            I => \N__35612\
        );

    \I__8259\ : CascadeMux
    port map (
            O => \N__35616\,
            I => \N__35605\
        );

    \I__8258\ : InMux
    port map (
            O => \N__35615\,
            I => \N__35595\
        );

    \I__8257\ : InMux
    port map (
            O => \N__35612\,
            I => \N__35595\
        );

    \I__8256\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35595\
        );

    \I__8255\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35592\
        );

    \I__8254\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35587\
        );

    \I__8253\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35587\
        );

    \I__8252\ : InMux
    port map (
            O => \N__35605\,
            I => \N__35582\
        );

    \I__8251\ : InMux
    port map (
            O => \N__35604\,
            I => \N__35582\
        );

    \I__8250\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35577\
        );

    \I__8249\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35577\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__35595\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_4\
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__35592\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_4\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__35587\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_4\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__35582\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_4\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__35577\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_4\
        );

    \I__8243\ : InMux
    port map (
            O => \N__35566\,
            I => \N__35563\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__35563\,
            I => \N__35560\
        );

    \I__8241\ : Odrv12
    port map (
            O => \N__35560\,
            I => \this_vga_signals.mult1_un47_sum_2_1\
        );

    \I__8240\ : InMux
    port map (
            O => \N__35557\,
            I => \N__35554\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__35554\,
            I => \N__35549\
        );

    \I__8238\ : InMux
    port map (
            O => \N__35553\,
            I => \N__35545\
        );

    \I__8237\ : InMux
    port map (
            O => \N__35552\,
            I => \N__35542\
        );

    \I__8236\ : Span4Mux_h
    port map (
            O => \N__35549\,
            I => \N__35539\
        );

    \I__8235\ : InMux
    port map (
            O => \N__35548\,
            I => \N__35536\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__35545\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__35542\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__35539\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__35536\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__8230\ : InMux
    port map (
            O => \N__35527\,
            I => \N__35524\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__35524\,
            I => \this_vga_signals.if_N_7_0_0\
        );

    \I__8228\ : CascadeMux
    port map (
            O => \N__35521\,
            I => \N__35511\
        );

    \I__8227\ : CascadeMux
    port map (
            O => \N__35520\,
            I => \N__35508\
        );

    \I__8226\ : CascadeMux
    port map (
            O => \N__35519\,
            I => \N__35505\
        );

    \I__8225\ : InMux
    port map (
            O => \N__35518\,
            I => \N__35498\
        );

    \I__8224\ : InMux
    port map (
            O => \N__35517\,
            I => \N__35498\
        );

    \I__8223\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35498\
        );

    \I__8222\ : InMux
    port map (
            O => \N__35515\,
            I => \N__35495\
        );

    \I__8221\ : InMux
    port map (
            O => \N__35514\,
            I => \N__35492\
        );

    \I__8220\ : InMux
    port map (
            O => \N__35511\,
            I => \N__35486\
        );

    \I__8219\ : InMux
    port map (
            O => \N__35508\,
            I => \N__35483\
        );

    \I__8218\ : InMux
    port map (
            O => \N__35505\,
            I => \N__35480\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__35498\,
            I => \N__35477\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__35495\,
            I => \N__35472\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__35492\,
            I => \N__35472\
        );

    \I__8214\ : CascadeMux
    port map (
            O => \N__35491\,
            I => \N__35469\
        );

    \I__8213\ : CascadeMux
    port map (
            O => \N__35490\,
            I => \N__35466\
        );

    \I__8212\ : InMux
    port map (
            O => \N__35489\,
            I => \N__35461\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__35486\,
            I => \N__35453\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__35483\,
            I => \N__35453\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__35480\,
            I => \N__35453\
        );

    \I__8208\ : Span4Mux_h
    port map (
            O => \N__35477\,
            I => \N__35448\
        );

    \I__8207\ : Span4Mux_h
    port map (
            O => \N__35472\,
            I => \N__35448\
        );

    \I__8206\ : InMux
    port map (
            O => \N__35469\,
            I => \N__35443\
        );

    \I__8205\ : InMux
    port map (
            O => \N__35466\,
            I => \N__35443\
        );

    \I__8204\ : InMux
    port map (
            O => \N__35465\,
            I => \N__35440\
        );

    \I__8203\ : InMux
    port map (
            O => \N__35464\,
            I => \N__35437\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__35461\,
            I => \N__35434\
        );

    \I__8201\ : InMux
    port map (
            O => \N__35460\,
            I => \N__35431\
        );

    \I__8200\ : Span12Mux_h
    port map (
            O => \N__35453\,
            I => \N__35426\
        );

    \I__8199\ : Sp12to4
    port map (
            O => \N__35448\,
            I => \N__35426\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__35443\,
            I => \N__35423\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__35440\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__35437\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__8195\ : Odrv4
    port map (
            O => \N__35434\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__35431\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__8193\ : Odrv12
    port map (
            O => \N__35426\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__8192\ : Odrv4
    port map (
            O => \N__35423\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__8191\ : InMux
    port map (
            O => \N__35410\,
            I => \N__35402\
        );

    \I__8190\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35393\
        );

    \I__8189\ : InMux
    port map (
            O => \N__35408\,
            I => \N__35393\
        );

    \I__8188\ : InMux
    port map (
            O => \N__35407\,
            I => \N__35387\
        );

    \I__8187\ : InMux
    port map (
            O => \N__35406\,
            I => \N__35387\
        );

    \I__8186\ : CascadeMux
    port map (
            O => \N__35405\,
            I => \N__35381\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__35402\,
            I => \N__35377\
        );

    \I__8184\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35370\
        );

    \I__8183\ : InMux
    port map (
            O => \N__35400\,
            I => \N__35370\
        );

    \I__8182\ : InMux
    port map (
            O => \N__35399\,
            I => \N__35370\
        );

    \I__8181\ : InMux
    port map (
            O => \N__35398\,
            I => \N__35367\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__35393\,
            I => \N__35364\
        );

    \I__8179\ : InMux
    port map (
            O => \N__35392\,
            I => \N__35361\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__35387\,
            I => \N__35358\
        );

    \I__8177\ : InMux
    port map (
            O => \N__35386\,
            I => \N__35353\
        );

    \I__8176\ : InMux
    port map (
            O => \N__35385\,
            I => \N__35353\
        );

    \I__8175\ : InMux
    port map (
            O => \N__35384\,
            I => \N__35346\
        );

    \I__8174\ : InMux
    port map (
            O => \N__35381\,
            I => \N__35346\
        );

    \I__8173\ : InMux
    port map (
            O => \N__35380\,
            I => \N__35346\
        );

    \I__8172\ : Odrv4
    port map (
            O => \N__35377\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__35370\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__35367\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__8169\ : Odrv12
    port map (
            O => \N__35364\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__35361\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__8167\ : Odrv4
    port map (
            O => \N__35358\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__35353\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__35346\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__8164\ : InMux
    port map (
            O => \N__35329\,
            I => \N__35326\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__35326\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_d_0_0\
        );

    \I__8162\ : InMux
    port map (
            O => \N__35323\,
            I => \N__35311\
        );

    \I__8161\ : InMux
    port map (
            O => \N__35322\,
            I => \N__35308\
        );

    \I__8160\ : InMux
    port map (
            O => \N__35321\,
            I => \N__35297\
        );

    \I__8159\ : InMux
    port map (
            O => \N__35320\,
            I => \N__35294\
        );

    \I__8158\ : InMux
    port map (
            O => \N__35319\,
            I => \N__35290\
        );

    \I__8157\ : InMux
    port map (
            O => \N__35318\,
            I => \N__35287\
        );

    \I__8156\ : InMux
    port map (
            O => \N__35317\,
            I => \N__35279\
        );

    \I__8155\ : InMux
    port map (
            O => \N__35316\,
            I => \N__35279\
        );

    \I__8154\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35279\
        );

    \I__8153\ : InMux
    port map (
            O => \N__35314\,
            I => \N__35276\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__35311\,
            I => \N__35271\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__35308\,
            I => \N__35271\
        );

    \I__8150\ : InMux
    port map (
            O => \N__35307\,
            I => \N__35266\
        );

    \I__8149\ : InMux
    port map (
            O => \N__35306\,
            I => \N__35266\
        );

    \I__8148\ : InMux
    port map (
            O => \N__35305\,
            I => \N__35263\
        );

    \I__8147\ : InMux
    port map (
            O => \N__35304\,
            I => \N__35260\
        );

    \I__8146\ : InMux
    port map (
            O => \N__35303\,
            I => \N__35257\
        );

    \I__8145\ : InMux
    port map (
            O => \N__35302\,
            I => \N__35252\
        );

    \I__8144\ : InMux
    port map (
            O => \N__35301\,
            I => \N__35252\
        );

    \I__8143\ : CascadeMux
    port map (
            O => \N__35300\,
            I => \N__35249\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__35297\,
            I => \N__35245\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__35294\,
            I => \N__35242\
        );

    \I__8140\ : CascadeMux
    port map (
            O => \N__35293\,
            I => \N__35237\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__35290\,
            I => \N__35232\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__35287\,
            I => \N__35232\
        );

    \I__8137\ : InMux
    port map (
            O => \N__35286\,
            I => \N__35229\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__35279\,
            I => \N__35220\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__35276\,
            I => \N__35220\
        );

    \I__8134\ : Span4Mux_v
    port map (
            O => \N__35271\,
            I => \N__35220\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__35266\,
            I => \N__35220\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__35263\,
            I => \N__35216\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__35260\,
            I => \N__35211\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__35257\,
            I => \N__35211\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__35252\,
            I => \N__35208\
        );

    \I__8128\ : InMux
    port map (
            O => \N__35249\,
            I => \N__35205\
        );

    \I__8127\ : InMux
    port map (
            O => \N__35248\,
            I => \N__35202\
        );

    \I__8126\ : Span4Mux_v
    port map (
            O => \N__35245\,
            I => \N__35197\
        );

    \I__8125\ : Span4Mux_v
    port map (
            O => \N__35242\,
            I => \N__35197\
        );

    \I__8124\ : InMux
    port map (
            O => \N__35241\,
            I => \N__35190\
        );

    \I__8123\ : InMux
    port map (
            O => \N__35240\,
            I => \N__35190\
        );

    \I__8122\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35190\
        );

    \I__8121\ : Sp12to4
    port map (
            O => \N__35232\,
            I => \N__35185\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__35229\,
            I => \N__35185\
        );

    \I__8119\ : Span4Mux_h
    port map (
            O => \N__35220\,
            I => \N__35182\
        );

    \I__8118\ : InMux
    port map (
            O => \N__35219\,
            I => \N__35179\
        );

    \I__8117\ : Span4Mux_h
    port map (
            O => \N__35216\,
            I => \N__35170\
        );

    \I__8116\ : Span4Mux_h
    port map (
            O => \N__35211\,
            I => \N__35170\
        );

    \I__8115\ : Span4Mux_h
    port map (
            O => \N__35208\,
            I => \N__35170\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__35205\,
            I => \N__35170\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__35202\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__8112\ : Odrv4
    port map (
            O => \N__35197\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__35190\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__8110\ : Odrv12
    port map (
            O => \N__35185\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__8109\ : Odrv4
    port map (
            O => \N__35182\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__35179\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__8107\ : Odrv4
    port map (
            O => \N__35170\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__8106\ : CascadeMux
    port map (
            O => \N__35155\,
            I => \N__35147\
        );

    \I__8105\ : CascadeMux
    port map (
            O => \N__35154\,
            I => \N__35143\
        );

    \I__8104\ : InMux
    port map (
            O => \N__35153\,
            I => \N__35138\
        );

    \I__8103\ : InMux
    port map (
            O => \N__35152\,
            I => \N__35130\
        );

    \I__8102\ : InMux
    port map (
            O => \N__35151\,
            I => \N__35127\
        );

    \I__8101\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35124\
        );

    \I__8100\ : InMux
    port map (
            O => \N__35147\,
            I => \N__35121\
        );

    \I__8099\ : InMux
    port map (
            O => \N__35146\,
            I => \N__35118\
        );

    \I__8098\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35115\
        );

    \I__8097\ : InMux
    port map (
            O => \N__35142\,
            I => \N__35110\
        );

    \I__8096\ : InMux
    port map (
            O => \N__35141\,
            I => \N__35110\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__35138\,
            I => \N__35107\
        );

    \I__8094\ : InMux
    port map (
            O => \N__35137\,
            I => \N__35104\
        );

    \I__8093\ : CascadeMux
    port map (
            O => \N__35136\,
            I => \N__35101\
        );

    \I__8092\ : CascadeMux
    port map (
            O => \N__35135\,
            I => \N__35096\
        );

    \I__8091\ : InMux
    port map (
            O => \N__35134\,
            I => \N__35093\
        );

    \I__8090\ : CascadeMux
    port map (
            O => \N__35133\,
            I => \N__35090\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__35130\,
            I => \N__35086\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__35127\,
            I => \N__35079\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__35124\,
            I => \N__35079\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__35121\,
            I => \N__35079\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__35118\,
            I => \N__35076\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__35115\,
            I => \N__35072\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__35110\,
            I => \N__35065\
        );

    \I__8082\ : Span4Mux_v
    port map (
            O => \N__35107\,
            I => \N__35065\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__35104\,
            I => \N__35065\
        );

    \I__8080\ : InMux
    port map (
            O => \N__35101\,
            I => \N__35060\
        );

    \I__8079\ : InMux
    port map (
            O => \N__35100\,
            I => \N__35060\
        );

    \I__8078\ : InMux
    port map (
            O => \N__35099\,
            I => \N__35057\
        );

    \I__8077\ : InMux
    port map (
            O => \N__35096\,
            I => \N__35054\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__35093\,
            I => \N__35051\
        );

    \I__8075\ : InMux
    port map (
            O => \N__35090\,
            I => \N__35046\
        );

    \I__8074\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35046\
        );

    \I__8073\ : Span4Mux_v
    port map (
            O => \N__35086\,
            I => \N__35039\
        );

    \I__8072\ : Span4Mux_h
    port map (
            O => \N__35079\,
            I => \N__35039\
        );

    \I__8071\ : Span4Mux_v
    port map (
            O => \N__35076\,
            I => \N__35039\
        );

    \I__8070\ : InMux
    port map (
            O => \N__35075\,
            I => \N__35036\
        );

    \I__8069\ : Span4Mux_h
    port map (
            O => \N__35072\,
            I => \N__35029\
        );

    \I__8068\ : Span4Mux_h
    port map (
            O => \N__35065\,
            I => \N__35029\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__35060\,
            I => \N__35029\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__35057\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__35054\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__8064\ : Odrv4
    port map (
            O => \N__35051\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__35046\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__8062\ : Odrv4
    port map (
            O => \N__35039\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__35036\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__8060\ : Odrv4
    port map (
            O => \N__35029\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__8059\ : InMux
    port map (
            O => \N__35014\,
            I => \N__35009\
        );

    \I__8058\ : CascadeMux
    port map (
            O => \N__35013\,
            I => \N__35006\
        );

    \I__8057\ : InMux
    port map (
            O => \N__35012\,
            I => \N__35001\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__35009\,
            I => \N__34996\
        );

    \I__8055\ : InMux
    port map (
            O => \N__35006\,
            I => \N__34987\
        );

    \I__8054\ : CascadeMux
    port map (
            O => \N__35005\,
            I => \N__34983\
        );

    \I__8053\ : InMux
    port map (
            O => \N__35004\,
            I => \N__34980\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__35001\,
            I => \N__34977\
        );

    \I__8051\ : InMux
    port map (
            O => \N__35000\,
            I => \N__34974\
        );

    \I__8050\ : CascadeMux
    port map (
            O => \N__34999\,
            I => \N__34968\
        );

    \I__8049\ : Span4Mux_h
    port map (
            O => \N__34996\,
            I => \N__34963\
        );

    \I__8048\ : InMux
    port map (
            O => \N__34995\,
            I => \N__34960\
        );

    \I__8047\ : InMux
    port map (
            O => \N__34994\,
            I => \N__34955\
        );

    \I__8046\ : InMux
    port map (
            O => \N__34993\,
            I => \N__34955\
        );

    \I__8045\ : InMux
    port map (
            O => \N__34992\,
            I => \N__34948\
        );

    \I__8044\ : InMux
    port map (
            O => \N__34991\,
            I => \N__34948\
        );

    \I__8043\ : InMux
    port map (
            O => \N__34990\,
            I => \N__34948\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__34987\,
            I => \N__34939\
        );

    \I__8041\ : InMux
    port map (
            O => \N__34986\,
            I => \N__34935\
        );

    \I__8040\ : InMux
    port map (
            O => \N__34983\,
            I => \N__34932\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__34980\,
            I => \N__34929\
        );

    \I__8038\ : Span4Mux_h
    port map (
            O => \N__34977\,
            I => \N__34924\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__34974\,
            I => \N__34924\
        );

    \I__8036\ : InMux
    port map (
            O => \N__34973\,
            I => \N__34921\
        );

    \I__8035\ : InMux
    port map (
            O => \N__34972\,
            I => \N__34916\
        );

    \I__8034\ : InMux
    port map (
            O => \N__34971\,
            I => \N__34916\
        );

    \I__8033\ : InMux
    port map (
            O => \N__34968\,
            I => \N__34913\
        );

    \I__8032\ : InMux
    port map (
            O => \N__34967\,
            I => \N__34908\
        );

    \I__8031\ : InMux
    port map (
            O => \N__34966\,
            I => \N__34908\
        );

    \I__8030\ : Span4Mux_h
    port map (
            O => \N__34963\,
            I => \N__34901\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__34960\,
            I => \N__34901\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__34955\,
            I => \N__34901\
        );

    \I__8027\ : LocalMux
    port map (
            O => \N__34948\,
            I => \N__34898\
        );

    \I__8026\ : InMux
    port map (
            O => \N__34947\,
            I => \N__34894\
        );

    \I__8025\ : CascadeMux
    port map (
            O => \N__34946\,
            I => \N__34891\
        );

    \I__8024\ : CascadeMux
    port map (
            O => \N__34945\,
            I => \N__34888\
        );

    \I__8023\ : CascadeMux
    port map (
            O => \N__34944\,
            I => \N__34885\
        );

    \I__8022\ : CascadeMux
    port map (
            O => \N__34943\,
            I => \N__34882\
        );

    \I__8021\ : CascadeMux
    port map (
            O => \N__34942\,
            I => \N__34876\
        );

    \I__8020\ : Span4Mux_v
    port map (
            O => \N__34939\,
            I => \N__34873\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__34938\,
            I => \N__34870\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__34935\,
            I => \N__34865\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__34932\,
            I => \N__34865\
        );

    \I__8016\ : Span4Mux_v
    port map (
            O => \N__34929\,
            I => \N__34858\
        );

    \I__8015\ : Span4Mux_v
    port map (
            O => \N__34924\,
            I => \N__34858\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__34921\,
            I => \N__34858\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__34916\,
            I => \N__34855\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__34913\,
            I => \N__34846\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__34908\,
            I => \N__34846\
        );

    \I__8010\ : Span4Mux_h
    port map (
            O => \N__34901\,
            I => \N__34846\
        );

    \I__8009\ : Span4Mux_v
    port map (
            O => \N__34898\,
            I => \N__34846\
        );

    \I__8008\ : CascadeMux
    port map (
            O => \N__34897\,
            I => \N__34843\
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__34894\,
            I => \N__34839\
        );

    \I__8006\ : InMux
    port map (
            O => \N__34891\,
            I => \N__34836\
        );

    \I__8005\ : InMux
    port map (
            O => \N__34888\,
            I => \N__34831\
        );

    \I__8004\ : InMux
    port map (
            O => \N__34885\,
            I => \N__34831\
        );

    \I__8003\ : InMux
    port map (
            O => \N__34882\,
            I => \N__34826\
        );

    \I__8002\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34826\
        );

    \I__8001\ : InMux
    port map (
            O => \N__34880\,
            I => \N__34823\
        );

    \I__8000\ : InMux
    port map (
            O => \N__34879\,
            I => \N__34820\
        );

    \I__7999\ : InMux
    port map (
            O => \N__34876\,
            I => \N__34817\
        );

    \I__7998\ : Span4Mux_h
    port map (
            O => \N__34873\,
            I => \N__34814\
        );

    \I__7997\ : InMux
    port map (
            O => \N__34870\,
            I => \N__34811\
        );

    \I__7996\ : Span4Mux_v
    port map (
            O => \N__34865\,
            I => \N__34804\
        );

    \I__7995\ : Span4Mux_h
    port map (
            O => \N__34858\,
            I => \N__34804\
        );

    \I__7994\ : Span4Mux_v
    port map (
            O => \N__34855\,
            I => \N__34804\
        );

    \I__7993\ : Span4Mux_h
    port map (
            O => \N__34846\,
            I => \N__34801\
        );

    \I__7992\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34796\
        );

    \I__7991\ : InMux
    port map (
            O => \N__34842\,
            I => \N__34796\
        );

    \I__7990\ : Span12Mux_v
    port map (
            O => \N__34839\,
            I => \N__34787\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__34836\,
            I => \N__34787\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__34831\,
            I => \N__34787\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__34826\,
            I => \N__34787\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__34823\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__34820\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__34817\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__7983\ : Odrv4
    port map (
            O => \N__34814\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__34811\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__7981\ : Odrv4
    port map (
            O => \N__34804\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__7980\ : Odrv4
    port map (
            O => \N__34801\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__34796\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__7978\ : Odrv12
    port map (
            O => \N__34787\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__7977\ : CascadeMux
    port map (
            O => \N__34768\,
            I => \N__34765\
        );

    \I__7976\ : InMux
    port map (
            O => \N__34765\,
            I => \N__34762\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__34762\,
            I => \N__34759\
        );

    \I__7974\ : Span4Mux_v
    port map (
            O => \N__34759\,
            I => \N__34755\
        );

    \I__7973\ : InMux
    port map (
            O => \N__34758\,
            I => \N__34752\
        );

    \I__7972\ : Span4Mux_h
    port map (
            O => \N__34755\,
            I => \N__34739\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__34752\,
            I => \N__34739\
        );

    \I__7970\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34736\
        );

    \I__7969\ : InMux
    port map (
            O => \N__34750\,
            I => \N__34732\
        );

    \I__7968\ : InMux
    port map (
            O => \N__34749\,
            I => \N__34729\
        );

    \I__7967\ : InMux
    port map (
            O => \N__34748\,
            I => \N__34726\
        );

    \I__7966\ : InMux
    port map (
            O => \N__34747\,
            I => \N__34723\
        );

    \I__7965\ : InMux
    port map (
            O => \N__34746\,
            I => \N__34720\
        );

    \I__7964\ : InMux
    port map (
            O => \N__34745\,
            I => \N__34717\
        );

    \I__7963\ : InMux
    port map (
            O => \N__34744\,
            I => \N__34713\
        );

    \I__7962\ : Span4Mux_v
    port map (
            O => \N__34739\,
            I => \N__34710\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__34736\,
            I => \N__34707\
        );

    \I__7960\ : InMux
    port map (
            O => \N__34735\,
            I => \N__34700\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__34732\,
            I => \N__34697\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__34729\,
            I => \N__34692\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__34726\,
            I => \N__34692\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__34723\,
            I => \N__34685\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__34720\,
            I => \N__34685\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__34717\,
            I => \N__34685\
        );

    \I__7953\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34682\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__34713\,
            I => \N__34679\
        );

    \I__7951\ : Span4Mux_h
    port map (
            O => \N__34710\,
            I => \N__34676\
        );

    \I__7950\ : Span12Mux_h
    port map (
            O => \N__34707\,
            I => \N__34673\
        );

    \I__7949\ : InMux
    port map (
            O => \N__34706\,
            I => \N__34670\
        );

    \I__7948\ : InMux
    port map (
            O => \N__34705\,
            I => \N__34667\
        );

    \I__7947\ : InMux
    port map (
            O => \N__34704\,
            I => \N__34662\
        );

    \I__7946\ : InMux
    port map (
            O => \N__34703\,
            I => \N__34662\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__34700\,
            I => \N__34651\
        );

    \I__7944\ : Span4Mux_h
    port map (
            O => \N__34697\,
            I => \N__34651\
        );

    \I__7943\ : Span4Mux_h
    port map (
            O => \N__34692\,
            I => \N__34651\
        );

    \I__7942\ : Span4Mux_v
    port map (
            O => \N__34685\,
            I => \N__34651\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__34682\,
            I => \N__34651\
        );

    \I__7940\ : Span4Mux_v
    port map (
            O => \N__34679\,
            I => \N__34648\
        );

    \I__7939\ : Odrv4
    port map (
            O => \N__34676\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__7938\ : Odrv12
    port map (
            O => \N__34673\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__34670\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__34667\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__34662\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__7934\ : Odrv4
    port map (
            O => \N__34651\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__7933\ : Odrv4
    port map (
            O => \N__34648\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__7932\ : CascadeMux
    port map (
            O => \N__34633\,
            I => \N__34630\
        );

    \I__7931\ : InMux
    port map (
            O => \N__34630\,
            I => \N__34627\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__34627\,
            I => \this_vga_signals.vaddress_0_0_7\
        );

    \I__7929\ : CascadeMux
    port map (
            O => \N__34624\,
            I => \N__34621\
        );

    \I__7928\ : InMux
    port map (
            O => \N__34621\,
            I => \N__34618\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__34618\,
            I => \N__34615\
        );

    \I__7926\ : Span4Mux_h
    port map (
            O => \N__34615\,
            I => \N__34611\
        );

    \I__7925\ : CascadeMux
    port map (
            O => \N__34614\,
            I => \N__34608\
        );

    \I__7924\ : Span4Mux_h
    port map (
            O => \N__34611\,
            I => \N__34605\
        );

    \I__7923\ : InMux
    port map (
            O => \N__34608\,
            I => \N__34602\
        );

    \I__7922\ : Odrv4
    port map (
            O => \N__34605\,
            I => \M_this_scroll_qZ0Z_6\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__34602\,
            I => \M_this_scroll_qZ0Z_6\
        );

    \I__7920\ : InMux
    port map (
            O => \N__34597\,
            I => \N__34594\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__34594\,
            I => \N__34591\
        );

    \I__7918\ : Span4Mux_h
    port map (
            O => \N__34591\,
            I => \N__34588\
        );

    \I__7917\ : Span4Mux_h
    port map (
            O => \N__34588\,
            I => \N__34585\
        );

    \I__7916\ : Odrv4
    port map (
            O => \N__34585\,
            I => \this_ppu.M_screen_y_q_esr_RNILD7F7Z0Z_6\
        );

    \I__7915\ : InMux
    port map (
            O => \N__34582\,
            I => \N__34579\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__34579\,
            I => \N__34573\
        );

    \I__7913\ : InMux
    port map (
            O => \N__34578\,
            I => \N__34570\
        );

    \I__7912\ : InMux
    port map (
            O => \N__34577\,
            I => \N__34567\
        );

    \I__7911\ : InMux
    port map (
            O => \N__34576\,
            I => \N__34562\
        );

    \I__7910\ : Span4Mux_s3_v
    port map (
            O => \N__34573\,
            I => \N__34557\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__34570\,
            I => \N__34557\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__34567\,
            I => \N__34554\
        );

    \I__7907\ : InMux
    port map (
            O => \N__34566\,
            I => \N__34550\
        );

    \I__7906\ : InMux
    port map (
            O => \N__34565\,
            I => \N__34547\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__34562\,
            I => \N__34544\
        );

    \I__7904\ : Span4Mux_v
    port map (
            O => \N__34557\,
            I => \N__34541\
        );

    \I__7903\ : Span4Mux_h
    port map (
            O => \N__34554\,
            I => \N__34538\
        );

    \I__7902\ : InMux
    port map (
            O => \N__34553\,
            I => \N__34535\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__34550\,
            I => \N__34532\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__34547\,
            I => \N__34529\
        );

    \I__7899\ : Span12Mux_s10_h
    port map (
            O => \N__34544\,
            I => \N__34525\
        );

    \I__7898\ : Sp12to4
    port map (
            O => \N__34541\,
            I => \N__34522\
        );

    \I__7897\ : Sp12to4
    port map (
            O => \N__34538\,
            I => \N__34519\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__34535\,
            I => \N__34516\
        );

    \I__7895\ : Span4Mux_v
    port map (
            O => \N__34532\,
            I => \N__34511\
        );

    \I__7894\ : Span4Mux_h
    port map (
            O => \N__34529\,
            I => \N__34511\
        );

    \I__7893\ : InMux
    port map (
            O => \N__34528\,
            I => \N__34508\
        );

    \I__7892\ : Span12Mux_v
    port map (
            O => \N__34525\,
            I => \N__34505\
        );

    \I__7891\ : Span12Mux_h
    port map (
            O => \N__34522\,
            I => \N__34498\
        );

    \I__7890\ : Span12Mux_v
    port map (
            O => \N__34519\,
            I => \N__34498\
        );

    \I__7889\ : Span12Mux_s10_h
    port map (
            O => \N__34516\,
            I => \N__34498\
        );

    \I__7888\ : Span4Mux_v
    port map (
            O => \N__34511\,
            I => \N__34493\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__34508\,
            I => \N__34493\
        );

    \I__7886\ : Odrv12
    port map (
            O => \N__34505\,
            I => \M_this_spr_ram_write_data_3\
        );

    \I__7885\ : Odrv12
    port map (
            O => \N__34498\,
            I => \M_this_spr_ram_write_data_3\
        );

    \I__7884\ : Odrv4
    port map (
            O => \N__34493\,
            I => \M_this_spr_ram_write_data_3\
        );

    \I__7883\ : InMux
    port map (
            O => \N__34486\,
            I => \N__34483\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__34483\,
            I => \N__34480\
        );

    \I__7881\ : Odrv4
    port map (
            O => \N__34480\,
            I => \this_ppu.M_this_state_q_srsts_0_0_a2_1_xZ0Z_0\
        );

    \I__7880\ : InMux
    port map (
            O => \N__34477\,
            I => \N__34473\
        );

    \I__7879\ : InMux
    port map (
            O => \N__34476\,
            I => \N__34470\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__34473\,
            I => \N__34464\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__34470\,
            I => \N__34464\
        );

    \I__7876\ : InMux
    port map (
            O => \N__34469\,
            I => \N__34461\
        );

    \I__7875\ : Span4Mux_v
    port map (
            O => \N__34464\,
            I => \N__34458\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__34461\,
            I => \N__34455\
        );

    \I__7873\ : Span4Mux_h
    port map (
            O => \N__34458\,
            I => \N__34451\
        );

    \I__7872\ : Span12Mux_h
    port map (
            O => \N__34455\,
            I => \N__34448\
        );

    \I__7871\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34445\
        );

    \I__7870\ : Odrv4
    port map (
            O => \N__34451\,
            I => \this_ppu.N_798_0\
        );

    \I__7869\ : Odrv12
    port map (
            O => \N__34448\,
            I => \this_ppu.N_798_0\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__34445\,
            I => \this_ppu.N_798_0\
        );

    \I__7867\ : InMux
    port map (
            O => \N__34438\,
            I => \N__34434\
        );

    \I__7866\ : InMux
    port map (
            O => \N__34437\,
            I => \N__34431\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__34434\,
            I => \N__34427\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__34431\,
            I => \N__34424\
        );

    \I__7863\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34421\
        );

    \I__7862\ : Span4Mux_v
    port map (
            O => \N__34427\,
            I => \N__34418\
        );

    \I__7861\ : Span4Mux_v
    port map (
            O => \N__34424\,
            I => \N__34413\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__34421\,
            I => \N__34413\
        );

    \I__7859\ : Span4Mux_h
    port map (
            O => \N__34418\,
            I => \N__34408\
        );

    \I__7858\ : Span4Mux_h
    port map (
            O => \N__34413\,
            I => \N__34408\
        );

    \I__7857\ : Odrv4
    port map (
            O => \N__34408\,
            I => \this_ppu.N_1426\
        );

    \I__7856\ : InMux
    port map (
            O => \N__34405\,
            I => \N__34402\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__34402\,
            I => \N__34399\
        );

    \I__7854\ : Span4Mux_h
    port map (
            O => \N__34399\,
            I => \N__34396\
        );

    \I__7853\ : Span4Mux_h
    port map (
            O => \N__34396\,
            I => \N__34393\
        );

    \I__7852\ : Span4Mux_h
    port map (
            O => \N__34393\,
            I => \N__34390\
        );

    \I__7851\ : Span4Mux_h
    port map (
            O => \N__34390\,
            I => \N__34387\
        );

    \I__7850\ : Odrv4
    port map (
            O => \N__34387\,
            I => \M_this_ppu_vram_data_3\
        );

    \I__7849\ : InMux
    port map (
            O => \N__34384\,
            I => \N__34381\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__34381\,
            I => \M_this_spr_ram_read_data_2\
        );

    \I__7847\ : CascadeMux
    port map (
            O => \N__34378\,
            I => \M_this_spr_ram_read_data_1_cascade_\
        );

    \I__7846\ : InMux
    port map (
            O => \N__34375\,
            I => \N__34371\
        );

    \I__7845\ : InMux
    port map (
            O => \N__34374\,
            I => \N__34365\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__34371\,
            I => \N__34362\
        );

    \I__7843\ : InMux
    port map (
            O => \N__34370\,
            I => \N__34357\
        );

    \I__7842\ : InMux
    port map (
            O => \N__34369\,
            I => \N__34357\
        );

    \I__7841\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34354\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__34365\,
            I => \N__34351\
        );

    \I__7839\ : Span12Mux_h
    port map (
            O => \N__34362\,
            I => \N__34348\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__34357\,
            I => \N__34341\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__34354\,
            I => \N__34341\
        );

    \I__7836\ : Span12Mux_v
    port map (
            O => \N__34351\,
            I => \N__34341\
        );

    \I__7835\ : Odrv12
    port map (
            O => \N__34348\,
            I => \this_ppu.N_1000_0\
        );

    \I__7834\ : Odrv12
    port map (
            O => \N__34341\,
            I => \this_ppu.N_1000_0\
        );

    \I__7833\ : InMux
    port map (
            O => \N__34336\,
            I => \N__34333\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__34333\,
            I => \M_this_spr_ram_read_data_1\
        );

    \I__7831\ : InMux
    port map (
            O => \N__34330\,
            I => \N__34327\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__34327\,
            I => \N__34324\
        );

    \I__7829\ : Span4Mux_v
    port map (
            O => \N__34324\,
            I => \N__34321\
        );

    \I__7828\ : Span4Mux_h
    port map (
            O => \N__34321\,
            I => \N__34318\
        );

    \I__7827\ : Sp12to4
    port map (
            O => \N__34318\,
            I => \N__34315\
        );

    \I__7826\ : Odrv12
    port map (
            O => \N__34315\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__7825\ : InMux
    port map (
            O => \N__34312\,
            I => \N__34309\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__34309\,
            I => \this_spr_ram.mem_mem_1_0_RNIMA1GZ0\
        );

    \I__7823\ : InMux
    port map (
            O => \N__34306\,
            I => \N__34303\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__34303\,
            I => \N__34300\
        );

    \I__7821\ : Span4Mux_h
    port map (
            O => \N__34300\,
            I => \N__34297\
        );

    \I__7820\ : Span4Mux_h
    port map (
            O => \N__34297\,
            I => \N__34293\
        );

    \I__7819\ : InMux
    port map (
            O => \N__34296\,
            I => \N__34290\
        );

    \I__7818\ : Odrv4
    port map (
            O => \N__34293\,
            I => \M_this_spr_ram_read_data_0\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__34290\,
            I => \M_this_spr_ram_read_data_0\
        );

    \I__7816\ : InMux
    port map (
            O => \N__34285\,
            I => \N__34281\
        );

    \I__7815\ : InMux
    port map (
            O => \N__34284\,
            I => \N__34278\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__34281\,
            I => \N__34274\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__34278\,
            I => \N__34271\
        );

    \I__7812\ : InMux
    port map (
            O => \N__34277\,
            I => \N__34268\
        );

    \I__7811\ : Span4Mux_h
    port map (
            O => \N__34274\,
            I => \N__34265\
        );

    \I__7810\ : Span4Mux_v
    port map (
            O => \N__34271\,
            I => \N__34262\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__34268\,
            I => \N__34259\
        );

    \I__7808\ : Odrv4
    port map (
            O => \N__34265\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__7807\ : Odrv4
    port map (
            O => \N__34262\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__7806\ : Odrv4
    port map (
            O => \N__34259\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__7805\ : CEMux
    port map (
            O => \N__34252\,
            I => \N__34231\
        );

    \I__7804\ : CEMux
    port map (
            O => \N__34251\,
            I => \N__34231\
        );

    \I__7803\ : CEMux
    port map (
            O => \N__34250\,
            I => \N__34231\
        );

    \I__7802\ : CEMux
    port map (
            O => \N__34249\,
            I => \N__34231\
        );

    \I__7801\ : CEMux
    port map (
            O => \N__34248\,
            I => \N__34231\
        );

    \I__7800\ : CEMux
    port map (
            O => \N__34247\,
            I => \N__34231\
        );

    \I__7799\ : CEMux
    port map (
            O => \N__34246\,
            I => \N__34231\
        );

    \I__7798\ : GlobalMux
    port map (
            O => \N__34231\,
            I => \N__34228\
        );

    \I__7797\ : gio2CtrlBuf
    port map (
            O => \N__34228\,
            I => \this_vga_signals.N_1307_0_g\
        );

    \I__7796\ : InMux
    port map (
            O => \N__34225\,
            I => \N__34222\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__34222\,
            I => \N__34211\
        );

    \I__7794\ : SRMux
    port map (
            O => \N__34221\,
            I => \N__34192\
        );

    \I__7793\ : SRMux
    port map (
            O => \N__34220\,
            I => \N__34192\
        );

    \I__7792\ : SRMux
    port map (
            O => \N__34219\,
            I => \N__34192\
        );

    \I__7791\ : SRMux
    port map (
            O => \N__34218\,
            I => \N__34192\
        );

    \I__7790\ : SRMux
    port map (
            O => \N__34217\,
            I => \N__34192\
        );

    \I__7789\ : SRMux
    port map (
            O => \N__34216\,
            I => \N__34192\
        );

    \I__7788\ : SRMux
    port map (
            O => \N__34215\,
            I => \N__34192\
        );

    \I__7787\ : SRMux
    port map (
            O => \N__34214\,
            I => \N__34192\
        );

    \I__7786\ : Glb2LocalMux
    port map (
            O => \N__34211\,
            I => \N__34192\
        );

    \I__7785\ : GlobalMux
    port map (
            O => \N__34192\,
            I => \N__34189\
        );

    \I__7784\ : gio2CtrlBuf
    port map (
            O => \N__34189\,
            I => \this_vga_signals.N_1637_g\
        );

    \I__7783\ : InMux
    port map (
            O => \N__34186\,
            I => \N__34183\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__34183\,
            I => \N__34180\
        );

    \I__7781\ : Odrv4
    port map (
            O => \N__34180\,
            I => \this_vga_signals.N_5_i_0\
        );

    \I__7780\ : CascadeMux
    port map (
            O => \N__34177\,
            I => \this_vga_signals.N_5_i_0_cascade_\
        );

    \I__7779\ : InMux
    port map (
            O => \N__34174\,
            I => \N__34171\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__34171\,
            I => \N__34168\
        );

    \I__7777\ : Span4Mux_v
    port map (
            O => \N__34168\,
            I => \N__34165\
        );

    \I__7776\ : Odrv4
    port map (
            O => \N__34165\,
            I => \this_vga_signals.mult1_un47_sum_0_1\
        );

    \I__7775\ : InMux
    port map (
            O => \N__34162\,
            I => \N__34159\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__34159\,
            I => \N__34156\
        );

    \I__7773\ : Odrv12
    port map (
            O => \N__34156\,
            I => \this_vga_signals.g0_21_1\
        );

    \I__7772\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34149\
        );

    \I__7771\ : InMux
    port map (
            O => \N__34152\,
            I => \N__34146\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__34149\,
            I => \this_vga_signals.mult1_un47_sum_axb1\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__34146\,
            I => \this_vga_signals.mult1_un47_sum_axb1\
        );

    \I__7768\ : InMux
    port map (
            O => \N__34141\,
            I => \N__34138\
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__34138\,
            I => \N__34133\
        );

    \I__7766\ : CascadeMux
    port map (
            O => \N__34137\,
            I => \N__34127\
        );

    \I__7765\ : CascadeMux
    port map (
            O => \N__34136\,
            I => \N__34120\
        );

    \I__7764\ : Span4Mux_h
    port map (
            O => \N__34133\,
            I => \N__34115\
        );

    \I__7763\ : InMux
    port map (
            O => \N__34132\,
            I => \N__34110\
        );

    \I__7762\ : InMux
    port map (
            O => \N__34131\,
            I => \N__34110\
        );

    \I__7761\ : InMux
    port map (
            O => \N__34130\,
            I => \N__34101\
        );

    \I__7760\ : InMux
    port map (
            O => \N__34127\,
            I => \N__34101\
        );

    \I__7759\ : InMux
    port map (
            O => \N__34126\,
            I => \N__34101\
        );

    \I__7758\ : InMux
    port map (
            O => \N__34125\,
            I => \N__34101\
        );

    \I__7757\ : InMux
    port map (
            O => \N__34124\,
            I => \N__34098\
        );

    \I__7756\ : InMux
    port map (
            O => \N__34123\,
            I => \N__34095\
        );

    \I__7755\ : InMux
    port map (
            O => \N__34120\,
            I => \N__34088\
        );

    \I__7754\ : InMux
    port map (
            O => \N__34119\,
            I => \N__34088\
        );

    \I__7753\ : InMux
    port map (
            O => \N__34118\,
            I => \N__34088\
        );

    \I__7752\ : Odrv4
    port map (
            O => \N__34115\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__34110\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__34101\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__34098\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__34095\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__34088\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__7746\ : InMux
    port map (
            O => \N__34075\,
            I => \N__34061\
        );

    \I__7745\ : InMux
    port map (
            O => \N__34074\,
            I => \N__34061\
        );

    \I__7744\ : InMux
    port map (
            O => \N__34073\,
            I => \N__34061\
        );

    \I__7743\ : InMux
    port map (
            O => \N__34072\,
            I => \N__34058\
        );

    \I__7742\ : InMux
    port map (
            O => \N__34071\,
            I => \N__34053\
        );

    \I__7741\ : InMux
    port map (
            O => \N__34070\,
            I => \N__34053\
        );

    \I__7740\ : InMux
    port map (
            O => \N__34069\,
            I => \N__34048\
        );

    \I__7739\ : InMux
    port map (
            O => \N__34068\,
            I => \N__34048\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__34061\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_3\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__34058\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_3\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__34053\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_3\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__34048\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_3\
        );

    \I__7734\ : InMux
    port map (
            O => \N__34039\,
            I => \N__34036\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__34036\,
            I => \N__34033\
        );

    \I__7732\ : Span4Mux_h
    port map (
            O => \N__34033\,
            I => \N__34030\
        );

    \I__7731\ : Odrv4
    port map (
            O => \N__34030\,
            I => \this_vga_signals.mult1_un47_sum_1_1\
        );

    \I__7730\ : InMux
    port map (
            O => \N__34027\,
            I => \N__34024\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__34024\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_6\
        );

    \I__7728\ : InMux
    port map (
            O => \N__34021\,
            I => \N__34018\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__34018\,
            I => \N__34015\
        );

    \I__7726\ : Span4Mux_h
    port map (
            O => \N__34015\,
            I => \N__34012\
        );

    \I__7725\ : Span4Mux_v
    port map (
            O => \N__34012\,
            I => \N__34009\
        );

    \I__7724\ : Odrv4
    port map (
            O => \N__34009\,
            I => \this_spr_ram.mem_out_bus4_2\
        );

    \I__7723\ : InMux
    port map (
            O => \N__34006\,
            I => \N__34003\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__34003\,
            I => \N__34000\
        );

    \I__7721\ : Span4Mux_h
    port map (
            O => \N__34000\,
            I => \N__33997\
        );

    \I__7720\ : Span4Mux_v
    port map (
            O => \N__33997\,
            I => \N__33994\
        );

    \I__7719\ : Span4Mux_v
    port map (
            O => \N__33994\,
            I => \N__33991\
        );

    \I__7718\ : Odrv4
    port map (
            O => \N__33991\,
            I => \this_spr_ram.mem_out_bus0_2\
        );

    \I__7717\ : CascadeMux
    port map (
            O => \N__33988\,
            I => \this_spr_ram.mem_mem_0_1_RNIM6VFZ0_cascade_\
        );

    \I__7716\ : CascadeMux
    port map (
            O => \N__33985\,
            I => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\
        );

    \I__7715\ : CascadeMux
    port map (
            O => \N__33982\,
            I => \M_this_spr_ram_read_data_2_cascade_\
        );

    \I__7714\ : InMux
    port map (
            O => \N__33979\,
            I => \N__33976\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__33976\,
            I => \N__33973\
        );

    \I__7712\ : Span12Mux_s9_h
    port map (
            O => \N__33973\,
            I => \N__33970\
        );

    \I__7711\ : Span12Mux_h
    port map (
            O => \N__33970\,
            I => \N__33967\
        );

    \I__7710\ : Odrv12
    port map (
            O => \N__33967\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__7709\ : InMux
    port map (
            O => \N__33964\,
            I => \N__33961\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__33961\,
            I => \N__33958\
        );

    \I__7707\ : Span4Mux_v
    port map (
            O => \N__33958\,
            I => \N__33955\
        );

    \I__7706\ : Span4Mux_h
    port map (
            O => \N__33955\,
            I => \N__33952\
        );

    \I__7705\ : Odrv4
    port map (
            O => \N__33952\,
            I => \this_spr_ram.mem_out_bus5_0\
        );

    \I__7704\ : InMux
    port map (
            O => \N__33949\,
            I => \N__33946\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__33946\,
            I => \N__33943\
        );

    \I__7702\ : Span4Mux_v
    port map (
            O => \N__33943\,
            I => \N__33940\
        );

    \I__7701\ : Span4Mux_h
    port map (
            O => \N__33940\,
            I => \N__33937\
        );

    \I__7700\ : Span4Mux_v
    port map (
            O => \N__33937\,
            I => \N__33934\
        );

    \I__7699\ : Odrv4
    port map (
            O => \N__33934\,
            I => \this_spr_ram.mem_out_bus1_0\
        );

    \I__7698\ : InMux
    port map (
            O => \N__33931\,
            I => \N__33928\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__33928\,
            I => \N__33925\
        );

    \I__7696\ : Span4Mux_h
    port map (
            O => \N__33925\,
            I => \N__33922\
        );

    \I__7695\ : Odrv4
    port map (
            O => \N__33922\,
            I => \this_spr_ram.mem_out_bus4_1\
        );

    \I__7694\ : InMux
    port map (
            O => \N__33919\,
            I => \N__33916\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__33916\,
            I => \N__33913\
        );

    \I__7692\ : Span4Mux_h
    port map (
            O => \N__33913\,
            I => \N__33910\
        );

    \I__7691\ : Span4Mux_v
    port map (
            O => \N__33910\,
            I => \N__33907\
        );

    \I__7690\ : Span4Mux_v
    port map (
            O => \N__33907\,
            I => \N__33904\
        );

    \I__7689\ : Span4Mux_v
    port map (
            O => \N__33904\,
            I => \N__33901\
        );

    \I__7688\ : Odrv4
    port map (
            O => \N__33901\,
            I => \this_spr_ram.mem_out_bus0_1\
        );

    \I__7687\ : CascadeMux
    port map (
            O => \N__33898\,
            I => \this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0_cascade_\
        );

    \I__7686\ : CascadeMux
    port map (
            O => \N__33895\,
            I => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\
        );

    \I__7685\ : CascadeMux
    port map (
            O => \N__33892\,
            I => \N__33887\
        );

    \I__7684\ : CascadeMux
    port map (
            O => \N__33891\,
            I => \N__33882\
        );

    \I__7683\ : CascadeMux
    port map (
            O => \N__33890\,
            I => \N__33877\
        );

    \I__7682\ : InMux
    port map (
            O => \N__33887\,
            I => \N__33873\
        );

    \I__7681\ : CascadeMux
    port map (
            O => \N__33886\,
            I => \N__33870\
        );

    \I__7680\ : CascadeMux
    port map (
            O => \N__33885\,
            I => \N__33867\
        );

    \I__7679\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33864\
        );

    \I__7678\ : CascadeMux
    port map (
            O => \N__33881\,
            I => \N__33861\
        );

    \I__7677\ : CascadeMux
    port map (
            O => \N__33880\,
            I => \N__33857\
        );

    \I__7676\ : InMux
    port map (
            O => \N__33877\,
            I => \N__33853\
        );

    \I__7675\ : CascadeMux
    port map (
            O => \N__33876\,
            I => \N__33850\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__33873\,
            I => \N__33846\
        );

    \I__7673\ : InMux
    port map (
            O => \N__33870\,
            I => \N__33843\
        );

    \I__7672\ : InMux
    port map (
            O => \N__33867\,
            I => \N__33840\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__33864\,
            I => \N__33837\
        );

    \I__7670\ : InMux
    port map (
            O => \N__33861\,
            I => \N__33834\
        );

    \I__7669\ : CascadeMux
    port map (
            O => \N__33860\,
            I => \N__33831\
        );

    \I__7668\ : InMux
    port map (
            O => \N__33857\,
            I => \N__33827\
        );

    \I__7667\ : CascadeMux
    port map (
            O => \N__33856\,
            I => \N__33824\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__33853\,
            I => \N__33821\
        );

    \I__7665\ : InMux
    port map (
            O => \N__33850\,
            I => \N__33818\
        );

    \I__7664\ : CascadeMux
    port map (
            O => \N__33849\,
            I => \N__33815\
        );

    \I__7663\ : Span4Mux_s1_v
    port map (
            O => \N__33846\,
            I => \N__33806\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__33843\,
            I => \N__33806\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__33840\,
            I => \N__33806\
        );

    \I__7660\ : Span4Mux_h
    port map (
            O => \N__33837\,
            I => \N__33801\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__33834\,
            I => \N__33801\
        );

    \I__7658\ : InMux
    port map (
            O => \N__33831\,
            I => \N__33798\
        );

    \I__7657\ : CascadeMux
    port map (
            O => \N__33830\,
            I => \N__33795\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__33827\,
            I => \N__33791\
        );

    \I__7655\ : InMux
    port map (
            O => \N__33824\,
            I => \N__33788\
        );

    \I__7654\ : Span4Mux_v
    port map (
            O => \N__33821\,
            I => \N__33783\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__33818\,
            I => \N__33783\
        );

    \I__7652\ : InMux
    port map (
            O => \N__33815\,
            I => \N__33780\
        );

    \I__7651\ : CascadeMux
    port map (
            O => \N__33814\,
            I => \N__33777\
        );

    \I__7650\ : CascadeMux
    port map (
            O => \N__33813\,
            I => \N__33774\
        );

    \I__7649\ : Span4Mux_v
    port map (
            O => \N__33806\,
            I => \N__33770\
        );

    \I__7648\ : Span4Mux_v
    port map (
            O => \N__33801\,
            I => \N__33765\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__33798\,
            I => \N__33765\
        );

    \I__7646\ : InMux
    port map (
            O => \N__33795\,
            I => \N__33762\
        );

    \I__7645\ : CascadeMux
    port map (
            O => \N__33794\,
            I => \N__33759\
        );

    \I__7644\ : Span4Mux_v
    port map (
            O => \N__33791\,
            I => \N__33754\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__33788\,
            I => \N__33754\
        );

    \I__7642\ : Span4Mux_v
    port map (
            O => \N__33783\,
            I => \N__33749\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__33780\,
            I => \N__33749\
        );

    \I__7640\ : InMux
    port map (
            O => \N__33777\,
            I => \N__33746\
        );

    \I__7639\ : InMux
    port map (
            O => \N__33774\,
            I => \N__33743\
        );

    \I__7638\ : CascadeMux
    port map (
            O => \N__33773\,
            I => \N__33740\
        );

    \I__7637\ : Sp12to4
    port map (
            O => \N__33770\,
            I => \N__33737\
        );

    \I__7636\ : Span4Mux_h
    port map (
            O => \N__33765\,
            I => \N__33732\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__33762\,
            I => \N__33732\
        );

    \I__7634\ : InMux
    port map (
            O => \N__33759\,
            I => \N__33729\
        );

    \I__7633\ : Span4Mux_v
    port map (
            O => \N__33754\,
            I => \N__33722\
        );

    \I__7632\ : Span4Mux_h
    port map (
            O => \N__33749\,
            I => \N__33722\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__33746\,
            I => \N__33722\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__33743\,
            I => \N__33719\
        );

    \I__7629\ : InMux
    port map (
            O => \N__33740\,
            I => \N__33716\
        );

    \I__7628\ : Span12Mux_h
    port map (
            O => \N__33737\,
            I => \N__33713\
        );

    \I__7627\ : Span4Mux_v
    port map (
            O => \N__33732\,
            I => \N__33708\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__33729\,
            I => \N__33708\
        );

    \I__7625\ : Span4Mux_v
    port map (
            O => \N__33722\,
            I => \N__33701\
        );

    \I__7624\ : Span4Mux_v
    port map (
            O => \N__33719\,
            I => \N__33701\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__33716\,
            I => \N__33701\
        );

    \I__7622\ : Span12Mux_v
    port map (
            O => \N__33713\,
            I => \N__33697\
        );

    \I__7621\ : Span4Mux_h
    port map (
            O => \N__33708\,
            I => \N__33692\
        );

    \I__7620\ : Span4Mux_h
    port map (
            O => \N__33701\,
            I => \N__33692\
        );

    \I__7619\ : InMux
    port map (
            O => \N__33700\,
            I => \N__33689\
        );

    \I__7618\ : Odrv12
    port map (
            O => \N__33697\,
            I => \M_this_spr_address_qZ0Z_8\
        );

    \I__7617\ : Odrv4
    port map (
            O => \N__33692\,
            I => \M_this_spr_address_qZ0Z_8\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__33689\,
            I => \M_this_spr_address_qZ0Z_8\
        );

    \I__7615\ : InMux
    port map (
            O => \N__33682\,
            I => \bfn_22_15_0_\
        );

    \I__7614\ : CascadeMux
    port map (
            O => \N__33679\,
            I => \N__33675\
        );

    \I__7613\ : CascadeMux
    port map (
            O => \N__33678\,
            I => \N__33670\
        );

    \I__7612\ : InMux
    port map (
            O => \N__33675\,
            I => \N__33666\
        );

    \I__7611\ : CascadeMux
    port map (
            O => \N__33674\,
            I => \N__33663\
        );

    \I__7610\ : CascadeMux
    port map (
            O => \N__33673\,
            I => \N__33659\
        );

    \I__7609\ : InMux
    port map (
            O => \N__33670\,
            I => \N__33655\
        );

    \I__7608\ : CascadeMux
    port map (
            O => \N__33669\,
            I => \N__33652\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__33666\,
            I => \N__33646\
        );

    \I__7606\ : InMux
    port map (
            O => \N__33663\,
            I => \N__33643\
        );

    \I__7605\ : CascadeMux
    port map (
            O => \N__33662\,
            I => \N__33640\
        );

    \I__7604\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33637\
        );

    \I__7603\ : CascadeMux
    port map (
            O => \N__33658\,
            I => \N__33634\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__33655\,
            I => \N__33630\
        );

    \I__7601\ : InMux
    port map (
            O => \N__33652\,
            I => \N__33627\
        );

    \I__7600\ : CascadeMux
    port map (
            O => \N__33651\,
            I => \N__33624\
        );

    \I__7599\ : CascadeMux
    port map (
            O => \N__33650\,
            I => \N__33621\
        );

    \I__7598\ : CascadeMux
    port map (
            O => \N__33649\,
            I => \N__33617\
        );

    \I__7597\ : Span4Mux_s1_v
    port map (
            O => \N__33646\,
            I => \N__33611\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__33643\,
            I => \N__33611\
        );

    \I__7595\ : InMux
    port map (
            O => \N__33640\,
            I => \N__33608\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__33637\,
            I => \N__33604\
        );

    \I__7593\ : InMux
    port map (
            O => \N__33634\,
            I => \N__33601\
        );

    \I__7592\ : CascadeMux
    port map (
            O => \N__33633\,
            I => \N__33598\
        );

    \I__7591\ : Span4Mux_h
    port map (
            O => \N__33630\,
            I => \N__33592\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__33627\,
            I => \N__33592\
        );

    \I__7589\ : InMux
    port map (
            O => \N__33624\,
            I => \N__33589\
        );

    \I__7588\ : InMux
    port map (
            O => \N__33621\,
            I => \N__33586\
        );

    \I__7587\ : CascadeMux
    port map (
            O => \N__33620\,
            I => \N__33583\
        );

    \I__7586\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33580\
        );

    \I__7585\ : CascadeMux
    port map (
            O => \N__33616\,
            I => \N__33577\
        );

    \I__7584\ : Span4Mux_v
    port map (
            O => \N__33611\,
            I => \N__33573\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__33608\,
            I => \N__33570\
        );

    \I__7582\ : CascadeMux
    port map (
            O => \N__33607\,
            I => \N__33567\
        );

    \I__7581\ : Span4Mux_v
    port map (
            O => \N__33604\,
            I => \N__33562\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__33601\,
            I => \N__33562\
        );

    \I__7579\ : InMux
    port map (
            O => \N__33598\,
            I => \N__33559\
        );

    \I__7578\ : CascadeMux
    port map (
            O => \N__33597\,
            I => \N__33556\
        );

    \I__7577\ : Span4Mux_v
    port map (
            O => \N__33592\,
            I => \N__33549\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__33589\,
            I => \N__33549\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__33586\,
            I => \N__33549\
        );

    \I__7574\ : InMux
    port map (
            O => \N__33583\,
            I => \N__33546\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__33580\,
            I => \N__33543\
        );

    \I__7572\ : InMux
    port map (
            O => \N__33577\,
            I => \N__33540\
        );

    \I__7571\ : CascadeMux
    port map (
            O => \N__33576\,
            I => \N__33537\
        );

    \I__7570\ : Sp12to4
    port map (
            O => \N__33573\,
            I => \N__33534\
        );

    \I__7569\ : Span12Mux_s9_h
    port map (
            O => \N__33570\,
            I => \N__33531\
        );

    \I__7568\ : InMux
    port map (
            O => \N__33567\,
            I => \N__33528\
        );

    \I__7567\ : Span4Mux_h
    port map (
            O => \N__33562\,
            I => \N__33523\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__33559\,
            I => \N__33523\
        );

    \I__7565\ : InMux
    port map (
            O => \N__33556\,
            I => \N__33520\
        );

    \I__7564\ : Span4Mux_v
    port map (
            O => \N__33549\,
            I => \N__33517\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__33546\,
            I => \N__33514\
        );

    \I__7562\ : Span4Mux_v
    port map (
            O => \N__33543\,
            I => \N__33509\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__33540\,
            I => \N__33509\
        );

    \I__7560\ : InMux
    port map (
            O => \N__33537\,
            I => \N__33506\
        );

    \I__7559\ : Span12Mux_h
    port map (
            O => \N__33534\,
            I => \N__33503\
        );

    \I__7558\ : Span12Mux_h
    port map (
            O => \N__33531\,
            I => \N__33500\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__33528\,
            I => \N__33497\
        );

    \I__7556\ : Span4Mux_v
    port map (
            O => \N__33523\,
            I => \N__33492\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__33520\,
            I => \N__33492\
        );

    \I__7554\ : Span4Mux_v
    port map (
            O => \N__33517\,
            I => \N__33483\
        );

    \I__7553\ : Span4Mux_v
    port map (
            O => \N__33514\,
            I => \N__33483\
        );

    \I__7552\ : Span4Mux_v
    port map (
            O => \N__33509\,
            I => \N__33483\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__33506\,
            I => \N__33483\
        );

    \I__7550\ : Span12Mux_v
    port map (
            O => \N__33503\,
            I => \N__33479\
        );

    \I__7549\ : Span12Mux_v
    port map (
            O => \N__33500\,
            I => \N__33474\
        );

    \I__7548\ : Span12Mux_s10_h
    port map (
            O => \N__33497\,
            I => \N__33474\
        );

    \I__7547\ : Span4Mux_h
    port map (
            O => \N__33492\,
            I => \N__33469\
        );

    \I__7546\ : Span4Mux_h
    port map (
            O => \N__33483\,
            I => \N__33469\
        );

    \I__7545\ : InMux
    port map (
            O => \N__33482\,
            I => \N__33466\
        );

    \I__7544\ : Odrv12
    port map (
            O => \N__33479\,
            I => \M_this_spr_address_qZ0Z_9\
        );

    \I__7543\ : Odrv12
    port map (
            O => \N__33474\,
            I => \M_this_spr_address_qZ0Z_9\
        );

    \I__7542\ : Odrv4
    port map (
            O => \N__33469\,
            I => \M_this_spr_address_qZ0Z_9\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__33466\,
            I => \M_this_spr_address_qZ0Z_9\
        );

    \I__7540\ : InMux
    port map (
            O => \N__33457\,
            I => \un1_M_this_spr_address_q_cry_8\
        );

    \I__7539\ : CascadeMux
    port map (
            O => \N__33454\,
            I => \N__33449\
        );

    \I__7538\ : CascadeMux
    port map (
            O => \N__33453\,
            I => \N__33445\
        );

    \I__7537\ : CascadeMux
    port map (
            O => \N__33452\,
            I => \N__33440\
        );

    \I__7536\ : InMux
    port map (
            O => \N__33449\,
            I => \N__33437\
        );

    \I__7535\ : CascadeMux
    port map (
            O => \N__33448\,
            I => \N__33434\
        );

    \I__7534\ : InMux
    port map (
            O => \N__33445\,
            I => \N__33427\
        );

    \I__7533\ : CascadeMux
    port map (
            O => \N__33444\,
            I => \N__33424\
        );

    \I__7532\ : CascadeMux
    port map (
            O => \N__33443\,
            I => \N__33420\
        );

    \I__7531\ : InMux
    port map (
            O => \N__33440\,
            I => \N__33416\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__33437\,
            I => \N__33413\
        );

    \I__7529\ : InMux
    port map (
            O => \N__33434\,
            I => \N__33410\
        );

    \I__7528\ : CascadeMux
    port map (
            O => \N__33433\,
            I => \N__33407\
        );

    \I__7527\ : CascadeMux
    port map (
            O => \N__33432\,
            I => \N__33404\
        );

    \I__7526\ : CascadeMux
    port map (
            O => \N__33431\,
            I => \N__33399\
        );

    \I__7525\ : CascadeMux
    port map (
            O => \N__33430\,
            I => \N__33396\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__33427\,
            I => \N__33393\
        );

    \I__7523\ : InMux
    port map (
            O => \N__33424\,
            I => \N__33390\
        );

    \I__7522\ : CascadeMux
    port map (
            O => \N__33423\,
            I => \N__33387\
        );

    \I__7521\ : InMux
    port map (
            O => \N__33420\,
            I => \N__33383\
        );

    \I__7520\ : CascadeMux
    port map (
            O => \N__33419\,
            I => \N__33380\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__33416\,
            I => \N__33373\
        );

    \I__7518\ : Span4Mux_s1_v
    port map (
            O => \N__33413\,
            I => \N__33373\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__33410\,
            I => \N__33373\
        );

    \I__7516\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33369\
        );

    \I__7515\ : InMux
    port map (
            O => \N__33404\,
            I => \N__33366\
        );

    \I__7514\ : CascadeMux
    port map (
            O => \N__33403\,
            I => \N__33363\
        );

    \I__7513\ : CascadeMux
    port map (
            O => \N__33402\,
            I => \N__33360\
        );

    \I__7512\ : InMux
    port map (
            O => \N__33399\,
            I => \N__33357\
        );

    \I__7511\ : InMux
    port map (
            O => \N__33396\,
            I => \N__33354\
        );

    \I__7510\ : Span4Mux_v
    port map (
            O => \N__33393\,
            I => \N__33349\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__33390\,
            I => \N__33349\
        );

    \I__7508\ : InMux
    port map (
            O => \N__33387\,
            I => \N__33346\
        );

    \I__7507\ : CascadeMux
    port map (
            O => \N__33386\,
            I => \N__33343\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__33383\,
            I => \N__33340\
        );

    \I__7505\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33337\
        );

    \I__7504\ : Span4Mux_v
    port map (
            O => \N__33373\,
            I => \N__33334\
        );

    \I__7503\ : CascadeMux
    port map (
            O => \N__33372\,
            I => \N__33331\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__33369\,
            I => \N__33328\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__33366\,
            I => \N__33325\
        );

    \I__7500\ : InMux
    port map (
            O => \N__33363\,
            I => \N__33322\
        );

    \I__7499\ : InMux
    port map (
            O => \N__33360\,
            I => \N__33319\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__33357\,
            I => \N__33316\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__33354\,
            I => \N__33313\
        );

    \I__7496\ : Span4Mux_h
    port map (
            O => \N__33349\,
            I => \N__33310\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__33346\,
            I => \N__33307\
        );

    \I__7494\ : InMux
    port map (
            O => \N__33343\,
            I => \N__33304\
        );

    \I__7493\ : Span4Mux_v
    port map (
            O => \N__33340\,
            I => \N__33299\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__33337\,
            I => \N__33299\
        );

    \I__7491\ : Span4Mux_h
    port map (
            O => \N__33334\,
            I => \N__33296\
        );

    \I__7490\ : InMux
    port map (
            O => \N__33331\,
            I => \N__33293\
        );

    \I__7489\ : Span4Mux_v
    port map (
            O => \N__33328\,
            I => \N__33286\
        );

    \I__7488\ : Span4Mux_v
    port map (
            O => \N__33325\,
            I => \N__33286\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__33322\,
            I => \N__33286\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__33319\,
            I => \N__33281\
        );

    \I__7485\ : Span4Mux_v
    port map (
            O => \N__33316\,
            I => \N__33281\
        );

    \I__7484\ : Span4Mux_h
    port map (
            O => \N__33313\,
            I => \N__33276\
        );

    \I__7483\ : Span4Mux_v
    port map (
            O => \N__33310\,
            I => \N__33276\
        );

    \I__7482\ : Span4Mux_v
    port map (
            O => \N__33307\,
            I => \N__33271\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__33304\,
            I => \N__33271\
        );

    \I__7480\ : Span4Mux_h
    port map (
            O => \N__33299\,
            I => \N__33268\
        );

    \I__7479\ : Sp12to4
    port map (
            O => \N__33296\,
            I => \N__33265\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__33293\,
            I => \N__33261\
        );

    \I__7477\ : Span4Mux_h
    port map (
            O => \N__33286\,
            I => \N__33254\
        );

    \I__7476\ : Span4Mux_h
    port map (
            O => \N__33281\,
            I => \N__33254\
        );

    \I__7475\ : Span4Mux_v
    port map (
            O => \N__33276\,
            I => \N__33254\
        );

    \I__7474\ : Span4Mux_h
    port map (
            O => \N__33271\,
            I => \N__33249\
        );

    \I__7473\ : Span4Mux_v
    port map (
            O => \N__33268\,
            I => \N__33249\
        );

    \I__7472\ : Span12Mux_v
    port map (
            O => \N__33265\,
            I => \N__33246\
        );

    \I__7471\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33243\
        );

    \I__7470\ : Span4Mux_h
    port map (
            O => \N__33261\,
            I => \N__33236\
        );

    \I__7469\ : Span4Mux_v
    port map (
            O => \N__33254\,
            I => \N__33236\
        );

    \I__7468\ : Span4Mux_v
    port map (
            O => \N__33249\,
            I => \N__33236\
        );

    \I__7467\ : Span12Mux_h
    port map (
            O => \N__33246\,
            I => \N__33233\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__33243\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__7465\ : Odrv4
    port map (
            O => \N__33236\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__7464\ : Odrv12
    port map (
            O => \N__33233\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__7463\ : InMux
    port map (
            O => \N__33226\,
            I => \un1_M_this_spr_address_q_cry_9\
        );

    \I__7462\ : InMux
    port map (
            O => \N__33223\,
            I => \un1_M_this_spr_address_q_cry_10\
        );

    \I__7461\ : InMux
    port map (
            O => \N__33220\,
            I => \un1_M_this_spr_address_q_cry_11\
        );

    \I__7460\ : InMux
    port map (
            O => \N__33217\,
            I => \N__33195\
        );

    \I__7459\ : InMux
    port map (
            O => \N__33216\,
            I => \N__33195\
        );

    \I__7458\ : InMux
    port map (
            O => \N__33215\,
            I => \N__33195\
        );

    \I__7457\ : InMux
    port map (
            O => \N__33214\,
            I => \N__33195\
        );

    \I__7456\ : InMux
    port map (
            O => \N__33213\,
            I => \N__33186\
        );

    \I__7455\ : InMux
    port map (
            O => \N__33212\,
            I => \N__33186\
        );

    \I__7454\ : InMux
    port map (
            O => \N__33211\,
            I => \N__33186\
        );

    \I__7453\ : InMux
    port map (
            O => \N__33210\,
            I => \N__33186\
        );

    \I__7452\ : InMux
    port map (
            O => \N__33209\,
            I => \N__33181\
        );

    \I__7451\ : InMux
    port map (
            O => \N__33208\,
            I => \N__33181\
        );

    \I__7450\ : InMux
    port map (
            O => \N__33207\,
            I => \N__33172\
        );

    \I__7449\ : InMux
    port map (
            O => \N__33206\,
            I => \N__33172\
        );

    \I__7448\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33172\
        );

    \I__7447\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33172\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__33195\,
            I => \N__33165\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__33186\,
            I => \N__33165\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__33181\,
            I => \N__33160\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__33172\,
            I => \N__33160\
        );

    \I__7442\ : CascadeMux
    port map (
            O => \N__33171\,
            I => \N__33157\
        );

    \I__7441\ : CascadeMux
    port map (
            O => \N__33170\,
            I => \N__33154\
        );

    \I__7440\ : Span4Mux_v
    port map (
            O => \N__33165\,
            I => \N__33151\
        );

    \I__7439\ : Span4Mux_h
    port map (
            O => \N__33160\,
            I => \N__33148\
        );

    \I__7438\ : InMux
    port map (
            O => \N__33157\,
            I => \N__33145\
        );

    \I__7437\ : InMux
    port map (
            O => \N__33154\,
            I => \N__33142\
        );

    \I__7436\ : Sp12to4
    port map (
            O => \N__33151\,
            I => \N__33139\
        );

    \I__7435\ : Span4Mux_v
    port map (
            O => \N__33148\,
            I => \N__33136\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__33145\,
            I => \N__33133\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__33142\,
            I => \N__33128\
        );

    \I__7432\ : Span12Mux_h
    port map (
            O => \N__33139\,
            I => \N__33128\
        );

    \I__7431\ : Span4Mux_h
    port map (
            O => \N__33136\,
            I => \N__33125\
        );

    \I__7430\ : Odrv12
    port map (
            O => \N__33133\,
            I => \N_1005_0\
        );

    \I__7429\ : Odrv12
    port map (
            O => \N__33128\,
            I => \N_1005_0\
        );

    \I__7428\ : Odrv4
    port map (
            O => \N__33125\,
            I => \N_1005_0\
        );

    \I__7427\ : InMux
    port map (
            O => \N__33118\,
            I => \un1_M_this_spr_address_q_cry_12\
        );

    \I__7426\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33112\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__33112\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_5\
        );

    \I__7424\ : InMux
    port map (
            O => \N__33109\,
            I => \N__33106\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__33106\,
            I => \N__33103\
        );

    \I__7422\ : Span4Mux_v
    port map (
            O => \N__33103\,
            I => \N__33100\
        );

    \I__7421\ : Sp12to4
    port map (
            O => \N__33100\,
            I => \N__33097\
        );

    \I__7420\ : Span12Mux_h
    port map (
            O => \N__33097\,
            I => \N__33094\
        );

    \I__7419\ : Odrv12
    port map (
            O => \N__33094\,
            I => \this_ppu.oam_cache.mem_6\
        );

    \I__7418\ : InMux
    port map (
            O => \N__33091\,
            I => \N__33084\
        );

    \I__7417\ : InMux
    port map (
            O => \N__33090\,
            I => \N__33081\
        );

    \I__7416\ : InMux
    port map (
            O => \N__33089\,
            I => \N__33076\
        );

    \I__7415\ : InMux
    port map (
            O => \N__33088\,
            I => \N__33076\
        );

    \I__7414\ : CascadeMux
    port map (
            O => \N__33087\,
            I => \N__33070\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__33084\,
            I => \N__33063\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__33081\,
            I => \N__33063\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__33076\,
            I => \N__33063\
        );

    \I__7410\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33056\
        );

    \I__7409\ : InMux
    port map (
            O => \N__33074\,
            I => \N__33056\
        );

    \I__7408\ : InMux
    port map (
            O => \N__33073\,
            I => \N__33056\
        );

    \I__7407\ : InMux
    port map (
            O => \N__33070\,
            I => \N__33053\
        );

    \I__7406\ : Span4Mux_v
    port map (
            O => \N__33063\,
            I => \N__33048\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__33056\,
            I => \N__33043\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__33053\,
            I => \N__33043\
        );

    \I__7403\ : InMux
    port map (
            O => \N__33052\,
            I => \N__33038\
        );

    \I__7402\ : InMux
    port map (
            O => \N__33051\,
            I => \N__33038\
        );

    \I__7401\ : Span4Mux_h
    port map (
            O => \N__33048\,
            I => \N__33031\
        );

    \I__7400\ : Span4Mux_v
    port map (
            O => \N__33043\,
            I => \N__33031\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__33038\,
            I => \N__33031\
        );

    \I__7398\ : Span4Mux_h
    port map (
            O => \N__33031\,
            I => \N__33028\
        );

    \I__7397\ : Span4Mux_h
    port map (
            O => \N__33028\,
            I => \N__33025\
        );

    \I__7396\ : Odrv4
    port map (
            O => \N__33025\,
            I => port_address_in_4
        );

    \I__7395\ : CascadeMux
    port map (
            O => \N__33022\,
            I => \N__33016\
        );

    \I__7394\ : InMux
    port map (
            O => \N__33021\,
            I => \N__33008\
        );

    \I__7393\ : InMux
    port map (
            O => \N__33020\,
            I => \N__33008\
        );

    \I__7392\ : InMux
    port map (
            O => \N__33019\,
            I => \N__33005\
        );

    \I__7391\ : InMux
    port map (
            O => \N__33016\,
            I => \N__33000\
        );

    \I__7390\ : InMux
    port map (
            O => \N__33015\,
            I => \N__33000\
        );

    \I__7389\ : InMux
    port map (
            O => \N__33014\,
            I => \N__32995\
        );

    \I__7388\ : InMux
    port map (
            O => \N__33013\,
            I => \N__32995\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__33008\,
            I => \N__32990\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__33005\,
            I => \N__32990\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__33000\,
            I => \N__32982\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__32995\,
            I => \N__32982\
        );

    \I__7383\ : Span4Mux_v
    port map (
            O => \N__32990\,
            I => \N__32977\
        );

    \I__7382\ : InMux
    port map (
            O => \N__32989\,
            I => \N__32970\
        );

    \I__7381\ : InMux
    port map (
            O => \N__32988\,
            I => \N__32970\
        );

    \I__7380\ : InMux
    port map (
            O => \N__32987\,
            I => \N__32970\
        );

    \I__7379\ : Span4Mux_v
    port map (
            O => \N__32982\,
            I => \N__32967\
        );

    \I__7378\ : InMux
    port map (
            O => \N__32981\,
            I => \N__32962\
        );

    \I__7377\ : InMux
    port map (
            O => \N__32980\,
            I => \N__32962\
        );

    \I__7376\ : Sp12to4
    port map (
            O => \N__32977\,
            I => \N__32953\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__32970\,
            I => \N__32953\
        );

    \I__7374\ : Sp12to4
    port map (
            O => \N__32967\,
            I => \N__32953\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__32962\,
            I => \N__32953\
        );

    \I__7372\ : Span12Mux_h
    port map (
            O => \N__32953\,
            I => \N__32950\
        );

    \I__7371\ : Odrv12
    port map (
            O => \N__32950\,
            I => port_address_in_0
        );

    \I__7370\ : CascadeMux
    port map (
            O => \N__32947\,
            I => \N__32944\
        );

    \I__7369\ : InMux
    port map (
            O => \N__32944\,
            I => \N__32939\
        );

    \I__7368\ : CascadeMux
    port map (
            O => \N__32943\,
            I => \N__32936\
        );

    \I__7367\ : CascadeMux
    port map (
            O => \N__32942\,
            I => \N__32929\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__32939\,
            I => \N__32924\
        );

    \I__7365\ : InMux
    port map (
            O => \N__32936\,
            I => \N__32921\
        );

    \I__7364\ : InMux
    port map (
            O => \N__32935\,
            I => \N__32916\
        );

    \I__7363\ : InMux
    port map (
            O => \N__32934\,
            I => \N__32916\
        );

    \I__7362\ : InMux
    port map (
            O => \N__32933\,
            I => \N__32913\
        );

    \I__7361\ : InMux
    port map (
            O => \N__32932\,
            I => \N__32908\
        );

    \I__7360\ : InMux
    port map (
            O => \N__32929\,
            I => \N__32908\
        );

    \I__7359\ : InMux
    port map (
            O => \N__32928\,
            I => \N__32903\
        );

    \I__7358\ : InMux
    port map (
            O => \N__32927\,
            I => \N__32903\
        );

    \I__7357\ : Span4Mux_h
    port map (
            O => \N__32924\,
            I => \N__32890\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__32921\,
            I => \N__32890\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__32916\,
            I => \N__32890\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__32913\,
            I => \N__32890\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__32908\,
            I => \N__32890\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__32903\,
            I => \N__32890\
        );

    \I__7351\ : Span4Mux_v
    port map (
            O => \N__32890\,
            I => \N__32887\
        );

    \I__7350\ : Span4Mux_h
    port map (
            O => \N__32887\,
            I => \N__32884\
        );

    \I__7349\ : Span4Mux_v
    port map (
            O => \N__32884\,
            I => \N__32881\
        );

    \I__7348\ : Sp12to4
    port map (
            O => \N__32881\,
            I => \N__32878\
        );

    \I__7347\ : Span12Mux_h
    port map (
            O => \N__32878\,
            I => \N__32874\
        );

    \I__7346\ : InMux
    port map (
            O => \N__32877\,
            I => \N__32871\
        );

    \I__7345\ : Odrv12
    port map (
            O => \N__32874\,
            I => port_rw_in
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__32871\,
            I => port_rw_in
        );

    \I__7343\ : CascadeMux
    port map (
            O => \N__32866\,
            I => \N__32863\
        );

    \I__7342\ : InMux
    port map (
            O => \N__32863\,
            I => \N__32860\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__32860\,
            I => \N__32857\
        );

    \I__7340\ : Span4Mux_h
    port map (
            O => \N__32857\,
            I => \N__32853\
        );

    \I__7339\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32850\
        );

    \I__7338\ : Odrv4
    port map (
            O => \N__32853\,
            I => \N_1422\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__32850\,
            I => \N_1422\
        );

    \I__7336\ : CascadeMux
    port map (
            O => \N__32845\,
            I => \N__32840\
        );

    \I__7335\ : CascadeMux
    port map (
            O => \N__32844\,
            I => \N__32834\
        );

    \I__7334\ : CascadeMux
    port map (
            O => \N__32843\,
            I => \N__32831\
        );

    \I__7333\ : InMux
    port map (
            O => \N__32840\,
            I => \N__32827\
        );

    \I__7332\ : CascadeMux
    port map (
            O => \N__32839\,
            I => \N__32824\
        );

    \I__7331\ : CascadeMux
    port map (
            O => \N__32838\,
            I => \N__32820\
        );

    \I__7330\ : CascadeMux
    port map (
            O => \N__32837\,
            I => \N__32817\
        );

    \I__7329\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32812\
        );

    \I__7328\ : InMux
    port map (
            O => \N__32831\,
            I => \N__32809\
        );

    \I__7327\ : CascadeMux
    port map (
            O => \N__32830\,
            I => \N__32806\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__32827\,
            I => \N__32803\
        );

    \I__7325\ : InMux
    port map (
            O => \N__32824\,
            I => \N__32800\
        );

    \I__7324\ : CascadeMux
    port map (
            O => \N__32823\,
            I => \N__32797\
        );

    \I__7323\ : InMux
    port map (
            O => \N__32820\,
            I => \N__32793\
        );

    \I__7322\ : InMux
    port map (
            O => \N__32817\,
            I => \N__32790\
        );

    \I__7321\ : CascadeMux
    port map (
            O => \N__32816\,
            I => \N__32787\
        );

    \I__7320\ : CascadeMux
    port map (
            O => \N__32815\,
            I => \N__32784\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__32812\,
            I => \N__32779\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__32809\,
            I => \N__32776\
        );

    \I__7317\ : InMux
    port map (
            O => \N__32806\,
            I => \N__32773\
        );

    \I__7316\ : Span4Mux_h
    port map (
            O => \N__32803\,
            I => \N__32768\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__32800\,
            I => \N__32768\
        );

    \I__7314\ : InMux
    port map (
            O => \N__32797\,
            I => \N__32765\
        );

    \I__7313\ : CascadeMux
    port map (
            O => \N__32796\,
            I => \N__32762\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__32793\,
            I => \N__32758\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__32790\,
            I => \N__32755\
        );

    \I__7310\ : InMux
    port map (
            O => \N__32787\,
            I => \N__32752\
        );

    \I__7309\ : InMux
    port map (
            O => \N__32784\,
            I => \N__32749\
        );

    \I__7308\ : CascadeMux
    port map (
            O => \N__32783\,
            I => \N__32746\
        );

    \I__7307\ : CascadeMux
    port map (
            O => \N__32782\,
            I => \N__32743\
        );

    \I__7306\ : Span4Mux_s2_v
    port map (
            O => \N__32779\,
            I => \N__32735\
        );

    \I__7305\ : Span4Mux_h
    port map (
            O => \N__32776\,
            I => \N__32735\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__32773\,
            I => \N__32735\
        );

    \I__7303\ : Span4Mux_v
    port map (
            O => \N__32768\,
            I => \N__32730\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__32765\,
            I => \N__32730\
        );

    \I__7301\ : InMux
    port map (
            O => \N__32762\,
            I => \N__32727\
        );

    \I__7300\ : CascadeMux
    port map (
            O => \N__32761\,
            I => \N__32724\
        );

    \I__7299\ : Span4Mux_v
    port map (
            O => \N__32758\,
            I => \N__32715\
        );

    \I__7298\ : Span4Mux_v
    port map (
            O => \N__32755\,
            I => \N__32715\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__32752\,
            I => \N__32715\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__32749\,
            I => \N__32715\
        );

    \I__7295\ : InMux
    port map (
            O => \N__32746\,
            I => \N__32712\
        );

    \I__7294\ : InMux
    port map (
            O => \N__32743\,
            I => \N__32709\
        );

    \I__7293\ : CascadeMux
    port map (
            O => \N__32742\,
            I => \N__32706\
        );

    \I__7292\ : Span4Mux_v
    port map (
            O => \N__32735\,
            I => \N__32703\
        );

    \I__7291\ : Span4Mux_h
    port map (
            O => \N__32730\,
            I => \N__32697\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__32727\,
            I => \N__32697\
        );

    \I__7289\ : InMux
    port map (
            O => \N__32724\,
            I => \N__32694\
        );

    \I__7288\ : Span4Mux_v
    port map (
            O => \N__32715\,
            I => \N__32687\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__32712\,
            I => \N__32687\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__32709\,
            I => \N__32687\
        );

    \I__7285\ : InMux
    port map (
            O => \N__32706\,
            I => \N__32684\
        );

    \I__7284\ : Sp12to4
    port map (
            O => \N__32703\,
            I => \N__32681\
        );

    \I__7283\ : CascadeMux
    port map (
            O => \N__32702\,
            I => \N__32678\
        );

    \I__7282\ : Span4Mux_v
    port map (
            O => \N__32697\,
            I => \N__32673\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__32694\,
            I => \N__32673\
        );

    \I__7280\ : Span4Mux_v
    port map (
            O => \N__32687\,
            I => \N__32668\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__32684\,
            I => \N__32668\
        );

    \I__7278\ : Span12Mux_h
    port map (
            O => \N__32681\,
            I => \N__32665\
        );

    \I__7277\ : InMux
    port map (
            O => \N__32678\,
            I => \N__32662\
        );

    \I__7276\ : Span4Mux_h
    port map (
            O => \N__32673\,
            I => \N__32656\
        );

    \I__7275\ : Span4Mux_h
    port map (
            O => \N__32668\,
            I => \N__32656\
        );

    \I__7274\ : Span12Mux_v
    port map (
            O => \N__32665\,
            I => \N__32651\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__32662\,
            I => \N__32651\
        );

    \I__7272\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32648\
        );

    \I__7271\ : Odrv4
    port map (
            O => \N__32656\,
            I => \M_this_spr_address_qZ0Z_0\
        );

    \I__7270\ : Odrv12
    port map (
            O => \N__32651\,
            I => \M_this_spr_address_qZ0Z_0\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__32648\,
            I => \M_this_spr_address_qZ0Z_0\
        );

    \I__7268\ : CascadeMux
    port map (
            O => \N__32641\,
            I => \N__32638\
        );

    \I__7267\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32627\
        );

    \I__7266\ : CascadeMux
    port map (
            O => \N__32637\,
            I => \N__32624\
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__32636\,
            I => \N__32620\
        );

    \I__7264\ : CascadeMux
    port map (
            O => \N__32635\,
            I => \N__32617\
        );

    \I__7263\ : CascadeMux
    port map (
            O => \N__32634\,
            I => \N__32614\
        );

    \I__7262\ : CascadeMux
    port map (
            O => \N__32633\,
            I => \N__32610\
        );

    \I__7261\ : CascadeMux
    port map (
            O => \N__32632\,
            I => \N__32606\
        );

    \I__7260\ : CascadeMux
    port map (
            O => \N__32631\,
            I => \N__32603\
        );

    \I__7259\ : CascadeMux
    port map (
            O => \N__32630\,
            I => \N__32598\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__32627\,
            I => \N__32595\
        );

    \I__7257\ : InMux
    port map (
            O => \N__32624\,
            I => \N__32592\
        );

    \I__7256\ : CascadeMux
    port map (
            O => \N__32623\,
            I => \N__32589\
        );

    \I__7255\ : InMux
    port map (
            O => \N__32620\,
            I => \N__32586\
        );

    \I__7254\ : InMux
    port map (
            O => \N__32617\,
            I => \N__32583\
        );

    \I__7253\ : InMux
    port map (
            O => \N__32614\,
            I => \N__32580\
        );

    \I__7252\ : CascadeMux
    port map (
            O => \N__32613\,
            I => \N__32576\
        );

    \I__7251\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32573\
        );

    \I__7250\ : CascadeMux
    port map (
            O => \N__32609\,
            I => \N__32570\
        );

    \I__7249\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32567\
        );

    \I__7248\ : InMux
    port map (
            O => \N__32603\,
            I => \N__32564\
        );

    \I__7247\ : CascadeMux
    port map (
            O => \N__32602\,
            I => \N__32561\
        );

    \I__7246\ : CascadeMux
    port map (
            O => \N__32601\,
            I => \N__32558\
        );

    \I__7245\ : InMux
    port map (
            O => \N__32598\,
            I => \N__32555\
        );

    \I__7244\ : Span4Mux_v
    port map (
            O => \N__32595\,
            I => \N__32550\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__32592\,
            I => \N__32550\
        );

    \I__7242\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32547\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__32586\,
            I => \N__32544\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__32583\,
            I => \N__32541\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__32580\,
            I => \N__32538\
        );

    \I__7238\ : CascadeMux
    port map (
            O => \N__32579\,
            I => \N__32534\
        );

    \I__7237\ : InMux
    port map (
            O => \N__32576\,
            I => \N__32531\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__32573\,
            I => \N__32528\
        );

    \I__7235\ : InMux
    port map (
            O => \N__32570\,
            I => \N__32525\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__32567\,
            I => \N__32520\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__32564\,
            I => \N__32520\
        );

    \I__7232\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32517\
        );

    \I__7231\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32514\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__32555\,
            I => \N__32511\
        );

    \I__7229\ : Span4Mux_h
    port map (
            O => \N__32550\,
            I => \N__32508\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__32547\,
            I => \N__32505\
        );

    \I__7227\ : Span4Mux_h
    port map (
            O => \N__32544\,
            I => \N__32502\
        );

    \I__7226\ : Span4Mux_h
    port map (
            O => \N__32541\,
            I => \N__32499\
        );

    \I__7225\ : Span4Mux_h
    port map (
            O => \N__32538\,
            I => \N__32496\
        );

    \I__7224\ : CascadeMux
    port map (
            O => \N__32537\,
            I => \N__32493\
        );

    \I__7223\ : InMux
    port map (
            O => \N__32534\,
            I => \N__32490\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__32531\,
            I => \N__32487\
        );

    \I__7221\ : Span4Mux_v
    port map (
            O => \N__32528\,
            I => \N__32482\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__32525\,
            I => \N__32482\
        );

    \I__7219\ : Span4Mux_v
    port map (
            O => \N__32520\,
            I => \N__32477\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__32517\,
            I => \N__32477\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__32514\,
            I => \N__32474\
        );

    \I__7216\ : Span4Mux_h
    port map (
            O => \N__32511\,
            I => \N__32471\
        );

    \I__7215\ : Span4Mux_h
    port map (
            O => \N__32508\,
            I => \N__32466\
        );

    \I__7214\ : Span4Mux_h
    port map (
            O => \N__32505\,
            I => \N__32466\
        );

    \I__7213\ : Sp12to4
    port map (
            O => \N__32502\,
            I => \N__32459\
        );

    \I__7212\ : Sp12to4
    port map (
            O => \N__32499\,
            I => \N__32459\
        );

    \I__7211\ : Sp12to4
    port map (
            O => \N__32496\,
            I => \N__32459\
        );

    \I__7210\ : InMux
    port map (
            O => \N__32493\,
            I => \N__32456\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__32490\,
            I => \N__32453\
        );

    \I__7208\ : Span4Mux_h
    port map (
            O => \N__32487\,
            I => \N__32448\
        );

    \I__7207\ : Span4Mux_h
    port map (
            O => \N__32482\,
            I => \N__32448\
        );

    \I__7206\ : Span4Mux_h
    port map (
            O => \N__32477\,
            I => \N__32445\
        );

    \I__7205\ : Span4Mux_h
    port map (
            O => \N__32474\,
            I => \N__32442\
        );

    \I__7204\ : Sp12to4
    port map (
            O => \N__32471\,
            I => \N__32436\
        );

    \I__7203\ : Sp12to4
    port map (
            O => \N__32466\,
            I => \N__32436\
        );

    \I__7202\ : Span12Mux_s9_v
    port map (
            O => \N__32459\,
            I => \N__32433\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__32456\,
            I => \N__32430\
        );

    \I__7200\ : Span4Mux_h
    port map (
            O => \N__32453\,
            I => \N__32425\
        );

    \I__7199\ : Span4Mux_v
    port map (
            O => \N__32448\,
            I => \N__32425\
        );

    \I__7198\ : Span4Mux_v
    port map (
            O => \N__32445\,
            I => \N__32422\
        );

    \I__7197\ : Sp12to4
    port map (
            O => \N__32442\,
            I => \N__32419\
        );

    \I__7196\ : InMux
    port map (
            O => \N__32441\,
            I => \N__32416\
        );

    \I__7195\ : Span12Mux_s9_v
    port map (
            O => \N__32436\,
            I => \N__32411\
        );

    \I__7194\ : Span12Mux_h
    port map (
            O => \N__32433\,
            I => \N__32411\
        );

    \I__7193\ : Odrv4
    port map (
            O => \N__32430\,
            I => \M_this_spr_address_qZ0Z_1\
        );

    \I__7192\ : Odrv4
    port map (
            O => \N__32425\,
            I => \M_this_spr_address_qZ0Z_1\
        );

    \I__7191\ : Odrv4
    port map (
            O => \N__32422\,
            I => \M_this_spr_address_qZ0Z_1\
        );

    \I__7190\ : Odrv12
    port map (
            O => \N__32419\,
            I => \M_this_spr_address_qZ0Z_1\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__32416\,
            I => \M_this_spr_address_qZ0Z_1\
        );

    \I__7188\ : Odrv12
    port map (
            O => \N__32411\,
            I => \M_this_spr_address_qZ0Z_1\
        );

    \I__7187\ : InMux
    port map (
            O => \N__32398\,
            I => \un1_M_this_spr_address_q_cry_0\
        );

    \I__7186\ : CascadeMux
    port map (
            O => \N__32395\,
            I => \N__32392\
        );

    \I__7185\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32387\
        );

    \I__7184\ : CascadeMux
    port map (
            O => \N__32391\,
            I => \N__32384\
        );

    \I__7183\ : CascadeMux
    port map (
            O => \N__32390\,
            I => \N__32381\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__32387\,
            I => \N__32376\
        );

    \I__7181\ : InMux
    port map (
            O => \N__32384\,
            I => \N__32373\
        );

    \I__7180\ : InMux
    port map (
            O => \N__32381\,
            I => \N__32369\
        );

    \I__7179\ : CascadeMux
    port map (
            O => \N__32380\,
            I => \N__32366\
        );

    \I__7178\ : CascadeMux
    port map (
            O => \N__32379\,
            I => \N__32362\
        );

    \I__7177\ : Span4Mux_h
    port map (
            O => \N__32376\,
            I => \N__32355\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__32373\,
            I => \N__32355\
        );

    \I__7175\ : CascadeMux
    port map (
            O => \N__32372\,
            I => \N__32352\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__32369\,
            I => \N__32349\
        );

    \I__7173\ : InMux
    port map (
            O => \N__32366\,
            I => \N__32346\
        );

    \I__7172\ : CascadeMux
    port map (
            O => \N__32365\,
            I => \N__32343\
        );

    \I__7171\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32339\
        );

    \I__7170\ : CascadeMux
    port map (
            O => \N__32361\,
            I => \N__32336\
        );

    \I__7169\ : CascadeMux
    port map (
            O => \N__32360\,
            I => \N__32333\
        );

    \I__7168\ : Span4Mux_v
    port map (
            O => \N__32355\,
            I => \N__32328\
        );

    \I__7167\ : InMux
    port map (
            O => \N__32352\,
            I => \N__32325\
        );

    \I__7166\ : Span4Mux_v
    port map (
            O => \N__32349\,
            I => \N__32320\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__32346\,
            I => \N__32320\
        );

    \I__7164\ : InMux
    port map (
            O => \N__32343\,
            I => \N__32317\
        );

    \I__7163\ : CascadeMux
    port map (
            O => \N__32342\,
            I => \N__32314\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__32339\,
            I => \N__32310\
        );

    \I__7161\ : InMux
    port map (
            O => \N__32336\,
            I => \N__32307\
        );

    \I__7160\ : InMux
    port map (
            O => \N__32333\,
            I => \N__32304\
        );

    \I__7159\ : CascadeMux
    port map (
            O => \N__32332\,
            I => \N__32301\
        );

    \I__7158\ : CascadeMux
    port map (
            O => \N__32331\,
            I => \N__32298\
        );

    \I__7157\ : Sp12to4
    port map (
            O => \N__32328\,
            I => \N__32293\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__32325\,
            I => \N__32290\
        );

    \I__7155\ : Span4Mux_h
    port map (
            O => \N__32320\,
            I => \N__32285\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__32317\,
            I => \N__32285\
        );

    \I__7153\ : InMux
    port map (
            O => \N__32314\,
            I => \N__32282\
        );

    \I__7152\ : CascadeMux
    port map (
            O => \N__32313\,
            I => \N__32279\
        );

    \I__7151\ : Span4Mux_v
    port map (
            O => \N__32310\,
            I => \N__32272\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__32307\,
            I => \N__32272\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__32304\,
            I => \N__32272\
        );

    \I__7148\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32269\
        );

    \I__7147\ : InMux
    port map (
            O => \N__32298\,
            I => \N__32266\
        );

    \I__7146\ : CascadeMux
    port map (
            O => \N__32297\,
            I => \N__32263\
        );

    \I__7145\ : CascadeMux
    port map (
            O => \N__32296\,
            I => \N__32260\
        );

    \I__7144\ : Span12Mux_h
    port map (
            O => \N__32293\,
            I => \N__32254\
        );

    \I__7143\ : Span12Mux_s9_h
    port map (
            O => \N__32290\,
            I => \N__32254\
        );

    \I__7142\ : Span4Mux_v
    port map (
            O => \N__32285\,
            I => \N__32249\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__32282\,
            I => \N__32249\
        );

    \I__7140\ : InMux
    port map (
            O => \N__32279\,
            I => \N__32246\
        );

    \I__7139\ : Span4Mux_v
    port map (
            O => \N__32272\,
            I => \N__32239\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__32269\,
            I => \N__32239\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__32266\,
            I => \N__32239\
        );

    \I__7136\ : InMux
    port map (
            O => \N__32263\,
            I => \N__32236\
        );

    \I__7135\ : InMux
    port map (
            O => \N__32260\,
            I => \N__32233\
        );

    \I__7134\ : CascadeMux
    port map (
            O => \N__32259\,
            I => \N__32230\
        );

    \I__7133\ : Span12Mux_v
    port map (
            O => \N__32254\,
            I => \N__32227\
        );

    \I__7132\ : Span4Mux_h
    port map (
            O => \N__32249\,
            I => \N__32222\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__32246\,
            I => \N__32222\
        );

    \I__7130\ : Span4Mux_v
    port map (
            O => \N__32239\,
            I => \N__32215\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__32236\,
            I => \N__32215\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__32233\,
            I => \N__32215\
        );

    \I__7127\ : InMux
    port map (
            O => \N__32230\,
            I => \N__32212\
        );

    \I__7126\ : Span12Mux_h
    port map (
            O => \N__32227\,
            I => \N__32208\
        );

    \I__7125\ : Span4Mux_v
    port map (
            O => \N__32222\,
            I => \N__32201\
        );

    \I__7124\ : Span4Mux_v
    port map (
            O => \N__32215\,
            I => \N__32201\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__32212\,
            I => \N__32201\
        );

    \I__7122\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32198\
        );

    \I__7121\ : Odrv12
    port map (
            O => \N__32208\,
            I => \M_this_spr_address_qZ0Z_2\
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__32201\,
            I => \M_this_spr_address_qZ0Z_2\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__32198\,
            I => \M_this_spr_address_qZ0Z_2\
        );

    \I__7118\ : InMux
    port map (
            O => \N__32191\,
            I => \un1_M_this_spr_address_q_cry_1\
        );

    \I__7117\ : CascadeMux
    port map (
            O => \N__32188\,
            I => \N__32184\
        );

    \I__7116\ : CascadeMux
    port map (
            O => \N__32187\,
            I => \N__32179\
        );

    \I__7115\ : InMux
    port map (
            O => \N__32184\,
            I => \N__32176\
        );

    \I__7114\ : CascadeMux
    port map (
            O => \N__32183\,
            I => \N__32173\
        );

    \I__7113\ : CascadeMux
    port map (
            O => \N__32182\,
            I => \N__32167\
        );

    \I__7112\ : InMux
    port map (
            O => \N__32179\,
            I => \N__32163\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__32176\,
            I => \N__32160\
        );

    \I__7110\ : InMux
    port map (
            O => \N__32173\,
            I => \N__32157\
        );

    \I__7109\ : CascadeMux
    port map (
            O => \N__32172\,
            I => \N__32154\
        );

    \I__7108\ : CascadeMux
    port map (
            O => \N__32171\,
            I => \N__32151\
        );

    \I__7107\ : CascadeMux
    port map (
            O => \N__32170\,
            I => \N__32146\
        );

    \I__7106\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32143\
        );

    \I__7105\ : CascadeMux
    port map (
            O => \N__32166\,
            I => \N__32140\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__32163\,
            I => \N__32135\
        );

    \I__7103\ : Span4Mux_h
    port map (
            O => \N__32160\,
            I => \N__32132\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__32157\,
            I => \N__32129\
        );

    \I__7101\ : InMux
    port map (
            O => \N__32154\,
            I => \N__32126\
        );

    \I__7100\ : InMux
    port map (
            O => \N__32151\,
            I => \N__32123\
        );

    \I__7099\ : CascadeMux
    port map (
            O => \N__32150\,
            I => \N__32120\
        );

    \I__7098\ : CascadeMux
    port map (
            O => \N__32149\,
            I => \N__32117\
        );

    \I__7097\ : InMux
    port map (
            O => \N__32146\,
            I => \N__32113\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__32143\,
            I => \N__32110\
        );

    \I__7095\ : InMux
    port map (
            O => \N__32140\,
            I => \N__32107\
        );

    \I__7094\ : CascadeMux
    port map (
            O => \N__32139\,
            I => \N__32104\
        );

    \I__7093\ : CascadeMux
    port map (
            O => \N__32138\,
            I => \N__32101\
        );

    \I__7092\ : Span4Mux_h
    port map (
            O => \N__32135\,
            I => \N__32096\
        );

    \I__7091\ : Span4Mux_v
    port map (
            O => \N__32132\,
            I => \N__32091\
        );

    \I__7090\ : Span4Mux_h
    port map (
            O => \N__32129\,
            I => \N__32091\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__32126\,
            I => \N__32088\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__32123\,
            I => \N__32085\
        );

    \I__7087\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32082\
        );

    \I__7086\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32079\
        );

    \I__7085\ : CascadeMux
    port map (
            O => \N__32116\,
            I => \N__32076\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__32113\,
            I => \N__32073\
        );

    \I__7083\ : Span4Mux_v
    port map (
            O => \N__32110\,
            I => \N__32068\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__32107\,
            I => \N__32068\
        );

    \I__7081\ : InMux
    port map (
            O => \N__32104\,
            I => \N__32065\
        );

    \I__7080\ : InMux
    port map (
            O => \N__32101\,
            I => \N__32062\
        );

    \I__7079\ : CascadeMux
    port map (
            O => \N__32100\,
            I => \N__32059\
        );

    \I__7078\ : CascadeMux
    port map (
            O => \N__32099\,
            I => \N__32056\
        );

    \I__7077\ : Sp12to4
    port map (
            O => \N__32096\,
            I => \N__32050\
        );

    \I__7076\ : Sp12to4
    port map (
            O => \N__32091\,
            I => \N__32050\
        );

    \I__7075\ : Span4Mux_v
    port map (
            O => \N__32088\,
            I => \N__32043\
        );

    \I__7074\ : Span4Mux_h
    port map (
            O => \N__32085\,
            I => \N__32043\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__32082\,
            I => \N__32043\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__32079\,
            I => \N__32040\
        );

    \I__7071\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32037\
        );

    \I__7070\ : Span4Mux_v
    port map (
            O => \N__32073\,
            I => \N__32028\
        );

    \I__7069\ : Span4Mux_v
    port map (
            O => \N__32068\,
            I => \N__32028\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__32065\,
            I => \N__32028\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__32062\,
            I => \N__32028\
        );

    \I__7066\ : InMux
    port map (
            O => \N__32059\,
            I => \N__32025\
        );

    \I__7065\ : InMux
    port map (
            O => \N__32056\,
            I => \N__32022\
        );

    \I__7064\ : CascadeMux
    port map (
            O => \N__32055\,
            I => \N__32019\
        );

    \I__7063\ : Span12Mux_v
    port map (
            O => \N__32050\,
            I => \N__32016\
        );

    \I__7062\ : Span4Mux_v
    port map (
            O => \N__32043\,
            I => \N__32009\
        );

    \I__7061\ : Span4Mux_h
    port map (
            O => \N__32040\,
            I => \N__32009\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__32037\,
            I => \N__32009\
        );

    \I__7059\ : Span4Mux_v
    port map (
            O => \N__32028\,
            I => \N__32002\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__32025\,
            I => \N__32002\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__32022\,
            I => \N__32002\
        );

    \I__7056\ : InMux
    port map (
            O => \N__32019\,
            I => \N__31999\
        );

    \I__7055\ : Span12Mux_h
    port map (
            O => \N__32016\,
            I => \N__31995\
        );

    \I__7054\ : Span4Mux_v
    port map (
            O => \N__32009\,
            I => \N__31990\
        );

    \I__7053\ : Span4Mux_v
    port map (
            O => \N__32002\,
            I => \N__31990\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__31999\,
            I => \N__31987\
        );

    \I__7051\ : InMux
    port map (
            O => \N__31998\,
            I => \N__31984\
        );

    \I__7050\ : Odrv12
    port map (
            O => \N__31995\,
            I => \M_this_spr_address_qZ0Z_3\
        );

    \I__7049\ : Odrv4
    port map (
            O => \N__31990\,
            I => \M_this_spr_address_qZ0Z_3\
        );

    \I__7048\ : Odrv12
    port map (
            O => \N__31987\,
            I => \M_this_spr_address_qZ0Z_3\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__31984\,
            I => \M_this_spr_address_qZ0Z_3\
        );

    \I__7046\ : InMux
    port map (
            O => \N__31975\,
            I => \un1_M_this_spr_address_q_cry_2\
        );

    \I__7045\ : CascadeMux
    port map (
            O => \N__31972\,
            I => \N__31967\
        );

    \I__7044\ : CascadeMux
    port map (
            O => \N__31971\,
            I => \N__31963\
        );

    \I__7043\ : CascadeMux
    port map (
            O => \N__31970\,
            I => \N__31958\
        );

    \I__7042\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31955\
        );

    \I__7041\ : CascadeMux
    port map (
            O => \N__31966\,
            I => \N__31952\
        );

    \I__7040\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31949\
        );

    \I__7039\ : CascadeMux
    port map (
            O => \N__31962\,
            I => \N__31946\
        );

    \I__7038\ : CascadeMux
    port map (
            O => \N__31961\,
            I => \N__31942\
        );

    \I__7037\ : InMux
    port map (
            O => \N__31958\,
            I => \N__31937\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__31955\,
            I => \N__31934\
        );

    \I__7035\ : InMux
    port map (
            O => \N__31952\,
            I => \N__31931\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__31949\,
            I => \N__31928\
        );

    \I__7033\ : InMux
    port map (
            O => \N__31946\,
            I => \N__31925\
        );

    \I__7032\ : CascadeMux
    port map (
            O => \N__31945\,
            I => \N__31922\
        );

    \I__7031\ : InMux
    port map (
            O => \N__31942\,
            I => \N__31918\
        );

    \I__7030\ : CascadeMux
    port map (
            O => \N__31941\,
            I => \N__31915\
        );

    \I__7029\ : CascadeMux
    port map (
            O => \N__31940\,
            I => \N__31912\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__31937\,
            I => \N__31906\
        );

    \I__7027\ : Span4Mux_h
    port map (
            O => \N__31934\,
            I => \N__31903\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__31931\,
            I => \N__31900\
        );

    \I__7025\ : Span4Mux_v
    port map (
            O => \N__31928\,
            I => \N__31895\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__31925\,
            I => \N__31895\
        );

    \I__7023\ : InMux
    port map (
            O => \N__31922\,
            I => \N__31892\
        );

    \I__7022\ : CascadeMux
    port map (
            O => \N__31921\,
            I => \N__31889\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__31918\,
            I => \N__31885\
        );

    \I__7020\ : InMux
    port map (
            O => \N__31915\,
            I => \N__31882\
        );

    \I__7019\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31879\
        );

    \I__7018\ : CascadeMux
    port map (
            O => \N__31911\,
            I => \N__31876\
        );

    \I__7017\ : CascadeMux
    port map (
            O => \N__31910\,
            I => \N__31873\
        );

    \I__7016\ : CascadeMux
    port map (
            O => \N__31909\,
            I => \N__31870\
        );

    \I__7015\ : Span4Mux_h
    port map (
            O => \N__31906\,
            I => \N__31866\
        );

    \I__7014\ : Span4Mux_v
    port map (
            O => \N__31903\,
            I => \N__31861\
        );

    \I__7013\ : Span4Mux_h
    port map (
            O => \N__31900\,
            I => \N__31861\
        );

    \I__7012\ : Span4Mux_h
    port map (
            O => \N__31895\,
            I => \N__31856\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__31892\,
            I => \N__31856\
        );

    \I__7010\ : InMux
    port map (
            O => \N__31889\,
            I => \N__31853\
        );

    \I__7009\ : CascadeMux
    port map (
            O => \N__31888\,
            I => \N__31850\
        );

    \I__7008\ : Span4Mux_v
    port map (
            O => \N__31885\,
            I => \N__31843\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__31882\,
            I => \N__31843\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__31879\,
            I => \N__31843\
        );

    \I__7005\ : InMux
    port map (
            O => \N__31876\,
            I => \N__31840\
        );

    \I__7004\ : InMux
    port map (
            O => \N__31873\,
            I => \N__31837\
        );

    \I__7003\ : InMux
    port map (
            O => \N__31870\,
            I => \N__31834\
        );

    \I__7002\ : CascadeMux
    port map (
            O => \N__31869\,
            I => \N__31831\
        );

    \I__7001\ : Sp12to4
    port map (
            O => \N__31866\,
            I => \N__31825\
        );

    \I__7000\ : Sp12to4
    port map (
            O => \N__31861\,
            I => \N__31825\
        );

    \I__6999\ : Span4Mux_v
    port map (
            O => \N__31856\,
            I => \N__31820\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__31853\,
            I => \N__31820\
        );

    \I__6997\ : InMux
    port map (
            O => \N__31850\,
            I => \N__31817\
        );

    \I__6996\ : Span4Mux_v
    port map (
            O => \N__31843\,
            I => \N__31812\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__31840\,
            I => \N__31812\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__31837\,
            I => \N__31809\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__31834\,
            I => \N__31806\
        );

    \I__6992\ : InMux
    port map (
            O => \N__31831\,
            I => \N__31803\
        );

    \I__6991\ : CascadeMux
    port map (
            O => \N__31830\,
            I => \N__31800\
        );

    \I__6990\ : Span12Mux_v
    port map (
            O => \N__31825\,
            I => \N__31797\
        );

    \I__6989\ : Span4Mux_h
    port map (
            O => \N__31820\,
            I => \N__31792\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__31817\,
            I => \N__31792\
        );

    \I__6987\ : Span4Mux_v
    port map (
            O => \N__31812\,
            I => \N__31783\
        );

    \I__6986\ : Span4Mux_v
    port map (
            O => \N__31809\,
            I => \N__31783\
        );

    \I__6985\ : Span4Mux_h
    port map (
            O => \N__31806\,
            I => \N__31783\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__31803\,
            I => \N__31783\
        );

    \I__6983\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31780\
        );

    \I__6982\ : Span12Mux_h
    port map (
            O => \N__31797\,
            I => \N__31776\
        );

    \I__6981\ : Span4Mux_v
    port map (
            O => \N__31792\,
            I => \N__31769\
        );

    \I__6980\ : Span4Mux_v
    port map (
            O => \N__31783\,
            I => \N__31769\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__31780\,
            I => \N__31769\
        );

    \I__6978\ : InMux
    port map (
            O => \N__31779\,
            I => \N__31766\
        );

    \I__6977\ : Odrv12
    port map (
            O => \N__31776\,
            I => \M_this_spr_address_qZ0Z_4\
        );

    \I__6976\ : Odrv4
    port map (
            O => \N__31769\,
            I => \M_this_spr_address_qZ0Z_4\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__31766\,
            I => \M_this_spr_address_qZ0Z_4\
        );

    \I__6974\ : InMux
    port map (
            O => \N__31759\,
            I => \un1_M_this_spr_address_q_cry_3\
        );

    \I__6973\ : CascadeMux
    port map (
            O => \N__31756\,
            I => \N__31752\
        );

    \I__6972\ : CascadeMux
    port map (
            O => \N__31755\,
            I => \N__31749\
        );

    \I__6971\ : InMux
    port map (
            O => \N__31752\,
            I => \N__31743\
        );

    \I__6970\ : InMux
    port map (
            O => \N__31749\,
            I => \N__31740\
        );

    \I__6969\ : CascadeMux
    port map (
            O => \N__31748\,
            I => \N__31737\
        );

    \I__6968\ : CascadeMux
    port map (
            O => \N__31747\,
            I => \N__31732\
        );

    \I__6967\ : CascadeMux
    port map (
            O => \N__31746\,
            I => \N__31729\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__31743\,
            I => \N__31724\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__31740\,
            I => \N__31721\
        );

    \I__6964\ : InMux
    port map (
            O => \N__31737\,
            I => \N__31718\
        );

    \I__6963\ : CascadeMux
    port map (
            O => \N__31736\,
            I => \N__31715\
        );

    \I__6962\ : CascadeMux
    port map (
            O => \N__31735\,
            I => \N__31709\
        );

    \I__6961\ : InMux
    port map (
            O => \N__31732\,
            I => \N__31704\
        );

    \I__6960\ : InMux
    port map (
            O => \N__31729\,
            I => \N__31701\
        );

    \I__6959\ : CascadeMux
    port map (
            O => \N__31728\,
            I => \N__31698\
        );

    \I__6958\ : CascadeMux
    port map (
            O => \N__31727\,
            I => \N__31695\
        );

    \I__6957\ : Span4Mux_s2_v
    port map (
            O => \N__31724\,
            I => \N__31687\
        );

    \I__6956\ : Span4Mux_h
    port map (
            O => \N__31721\,
            I => \N__31687\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__31718\,
            I => \N__31687\
        );

    \I__6954\ : InMux
    port map (
            O => \N__31715\,
            I => \N__31684\
        );

    \I__6953\ : CascadeMux
    port map (
            O => \N__31714\,
            I => \N__31681\
        );

    \I__6952\ : CascadeMux
    port map (
            O => \N__31713\,
            I => \N__31678\
        );

    \I__6951\ : CascadeMux
    port map (
            O => \N__31712\,
            I => \N__31675\
        );

    \I__6950\ : InMux
    port map (
            O => \N__31709\,
            I => \N__31672\
        );

    \I__6949\ : CascadeMux
    port map (
            O => \N__31708\,
            I => \N__31669\
        );

    \I__6948\ : CascadeMux
    port map (
            O => \N__31707\,
            I => \N__31666\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__31704\,
            I => \N__31661\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__31701\,
            I => \N__31661\
        );

    \I__6945\ : InMux
    port map (
            O => \N__31698\,
            I => \N__31658\
        );

    \I__6944\ : InMux
    port map (
            O => \N__31695\,
            I => \N__31655\
        );

    \I__6943\ : CascadeMux
    port map (
            O => \N__31694\,
            I => \N__31652\
        );

    \I__6942\ : Span4Mux_v
    port map (
            O => \N__31687\,
            I => \N__31649\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__31684\,
            I => \N__31645\
        );

    \I__6940\ : InMux
    port map (
            O => \N__31681\,
            I => \N__31642\
        );

    \I__6939\ : InMux
    port map (
            O => \N__31678\,
            I => \N__31639\
        );

    \I__6938\ : InMux
    port map (
            O => \N__31675\,
            I => \N__31636\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__31672\,
            I => \N__31633\
        );

    \I__6936\ : InMux
    port map (
            O => \N__31669\,
            I => \N__31630\
        );

    \I__6935\ : InMux
    port map (
            O => \N__31666\,
            I => \N__31627\
        );

    \I__6934\ : Span4Mux_v
    port map (
            O => \N__31661\,
            I => \N__31620\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__31658\,
            I => \N__31620\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__31655\,
            I => \N__31620\
        );

    \I__6931\ : InMux
    port map (
            O => \N__31652\,
            I => \N__31617\
        );

    \I__6930\ : Sp12to4
    port map (
            O => \N__31649\,
            I => \N__31614\
        );

    \I__6929\ : CascadeMux
    port map (
            O => \N__31648\,
            I => \N__31611\
        );

    \I__6928\ : Span12Mux_s6_v
    port map (
            O => \N__31645\,
            I => \N__31606\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__31642\,
            I => \N__31606\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__31639\,
            I => \N__31601\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__31636\,
            I => \N__31601\
        );

    \I__6924\ : Span4Mux_v
    port map (
            O => \N__31633\,
            I => \N__31596\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__31630\,
            I => \N__31596\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__31627\,
            I => \N__31593\
        );

    \I__6921\ : Span4Mux_v
    port map (
            O => \N__31620\,
            I => \N__31588\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__31617\,
            I => \N__31588\
        );

    \I__6919\ : Span12Mux_h
    port map (
            O => \N__31614\,
            I => \N__31585\
        );

    \I__6918\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31582\
        );

    \I__6917\ : Span12Mux_v
    port map (
            O => \N__31606\,
            I => \N__31576\
        );

    \I__6916\ : Span12Mux_v
    port map (
            O => \N__31601\,
            I => \N__31576\
        );

    \I__6915\ : Span4Mux_h
    port map (
            O => \N__31596\,
            I => \N__31573\
        );

    \I__6914\ : Span4Mux_h
    port map (
            O => \N__31593\,
            I => \N__31568\
        );

    \I__6913\ : Span4Mux_h
    port map (
            O => \N__31588\,
            I => \N__31568\
        );

    \I__6912\ : Span12Mux_v
    port map (
            O => \N__31585\,
            I => \N__31563\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__31582\,
            I => \N__31563\
        );

    \I__6910\ : InMux
    port map (
            O => \N__31581\,
            I => \N__31560\
        );

    \I__6909\ : Odrv12
    port map (
            O => \N__31576\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__6908\ : Odrv4
    port map (
            O => \N__31573\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__31568\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__6906\ : Odrv12
    port map (
            O => \N__31563\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__31560\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__6904\ : InMux
    port map (
            O => \N__31549\,
            I => \un1_M_this_spr_address_q_cry_4\
        );

    \I__6903\ : CascadeMux
    port map (
            O => \N__31546\,
            I => \N__31540\
        );

    \I__6902\ : CascadeMux
    port map (
            O => \N__31545\,
            I => \N__31535\
        );

    \I__6901\ : CascadeMux
    port map (
            O => \N__31544\,
            I => \N__31530\
        );

    \I__6900\ : CascadeMux
    port map (
            O => \N__31543\,
            I => \N__31527\
        );

    \I__6899\ : InMux
    port map (
            O => \N__31540\,
            I => \N__31522\
        );

    \I__6898\ : CascadeMux
    port map (
            O => \N__31539\,
            I => \N__31519\
        );

    \I__6897\ : CascadeMux
    port map (
            O => \N__31538\,
            I => \N__31516\
        );

    \I__6896\ : InMux
    port map (
            O => \N__31535\,
            I => \N__31511\
        );

    \I__6895\ : CascadeMux
    port map (
            O => \N__31534\,
            I => \N__31508\
        );

    \I__6894\ : CascadeMux
    port map (
            O => \N__31533\,
            I => \N__31505\
        );

    \I__6893\ : InMux
    port map (
            O => \N__31530\,
            I => \N__31502\
        );

    \I__6892\ : InMux
    port map (
            O => \N__31527\,
            I => \N__31499\
        );

    \I__6891\ : CascadeMux
    port map (
            O => \N__31526\,
            I => \N__31496\
        );

    \I__6890\ : CascadeMux
    port map (
            O => \N__31525\,
            I => \N__31493\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__31522\,
            I => \N__31489\
        );

    \I__6888\ : InMux
    port map (
            O => \N__31519\,
            I => \N__31486\
        );

    \I__6887\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31483\
        );

    \I__6886\ : CascadeMux
    port map (
            O => \N__31515\,
            I => \N__31480\
        );

    \I__6885\ : CascadeMux
    port map (
            O => \N__31514\,
            I => \N__31477\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__31511\,
            I => \N__31472\
        );

    \I__6883\ : InMux
    port map (
            O => \N__31508\,
            I => \N__31469\
        );

    \I__6882\ : InMux
    port map (
            O => \N__31505\,
            I => \N__31466\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__31502\,
            I => \N__31463\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__31499\,
            I => \N__31460\
        );

    \I__6879\ : InMux
    port map (
            O => \N__31496\,
            I => \N__31457\
        );

    \I__6878\ : InMux
    port map (
            O => \N__31493\,
            I => \N__31454\
        );

    \I__6877\ : CascadeMux
    port map (
            O => \N__31492\,
            I => \N__31451\
        );

    \I__6876\ : Span4Mux_v
    port map (
            O => \N__31489\,
            I => \N__31444\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__31486\,
            I => \N__31444\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__31483\,
            I => \N__31444\
        );

    \I__6873\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31441\
        );

    \I__6872\ : InMux
    port map (
            O => \N__31477\,
            I => \N__31438\
        );

    \I__6871\ : CascadeMux
    port map (
            O => \N__31476\,
            I => \N__31435\
        );

    \I__6870\ : CascadeMux
    port map (
            O => \N__31475\,
            I => \N__31432\
        );

    \I__6869\ : Sp12to4
    port map (
            O => \N__31472\,
            I => \N__31425\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__31469\,
            I => \N__31425\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__31466\,
            I => \N__31425\
        );

    \I__6866\ : Span4Mux_v
    port map (
            O => \N__31463\,
            I => \N__31417\
        );

    \I__6865\ : Span4Mux_h
    port map (
            O => \N__31460\,
            I => \N__31417\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__31457\,
            I => \N__31417\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__31454\,
            I => \N__31414\
        );

    \I__6862\ : InMux
    port map (
            O => \N__31451\,
            I => \N__31411\
        );

    \I__6861\ : Span4Mux_v
    port map (
            O => \N__31444\,
            I => \N__31404\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__31441\,
            I => \N__31404\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__31438\,
            I => \N__31404\
        );

    \I__6858\ : InMux
    port map (
            O => \N__31435\,
            I => \N__31401\
        );

    \I__6857\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31398\
        );

    \I__6856\ : Span12Mux_s6_v
    port map (
            O => \N__31425\,
            I => \N__31395\
        );

    \I__6855\ : CascadeMux
    port map (
            O => \N__31424\,
            I => \N__31392\
        );

    \I__6854\ : Span4Mux_v
    port map (
            O => \N__31417\,
            I => \N__31385\
        );

    \I__6853\ : Span4Mux_h
    port map (
            O => \N__31414\,
            I => \N__31385\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__31411\,
            I => \N__31385\
        );

    \I__6851\ : Span4Mux_v
    port map (
            O => \N__31404\,
            I => \N__31378\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__31401\,
            I => \N__31378\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__31398\,
            I => \N__31378\
        );

    \I__6848\ : Span12Mux_v
    port map (
            O => \N__31395\,
            I => \N__31375\
        );

    \I__6847\ : InMux
    port map (
            O => \N__31392\,
            I => \N__31372\
        );

    \I__6846\ : Span4Mux_v
    port map (
            O => \N__31385\,
            I => \N__31366\
        );

    \I__6845\ : Span4Mux_v
    port map (
            O => \N__31378\,
            I => \N__31366\
        );

    \I__6844\ : Span12Mux_h
    port map (
            O => \N__31375\,
            I => \N__31361\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__31372\,
            I => \N__31361\
        );

    \I__6842\ : InMux
    port map (
            O => \N__31371\,
            I => \N__31358\
        );

    \I__6841\ : Odrv4
    port map (
            O => \N__31366\,
            I => \M_this_spr_address_qZ0Z_6\
        );

    \I__6840\ : Odrv12
    port map (
            O => \N__31361\,
            I => \M_this_spr_address_qZ0Z_6\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__31358\,
            I => \M_this_spr_address_qZ0Z_6\
        );

    \I__6838\ : InMux
    port map (
            O => \N__31351\,
            I => \un1_M_this_spr_address_q_cry_5\
        );

    \I__6837\ : CascadeMux
    port map (
            O => \N__31348\,
            I => \N__31344\
        );

    \I__6836\ : CascadeMux
    port map (
            O => \N__31347\,
            I => \N__31341\
        );

    \I__6835\ : InMux
    port map (
            O => \N__31344\,
            I => \N__31334\
        );

    \I__6834\ : InMux
    port map (
            O => \N__31341\,
            I => \N__31331\
        );

    \I__6833\ : CascadeMux
    port map (
            O => \N__31340\,
            I => \N__31328\
        );

    \I__6832\ : CascadeMux
    port map (
            O => \N__31339\,
            I => \N__31325\
        );

    \I__6831\ : CascadeMux
    port map (
            O => \N__31338\,
            I => \N__31320\
        );

    \I__6830\ : CascadeMux
    port map (
            O => \N__31337\,
            I => \N__31317\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__31334\,
            I => \N__31312\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__31331\,
            I => \N__31309\
        );

    \I__6827\ : InMux
    port map (
            O => \N__31328\,
            I => \N__31306\
        );

    \I__6826\ : InMux
    port map (
            O => \N__31325\,
            I => \N__31303\
        );

    \I__6825\ : CascadeMux
    port map (
            O => \N__31324\,
            I => \N__31300\
        );

    \I__6824\ : CascadeMux
    port map (
            O => \N__31323\,
            I => \N__31297\
        );

    \I__6823\ : InMux
    port map (
            O => \N__31320\,
            I => \N__31292\
        );

    \I__6822\ : InMux
    port map (
            O => \N__31317\,
            I => \N__31289\
        );

    \I__6821\ : CascadeMux
    port map (
            O => \N__31316\,
            I => \N__31286\
        );

    \I__6820\ : CascadeMux
    port map (
            O => \N__31315\,
            I => \N__31283\
        );

    \I__6819\ : Span4Mux_s2_v
    port map (
            O => \N__31312\,
            I => \N__31277\
        );

    \I__6818\ : Span4Mux_h
    port map (
            O => \N__31309\,
            I => \N__31277\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__31306\,
            I => \N__31274\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__31303\,
            I => \N__31271\
        );

    \I__6815\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31268\
        );

    \I__6814\ : InMux
    port map (
            O => \N__31297\,
            I => \N__31265\
        );

    \I__6813\ : CascadeMux
    port map (
            O => \N__31296\,
            I => \N__31262\
        );

    \I__6812\ : CascadeMux
    port map (
            O => \N__31295\,
            I => \N__31259\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__31292\,
            I => \N__31255\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__31289\,
            I => \N__31252\
        );

    \I__6809\ : InMux
    port map (
            O => \N__31286\,
            I => \N__31249\
        );

    \I__6808\ : InMux
    port map (
            O => \N__31283\,
            I => \N__31246\
        );

    \I__6807\ : CascadeMux
    port map (
            O => \N__31282\,
            I => \N__31243\
        );

    \I__6806\ : Span4Mux_v
    port map (
            O => \N__31277\,
            I => \N__31236\
        );

    \I__6805\ : Span4Mux_v
    port map (
            O => \N__31274\,
            I => \N__31236\
        );

    \I__6804\ : Span4Mux_v
    port map (
            O => \N__31271\,
            I => \N__31229\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__31268\,
            I => \N__31229\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__31265\,
            I => \N__31229\
        );

    \I__6801\ : InMux
    port map (
            O => \N__31262\,
            I => \N__31226\
        );

    \I__6800\ : InMux
    port map (
            O => \N__31259\,
            I => \N__31223\
        );

    \I__6799\ : CascadeMux
    port map (
            O => \N__31258\,
            I => \N__31220\
        );

    \I__6798\ : Span4Mux_v
    port map (
            O => \N__31255\,
            I => \N__31213\
        );

    \I__6797\ : Span4Mux_h
    port map (
            O => \N__31252\,
            I => \N__31213\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__31249\,
            I => \N__31213\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__31246\,
            I => \N__31210\
        );

    \I__6794\ : InMux
    port map (
            O => \N__31243\,
            I => \N__31207\
        );

    \I__6793\ : CascadeMux
    port map (
            O => \N__31242\,
            I => \N__31204\
        );

    \I__6792\ : CascadeMux
    port map (
            O => \N__31241\,
            I => \N__31201\
        );

    \I__6791\ : Sp12to4
    port map (
            O => \N__31236\,
            I => \N__31198\
        );

    \I__6790\ : Span4Mux_v
    port map (
            O => \N__31229\,
            I => \N__31191\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__31226\,
            I => \N__31191\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__31223\,
            I => \N__31191\
        );

    \I__6787\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31188\
        );

    \I__6786\ : Span4Mux_v
    port map (
            O => \N__31213\,
            I => \N__31181\
        );

    \I__6785\ : Span4Mux_h
    port map (
            O => \N__31210\,
            I => \N__31181\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__31207\,
            I => \N__31181\
        );

    \I__6783\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31178\
        );

    \I__6782\ : InMux
    port map (
            O => \N__31201\,
            I => \N__31175\
        );

    \I__6781\ : Span12Mux_h
    port map (
            O => \N__31198\,
            I => \N__31172\
        );

    \I__6780\ : Span4Mux_v
    port map (
            O => \N__31191\,
            I => \N__31163\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__31188\,
            I => \N__31163\
        );

    \I__6778\ : Span4Mux_v
    port map (
            O => \N__31181\,
            I => \N__31163\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__31178\,
            I => \N__31163\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__31175\,
            I => \N__31160\
        );

    \I__6775\ : Span12Mux_v
    port map (
            O => \N__31172\,
            I => \N__31156\
        );

    \I__6774\ : Span4Mux_v
    port map (
            O => \N__31163\,
            I => \N__31151\
        );

    \I__6773\ : Span4Mux_h
    port map (
            O => \N__31160\,
            I => \N__31151\
        );

    \I__6772\ : InMux
    port map (
            O => \N__31159\,
            I => \N__31148\
        );

    \I__6771\ : Odrv12
    port map (
            O => \N__31156\,
            I => \M_this_spr_address_qZ0Z_7\
        );

    \I__6770\ : Odrv4
    port map (
            O => \N__31151\,
            I => \M_this_spr_address_qZ0Z_7\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__31148\,
            I => \M_this_spr_address_qZ0Z_7\
        );

    \I__6768\ : InMux
    port map (
            O => \N__31141\,
            I => \un1_M_this_spr_address_q_cry_6\
        );

    \I__6767\ : InMux
    port map (
            O => \N__31138\,
            I => \N__31132\
        );

    \I__6766\ : InMux
    port map (
            O => \N__31137\,
            I => \N__31132\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__31132\,
            I => \this_ppu.N_1176_1\
        );

    \I__6764\ : InMux
    port map (
            O => \N__31129\,
            I => \N__31126\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__31126\,
            I => \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_3\
        );

    \I__6762\ : CascadeMux
    port map (
            O => \N__31123\,
            I => \N__31120\
        );

    \I__6761\ : InMux
    port map (
            O => \N__31120\,
            I => \N__31117\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__31117\,
            I => \N__31114\
        );

    \I__6759\ : Odrv4
    port map (
            O => \N__31114\,
            I => \this_ppu.N_893\
        );

    \I__6758\ : CascadeMux
    port map (
            O => \N__31111\,
            I => \N__31108\
        );

    \I__6757\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31105\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__31105\,
            I => \this_ppu.N_969\
        );

    \I__6755\ : CascadeMux
    port map (
            O => \N__31102\,
            I => \un1_M_this_state_q_11_0_0_cascade_\
        );

    \I__6754\ : CascadeMux
    port map (
            O => \N__31099\,
            I => \this_ppu.un1_M_this_state_q_11_0_0Z0Z_0_cascade_\
        );

    \I__6753\ : InMux
    port map (
            O => \N__31096\,
            I => \N__31093\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__31093\,
            I => \this_ppu.un1_M_this_state_q_11_0_0Z0Z_1\
        );

    \I__6751\ : CascadeMux
    port map (
            O => \N__31090\,
            I => \N__31085\
        );

    \I__6750\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31080\
        );

    \I__6749\ : InMux
    port map (
            O => \N__31088\,
            I => \N__31080\
        );

    \I__6748\ : InMux
    port map (
            O => \N__31085\,
            I => \N__31076\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__31080\,
            I => \N__31072\
        );

    \I__6746\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31069\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__31076\,
            I => \N__31060\
        );

    \I__6744\ : CascadeMux
    port map (
            O => \N__31075\,
            I => \N__31056\
        );

    \I__6743\ : Span4Mux_v
    port map (
            O => \N__31072\,
            I => \N__31049\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__31069\,
            I => \N__31049\
        );

    \I__6741\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31040\
        );

    \I__6740\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31040\
        );

    \I__6739\ : InMux
    port map (
            O => \N__31066\,
            I => \N__31040\
        );

    \I__6738\ : InMux
    port map (
            O => \N__31065\,
            I => \N__31040\
        );

    \I__6737\ : InMux
    port map (
            O => \N__31064\,
            I => \N__31035\
        );

    \I__6736\ : InMux
    port map (
            O => \N__31063\,
            I => \N__31035\
        );

    \I__6735\ : Span4Mux_v
    port map (
            O => \N__31060\,
            I => \N__31031\
        );

    \I__6734\ : InMux
    port map (
            O => \N__31059\,
            I => \N__31028\
        );

    \I__6733\ : InMux
    port map (
            O => \N__31056\,
            I => \N__31025\
        );

    \I__6732\ : InMux
    port map (
            O => \N__31055\,
            I => \N__31020\
        );

    \I__6731\ : InMux
    port map (
            O => \N__31054\,
            I => \N__31020\
        );

    \I__6730\ : Span4Mux_h
    port map (
            O => \N__31049\,
            I => \N__31017\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__31040\,
            I => \N__31012\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__31035\,
            I => \N__31012\
        );

    \I__6727\ : InMux
    port map (
            O => \N__31034\,
            I => \N__31009\
        );

    \I__6726\ : Odrv4
    port map (
            O => \N__31031\,
            I => \this_ppu.N_430_1_0\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__31028\,
            I => \this_ppu.N_430_1_0\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__31025\,
            I => \this_ppu.N_430_1_0\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__31020\,
            I => \this_ppu.N_430_1_0\
        );

    \I__6722\ : Odrv4
    port map (
            O => \N__31017\,
            I => \this_ppu.N_430_1_0\
        );

    \I__6721\ : Odrv12
    port map (
            O => \N__31012\,
            I => \this_ppu.N_430_1_0\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__31009\,
            I => \this_ppu.N_430_1_0\
        );

    \I__6719\ : CascadeMux
    port map (
            O => \N__30994\,
            I => \N__30991\
        );

    \I__6718\ : InMux
    port map (
            O => \N__30991\,
            I => \N__30987\
        );

    \I__6717\ : InMux
    port map (
            O => \N__30990\,
            I => \N__30984\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__30987\,
            I => \N__30981\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__30984\,
            I => \N__30978\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__30981\,
            I => \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_2\
        );

    \I__6713\ : Odrv4
    port map (
            O => \N__30978\,
            I => \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_2\
        );

    \I__6712\ : CascadeMux
    port map (
            O => \N__30973\,
            I => \this_ppu.N_1158_cascade_\
        );

    \I__6711\ : InMux
    port map (
            O => \N__30970\,
            I => \N__30966\
        );

    \I__6710\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30963\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__30966\,
            I => \N__30960\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__30963\,
            I => \this_ppu.N_1263\
        );

    \I__6707\ : Odrv4
    port map (
            O => \N__30960\,
            I => \this_ppu.N_1263\
        );

    \I__6706\ : CascadeMux
    port map (
            O => \N__30955\,
            I => \N__30952\
        );

    \I__6705\ : InMux
    port map (
            O => \N__30952\,
            I => \N__30949\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__30949\,
            I => \N__30946\
        );

    \I__6703\ : Odrv4
    port map (
            O => \N__30946\,
            I => \this_ppu.M_this_state_q_srsts_0_0_a3_1_2_1Z0Z_0\
        );

    \I__6702\ : InMux
    port map (
            O => \N__30943\,
            I => \N__30940\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__30940\,
            I => \this_ppu.M_this_state_q_srsts_0_0_0_tz_0_0\
        );

    \I__6700\ : InMux
    port map (
            O => \N__30937\,
            I => \N__30933\
        );

    \I__6699\ : InMux
    port map (
            O => \N__30936\,
            I => \N__30930\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__30933\,
            I => \N__30925\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__30930\,
            I => \N__30922\
        );

    \I__6696\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30919\
        );

    \I__6695\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30915\
        );

    \I__6694\ : Span4Mux_v
    port map (
            O => \N__30925\,
            I => \N__30910\
        );

    \I__6693\ : Span4Mux_v
    port map (
            O => \N__30922\,
            I => \N__30910\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__30919\,
            I => \N__30907\
        );

    \I__6691\ : InMux
    port map (
            O => \N__30918\,
            I => \N__30904\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__30915\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6689\ : Odrv4
    port map (
            O => \N__30910\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6688\ : Odrv4
    port map (
            O => \N__30907\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__30904\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6686\ : InMux
    port map (
            O => \N__30895\,
            I => \N__30892\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__30892\,
            I => \N__30889\
        );

    \I__6684\ : Span4Mux_h
    port map (
            O => \N__30889\,
            I => \N__30884\
        );

    \I__6683\ : InMux
    port map (
            O => \N__30888\,
            I => \N__30881\
        );

    \I__6682\ : InMux
    port map (
            O => \N__30887\,
            I => \N__30878\
        );

    \I__6681\ : Odrv4
    port map (
            O => \N__30884\,
            I => \N_815_0\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__30881\,
            I => \N_815_0\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__30878\,
            I => \N_815_0\
        );

    \I__6678\ : IoInMux
    port map (
            O => \N__30871\,
            I => \N__30868\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__30868\,
            I => \N__30865\
        );

    \I__6676\ : IoSpan4Mux
    port map (
            O => \N__30865\,
            I => \N__30862\
        );

    \I__6675\ : Span4Mux_s3_h
    port map (
            O => \N__30862\,
            I => \N__30859\
        );

    \I__6674\ : Sp12to4
    port map (
            O => \N__30859\,
            I => \N__30856\
        );

    \I__6673\ : Span12Mux_s11_h
    port map (
            O => \N__30856\,
            I => \N__30853\
        );

    \I__6672\ : Span12Mux_v
    port map (
            O => \N__30853\,
            I => \N__30850\
        );

    \I__6671\ : Odrv12
    port map (
            O => \N__30850\,
            I => led_c_7
        );

    \I__6670\ : CascadeMux
    port map (
            O => \N__30847\,
            I => \N__30844\
        );

    \I__6669\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30841\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__30841\,
            I => \this_ppu.N_807_0\
        );

    \I__6667\ : InMux
    port map (
            O => \N__30838\,
            I => \N__30828\
        );

    \I__6666\ : InMux
    port map (
            O => \N__30837\,
            I => \N__30828\
        );

    \I__6665\ : InMux
    port map (
            O => \N__30836\,
            I => \N__30825\
        );

    \I__6664\ : InMux
    port map (
            O => \N__30835\,
            I => \N__30822\
        );

    \I__6663\ : InMux
    port map (
            O => \N__30834\,
            I => \N__30819\
        );

    \I__6662\ : InMux
    port map (
            O => \N__30833\,
            I => \N__30816\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__30828\,
            I => \M_this_state_qZ0Z_16\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__30825\,
            I => \M_this_state_qZ0Z_16\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__30822\,
            I => \M_this_state_qZ0Z_16\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__30819\,
            I => \M_this_state_qZ0Z_16\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__30816\,
            I => \M_this_state_qZ0Z_16\
        );

    \I__6656\ : InMux
    port map (
            O => \N__30805\,
            I => \N__30802\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__30802\,
            I => \N__30799\
        );

    \I__6654\ : Odrv12
    port map (
            O => \N__30799\,
            I => \N_1415\
        );

    \I__6653\ : CascadeMux
    port map (
            O => \N__30796\,
            I => \N_1415_cascade_\
        );

    \I__6652\ : InMux
    port map (
            O => \N__30793\,
            I => \N__30785\
        );

    \I__6651\ : InMux
    port map (
            O => \N__30792\,
            I => \N__30785\
        );

    \I__6650\ : InMux
    port map (
            O => \N__30791\,
            I => \N__30780\
        );

    \I__6649\ : InMux
    port map (
            O => \N__30790\,
            I => \N__30780\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__30785\,
            I => \this_ppu.N_1278\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__30780\,
            I => \this_ppu.N_1278\
        );

    \I__6646\ : InMux
    port map (
            O => \N__30775\,
            I => \N__30772\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__30772\,
            I => \this_ppu.N_1166\
        );

    \I__6644\ : CascadeMux
    port map (
            O => \N__30769\,
            I => \this_ppu.N_1263_cascade_\
        );

    \I__6643\ : InMux
    port map (
            O => \N__30766\,
            I => \N__30763\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__30763\,
            I => \N__30759\
        );

    \I__6641\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30756\
        );

    \I__6640\ : Span4Mux_h
    port map (
            O => \N__30759\,
            I => \N__30752\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__30756\,
            I => \N__30749\
        );

    \I__6638\ : InMux
    port map (
            O => \N__30755\,
            I => \N__30746\
        );

    \I__6637\ : Span4Mux_v
    port map (
            O => \N__30752\,
            I => \N__30743\
        );

    \I__6636\ : Span4Mux_v
    port map (
            O => \N__30749\,
            I => \N__30740\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__30746\,
            I => \N__30737\
        );

    \I__6634\ : Odrv4
    port map (
            O => \N__30743\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__6633\ : Odrv4
    port map (
            O => \N__30740\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__6632\ : Odrv12
    port map (
            O => \N__30737\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__6631\ : InMux
    port map (
            O => \N__30730\,
            I => \N__30727\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__30727\,
            I => \N__30722\
        );

    \I__6629\ : InMux
    port map (
            O => \N__30726\,
            I => \N__30719\
        );

    \I__6628\ : InMux
    port map (
            O => \N__30725\,
            I => \N__30716\
        );

    \I__6627\ : Span4Mux_v
    port map (
            O => \N__30722\,
            I => \N__30711\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__30719\,
            I => \N__30711\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__30716\,
            I => \N__30708\
        );

    \I__6624\ : Span4Mux_v
    port map (
            O => \N__30711\,
            I => \N__30705\
        );

    \I__6623\ : Odrv12
    port map (
            O => \N__30708\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__6622\ : Odrv4
    port map (
            O => \N__30705\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__6621\ : InMux
    port map (
            O => \N__30700\,
            I => \N__30694\
        );

    \I__6620\ : InMux
    port map (
            O => \N__30699\,
            I => \N__30694\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__30694\,
            I => \N__30689\
        );

    \I__6618\ : InMux
    port map (
            O => \N__30693\,
            I => \N__30680\
        );

    \I__6617\ : InMux
    port map (
            O => \N__30692\,
            I => \N__30677\
        );

    \I__6616\ : Span4Mux_v
    port map (
            O => \N__30689\,
            I => \N__30674\
        );

    \I__6615\ : InMux
    port map (
            O => \N__30688\,
            I => \N__30671\
        );

    \I__6614\ : InMux
    port map (
            O => \N__30687\,
            I => \N__30664\
        );

    \I__6613\ : InMux
    port map (
            O => \N__30686\,
            I => \N__30664\
        );

    \I__6612\ : InMux
    port map (
            O => \N__30685\,
            I => \N__30661\
        );

    \I__6611\ : InMux
    port map (
            O => \N__30684\,
            I => \N__30656\
        );

    \I__6610\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30656\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__30680\,
            I => \N__30653\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__30677\,
            I => \N__30648\
        );

    \I__6607\ : Span4Mux_h
    port map (
            O => \N__30674\,
            I => \N__30645\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__30671\,
            I => \N__30642\
        );

    \I__6605\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30639\
        );

    \I__6604\ : InMux
    port map (
            O => \N__30669\,
            I => \N__30634\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__30664\,
            I => \N__30627\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__30661\,
            I => \N__30627\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__30656\,
            I => \N__30627\
        );

    \I__6600\ : Span4Mux_v
    port map (
            O => \N__30653\,
            I => \N__30624\
        );

    \I__6599\ : InMux
    port map (
            O => \N__30652\,
            I => \N__30619\
        );

    \I__6598\ : InMux
    port map (
            O => \N__30651\,
            I => \N__30619\
        );

    \I__6597\ : Span4Mux_v
    port map (
            O => \N__30648\,
            I => \N__30610\
        );

    \I__6596\ : Span4Mux_h
    port map (
            O => \N__30645\,
            I => \N__30610\
        );

    \I__6595\ : Span4Mux_v
    port map (
            O => \N__30642\,
            I => \N__30610\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__30639\,
            I => \N__30610\
        );

    \I__6593\ : InMux
    port map (
            O => \N__30638\,
            I => \N__30605\
        );

    \I__6592\ : InMux
    port map (
            O => \N__30637\,
            I => \N__30605\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__30634\,
            I => \N__30600\
        );

    \I__6590\ : Span4Mux_h
    port map (
            O => \N__30627\,
            I => \N__30600\
        );

    \I__6589\ : Odrv4
    port map (
            O => \N__30624\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__30619\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__6587\ : Odrv4
    port map (
            O => \N__30610\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__30605\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__6585\ : Odrv4
    port map (
            O => \N__30600\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__6584\ : InMux
    port map (
            O => \N__30589\,
            I => \N__30585\
        );

    \I__6583\ : InMux
    port map (
            O => \N__30588\,
            I => \N__30582\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__30585\,
            I => \N__30578\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__30582\,
            I => \N__30575\
        );

    \I__6580\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30572\
        );

    \I__6579\ : Span4Mux_v
    port map (
            O => \N__30578\,
            I => \N__30568\
        );

    \I__6578\ : Span4Mux_h
    port map (
            O => \N__30575\,
            I => \N__30562\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__30572\,
            I => \N__30562\
        );

    \I__6576\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30559\
        );

    \I__6575\ : Span4Mux_h
    port map (
            O => \N__30568\,
            I => \N__30556\
        );

    \I__6574\ : InMux
    port map (
            O => \N__30567\,
            I => \N__30553\
        );

    \I__6573\ : Span4Mux_v
    port map (
            O => \N__30562\,
            I => \N__30548\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__30559\,
            I => \N__30548\
        );

    \I__6571\ : Odrv4
    port map (
            O => \N__30556\,
            I => \N_1001_0\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__30553\,
            I => \N_1001_0\
        );

    \I__6569\ : Odrv4
    port map (
            O => \N__30548\,
            I => \N_1001_0\
        );

    \I__6568\ : InMux
    port map (
            O => \N__30541\,
            I => \N__30536\
        );

    \I__6567\ : InMux
    port map (
            O => \N__30540\,
            I => \N__30527\
        );

    \I__6566\ : InMux
    port map (
            O => \N__30539\,
            I => \N__30527\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__30536\,
            I => \N__30524\
        );

    \I__6564\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30521\
        );

    \I__6563\ : InMux
    port map (
            O => \N__30534\,
            I => \N__30517\
        );

    \I__6562\ : InMux
    port map (
            O => \N__30533\,
            I => \N__30514\
        );

    \I__6561\ : InMux
    port map (
            O => \N__30532\,
            I => \N__30511\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__30527\,
            I => \N__30508\
        );

    \I__6559\ : Span4Mux_v
    port map (
            O => \N__30524\,
            I => \N__30503\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__30521\,
            I => \N__30503\
        );

    \I__6557\ : InMux
    port map (
            O => \N__30520\,
            I => \N__30498\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__30517\,
            I => \N__30487\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__30514\,
            I => \N__30487\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__30511\,
            I => \N__30487\
        );

    \I__6553\ : Span4Mux_h
    port map (
            O => \N__30508\,
            I => \N__30487\
        );

    \I__6552\ : Span4Mux_h
    port map (
            O => \N__30503\,
            I => \N__30487\
        );

    \I__6551\ : InMux
    port map (
            O => \N__30502\,
            I => \N__30482\
        );

    \I__6550\ : InMux
    port map (
            O => \N__30501\,
            I => \N__30482\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__30498\,
            I => \N_814_0\
        );

    \I__6548\ : Odrv4
    port map (
            O => \N__30487\,
            I => \N_814_0\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__30482\,
            I => \N_814_0\
        );

    \I__6546\ : CascadeMux
    port map (
            O => \N__30475\,
            I => \N_1001_0_cascade_\
        );

    \I__6545\ : CascadeMux
    port map (
            O => \N__30472\,
            I => \N__30469\
        );

    \I__6544\ : InMux
    port map (
            O => \N__30469\,
            I => \N__30463\
        );

    \I__6543\ : InMux
    port map (
            O => \N__30468\,
            I => \N__30460\
        );

    \I__6542\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30448\
        );

    \I__6541\ : InMux
    port map (
            O => \N__30466\,
            I => \N__30445\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__30463\,
            I => \N__30442\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__30460\,
            I => \N__30439\
        );

    \I__6538\ : InMux
    port map (
            O => \N__30459\,
            I => \N__30436\
        );

    \I__6537\ : InMux
    port map (
            O => \N__30458\,
            I => \N__30433\
        );

    \I__6536\ : InMux
    port map (
            O => \N__30457\,
            I => \N__30430\
        );

    \I__6535\ : InMux
    port map (
            O => \N__30456\,
            I => \N__30425\
        );

    \I__6534\ : InMux
    port map (
            O => \N__30455\,
            I => \N__30422\
        );

    \I__6533\ : InMux
    port map (
            O => \N__30454\,
            I => \N__30415\
        );

    \I__6532\ : InMux
    port map (
            O => \N__30453\,
            I => \N__30415\
        );

    \I__6531\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30412\
        );

    \I__6530\ : CascadeMux
    port map (
            O => \N__30451\,
            I => \N__30409\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__30448\,
            I => \N__30406\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__30445\,
            I => \N__30403\
        );

    \I__6527\ : Span4Mux_h
    port map (
            O => \N__30442\,
            I => \N__30398\
        );

    \I__6526\ : Span4Mux_v
    port map (
            O => \N__30439\,
            I => \N__30398\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__30436\,
            I => \N__30393\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__30433\,
            I => \N__30393\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__30430\,
            I => \N__30390\
        );

    \I__6522\ : InMux
    port map (
            O => \N__30429\,
            I => \N__30385\
        );

    \I__6521\ : InMux
    port map (
            O => \N__30428\,
            I => \N__30385\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__30425\,
            I => \N__30380\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__30422\,
            I => \N__30380\
        );

    \I__6518\ : InMux
    port map (
            O => \N__30421\,
            I => \N__30377\
        );

    \I__6517\ : InMux
    port map (
            O => \N__30420\,
            I => \N__30374\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__30415\,
            I => \N__30371\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__30412\,
            I => \N__30368\
        );

    \I__6514\ : InMux
    port map (
            O => \N__30409\,
            I => \N__30365\
        );

    \I__6513\ : Span4Mux_v
    port map (
            O => \N__30406\,
            I => \N__30356\
        );

    \I__6512\ : Span4Mux_v
    port map (
            O => \N__30403\,
            I => \N__30356\
        );

    \I__6511\ : Span4Mux_h
    port map (
            O => \N__30398\,
            I => \N__30356\
        );

    \I__6510\ : Span4Mux_v
    port map (
            O => \N__30393\,
            I => \N__30356\
        );

    \I__6509\ : Span4Mux_v
    port map (
            O => \N__30390\,
            I => \N__30349\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__30385\,
            I => \N__30349\
        );

    \I__6507\ : Span4Mux_h
    port map (
            O => \N__30380\,
            I => \N__30349\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__30377\,
            I => \N__30346\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__30374\,
            I => \N__30343\
        );

    \I__6504\ : Odrv4
    port map (
            O => \N__30371\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__6503\ : Odrv12
    port map (
            O => \N__30368\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__30365\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__6501\ : Odrv4
    port map (
            O => \N__30356\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__6500\ : Odrv4
    port map (
            O => \N__30349\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__6499\ : Odrv12
    port map (
            O => \N__30346\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__6498\ : Odrv4
    port map (
            O => \N__30343\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__6497\ : InMux
    port map (
            O => \N__30328\,
            I => \N__30325\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__30325\,
            I => \N__30322\
        );

    \I__6495\ : Odrv12
    port map (
            O => \N__30322\,
            I => \this_vga_signals.g4\
        );

    \I__6494\ : CascadeMux
    port map (
            O => \N__30319\,
            I => \this_ppu.N_1278_cascade_\
        );

    \I__6493\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30310\
        );

    \I__6492\ : InMux
    port map (
            O => \N__30315\,
            I => \N__30310\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__30310\,
            I => \N__30307\
        );

    \I__6490\ : Span4Mux_h
    port map (
            O => \N__30307\,
            I => \N__30304\
        );

    \I__6489\ : Odrv4
    port map (
            O => \N__30304\,
            I => \this_ppu.N_767_0\
        );

    \I__6488\ : InMux
    port map (
            O => \N__30301\,
            I => \N__30298\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__30298\,
            I => \N__30293\
        );

    \I__6486\ : InMux
    port map (
            O => \N__30297\,
            I => \N__30288\
        );

    \I__6485\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30288\
        );

    \I__6484\ : Odrv4
    port map (
            O => \N__30293\,
            I => \this_ppu.N_1425\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__30288\,
            I => \this_ppu.N_1425\
        );

    \I__6482\ : CascadeMux
    port map (
            O => \N__30283\,
            I => \this_ppu.N_1149_cascade_\
        );

    \I__6481\ : CascadeMux
    port map (
            O => \N__30280\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_3_cascade_\
        );

    \I__6480\ : CascadeMux
    port map (
            O => \N__30277\,
            I => \this_vga_signals.g1_0_0_0_cascade_\
        );

    \I__6479\ : InMux
    port map (
            O => \N__30274\,
            I => \N__30271\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__30271\,
            I => \N__30268\
        );

    \I__6477\ : Span4Mux_v
    port map (
            O => \N__30268\,
            I => \N__30265\
        );

    \I__6476\ : Sp12to4
    port map (
            O => \N__30265\,
            I => \N__30262\
        );

    \I__6475\ : Odrv12
    port map (
            O => \N__30262\,
            I => \this_vga_signals.SUM_2_i_i_1_0_3\
        );

    \I__6474\ : InMux
    port map (
            O => \N__30259\,
            I => \N__30256\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__30256\,
            I => \N__30253\
        );

    \I__6472\ : Odrv4
    port map (
            O => \N__30253\,
            I => \this_vga_signals.N_5_0_0\
        );

    \I__6471\ : InMux
    port map (
            O => \N__30250\,
            I => \N__30247\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__30247\,
            I => \N__30244\
        );

    \I__6469\ : Odrv4
    port map (
            O => \N__30244\,
            I => \this_vga_signals.g1_0_1\
        );

    \I__6468\ : InMux
    port map (
            O => \N__30241\,
            I => \N__30235\
        );

    \I__6467\ : InMux
    port map (
            O => \N__30240\,
            I => \N__30235\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__30235\,
            I => \N__30232\
        );

    \I__6465\ : Odrv4
    port map (
            O => \N__30232\,
            I => \this_vga_signals.N_39_0_0\
        );

    \I__6464\ : CascadeMux
    port map (
            O => \N__30229\,
            I => \this_vga_signals.g1_3_0_0_cascade_\
        );

    \I__6463\ : InMux
    port map (
            O => \N__30226\,
            I => \N__30223\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__30223\,
            I => \this_vga_signals.N_4_1\
        );

    \I__6461\ : CascadeMux
    port map (
            O => \N__30220\,
            I => \this_vga_signals.g3_cascade_\
        );

    \I__6460\ : InMux
    port map (
            O => \N__30217\,
            I => \N__30214\
        );

    \I__6459\ : LocalMux
    port map (
            O => \N__30214\,
            I => \this_vga_signals.N_5_1\
        );

    \I__6458\ : InMux
    port map (
            O => \N__30211\,
            I => \N__30208\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__30208\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_0_0_1\
        );

    \I__6456\ : InMux
    port map (
            O => \N__30205\,
            I => \N__30202\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__30202\,
            I => \N__30199\
        );

    \I__6454\ : Odrv4
    port map (
            O => \N__30199\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__6453\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30193\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__30193\,
            I => \N__30190\
        );

    \I__6451\ : Odrv4
    port map (
            O => \N__30190\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_0_0_1\
        );

    \I__6450\ : InMux
    port map (
            O => \N__30187\,
            I => \N__30183\
        );

    \I__6449\ : CascadeMux
    port map (
            O => \N__30186\,
            I => \N__30180\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__30183\,
            I => \N__30177\
        );

    \I__6447\ : InMux
    port map (
            O => \N__30180\,
            I => \N__30174\
        );

    \I__6446\ : Span4Mux_v
    port map (
            O => \N__30177\,
            I => \N__30168\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__30174\,
            I => \N__30168\
        );

    \I__6444\ : InMux
    port map (
            O => \N__30173\,
            I => \N__30165\
        );

    \I__6443\ : Span4Mux_h
    port map (
            O => \N__30168\,
            I => \N__30162\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__30165\,
            I => \this_vga_signals.N_1264\
        );

    \I__6441\ : Odrv4
    port map (
            O => \N__30162\,
            I => \this_vga_signals.N_1264\
        );

    \I__6440\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30153\
        );

    \I__6439\ : InMux
    port map (
            O => \N__30156\,
            I => \N__30150\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__30153\,
            I => \N__30147\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__30150\,
            I => \N__30144\
        );

    \I__6436\ : Span4Mux_v
    port map (
            O => \N__30147\,
            I => \N__30141\
        );

    \I__6435\ : Span4Mux_h
    port map (
            O => \N__30144\,
            I => \N__30138\
        );

    \I__6434\ : Odrv4
    port map (
            O => \N__30141\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1\
        );

    \I__6433\ : Odrv4
    port map (
            O => \N__30138\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1\
        );

    \I__6432\ : CascadeMux
    port map (
            O => \N__30133\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_x1_cascade_\
        );

    \I__6431\ : InMux
    port map (
            O => \N__30130\,
            I => \N__30127\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__30127\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_x0\
        );

    \I__6429\ : InMux
    port map (
            O => \N__30124\,
            I => \N__30121\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__30121\,
            I => \N__30118\
        );

    \I__6427\ : Span4Mux_h
    port map (
            O => \N__30118\,
            I => \N__30115\
        );

    \I__6426\ : Odrv4
    port map (
            O => \N__30115\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_1\
        );

    \I__6425\ : InMux
    port map (
            O => \N__30112\,
            I => \N__30109\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__30109\,
            I => \N__30104\
        );

    \I__6423\ : InMux
    port map (
            O => \N__30108\,
            I => \N__30098\
        );

    \I__6422\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30098\
        );

    \I__6421\ : Span4Mux_v
    port map (
            O => \N__30104\,
            I => \N__30095\
        );

    \I__6420\ : InMux
    port map (
            O => \N__30103\,
            I => \N__30092\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__30098\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__6418\ : Odrv4
    port map (
            O => \N__30095\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__30092\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__6416\ : CascadeMux
    port map (
            O => \N__30085\,
            I => \this_vga_signals.mult1_un47_sum_c2_0_cascade_\
        );

    \I__6415\ : CascadeMux
    port map (
            O => \N__30082\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_\
        );

    \I__6414\ : InMux
    port map (
            O => \N__30079\,
            I => \N__30076\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__30076\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3\
        );

    \I__6412\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30069\
        );

    \I__6411\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30066\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__30069\,
            I => \N__30063\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__30066\,
            I => \N__30060\
        );

    \I__6408\ : Span4Mux_h
    port map (
            O => \N__30063\,
            I => \N__30057\
        );

    \I__6407\ : Odrv4
    port map (
            O => \N__30060\,
            I => \this_vga_signals.g1_0\
        );

    \I__6406\ : Odrv4
    port map (
            O => \N__30057\,
            I => \this_vga_signals.g1_0\
        );

    \I__6405\ : CascadeMux
    port map (
            O => \N__30052\,
            I => \N__30049\
        );

    \I__6404\ : InMux
    port map (
            O => \N__30049\,
            I => \N__30046\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__30046\,
            I => \N__30043\
        );

    \I__6402\ : Span4Mux_h
    port map (
            O => \N__30043\,
            I => \N__30040\
        );

    \I__6401\ : Odrv4
    port map (
            O => \N__30040\,
            I => \this_vga_signals.g0_0_1\
        );

    \I__6400\ : InMux
    port map (
            O => \N__30037\,
            I => \N__30034\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__30034\,
            I => \this_vga_signals.g0_3_0\
        );

    \I__6398\ : InMux
    port map (
            O => \N__30031\,
            I => \N__30025\
        );

    \I__6397\ : InMux
    port map (
            O => \N__30030\,
            I => \N__30020\
        );

    \I__6396\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30020\
        );

    \I__6395\ : InMux
    port map (
            O => \N__30028\,
            I => \N__30013\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__30025\,
            I => \N__30008\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__30020\,
            I => \N__30008\
        );

    \I__6392\ : InMux
    port map (
            O => \N__30019\,
            I => \N__30003\
        );

    \I__6391\ : InMux
    port map (
            O => \N__30018\,
            I => \N__30003\
        );

    \I__6390\ : InMux
    port map (
            O => \N__30017\,
            I => \N__29998\
        );

    \I__6389\ : InMux
    port map (
            O => \N__30016\,
            I => \N__29998\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__30013\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__6387\ : Odrv4
    port map (
            O => \N__30008\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__30003\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__29998\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__6384\ : InMux
    port map (
            O => \N__29989\,
            I => \N__29984\
        );

    \I__6383\ : CascadeMux
    port map (
            O => \N__29988\,
            I => \N__29975\
        );

    \I__6382\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29972\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__29984\,
            I => \N__29969\
        );

    \I__6380\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29964\
        );

    \I__6379\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29964\
        );

    \I__6378\ : InMux
    port map (
            O => \N__29981\,
            I => \N__29959\
        );

    \I__6377\ : InMux
    port map (
            O => \N__29980\,
            I => \N__29959\
        );

    \I__6376\ : InMux
    port map (
            O => \N__29979\,
            I => \N__29954\
        );

    \I__6375\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29954\
        );

    \I__6374\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29951\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__29972\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__6372\ : Odrv4
    port map (
            O => \N__29969\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__29964\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__29959\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__29954\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__29951\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__6367\ : InMux
    port map (
            O => \N__29938\,
            I => \N__29934\
        );

    \I__6366\ : CascadeMux
    port map (
            O => \N__29937\,
            I => \N__29931\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__29934\,
            I => \N__29926\
        );

    \I__6364\ : InMux
    port map (
            O => \N__29931\,
            I => \N__29923\
        );

    \I__6363\ : CascadeMux
    port map (
            O => \N__29930\,
            I => \N__29920\
        );

    \I__6362\ : InMux
    port map (
            O => \N__29929\,
            I => \N__29917\
        );

    \I__6361\ : Span4Mux_v
    port map (
            O => \N__29926\,
            I => \N__29912\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__29923\,
            I => \N__29912\
        );

    \I__6359\ : InMux
    port map (
            O => \N__29920\,
            I => \N__29909\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__29917\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__6357\ : Odrv4
    port map (
            O => \N__29912\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__29909\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__6355\ : CascadeMux
    port map (
            O => \N__29902\,
            I => \N__29899\
        );

    \I__6354\ : InMux
    port map (
            O => \N__29899\,
            I => \N__29896\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__29896\,
            I => \N__29893\
        );

    \I__6352\ : Span4Mux_h
    port map (
            O => \N__29893\,
            I => \N__29890\
        );

    \I__6351\ : Odrv4
    port map (
            O => \N__29890\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_4_1_0\
        );

    \I__6350\ : InMux
    port map (
            O => \N__29887\,
            I => \N__29881\
        );

    \I__6349\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29881\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__29881\,
            I => \N__29877\
        );

    \I__6347\ : InMux
    port map (
            O => \N__29880\,
            I => \N__29873\
        );

    \I__6346\ : Span4Mux_h
    port map (
            O => \N__29877\,
            I => \N__29869\
        );

    \I__6345\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29866\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__29873\,
            I => \N__29863\
        );

    \I__6343\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29860\
        );

    \I__6342\ : Odrv4
    port map (
            O => \N__29869\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__29866\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__6340\ : Odrv12
    port map (
            O => \N__29863\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__29860\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__6338\ : InMux
    port map (
            O => \N__29851\,
            I => \N__29844\
        );

    \I__6337\ : InMux
    port map (
            O => \N__29850\,
            I => \N__29844\
        );

    \I__6336\ : CascadeMux
    port map (
            O => \N__29849\,
            I => \N__29839\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__29844\,
            I => \N__29835\
        );

    \I__6334\ : InMux
    port map (
            O => \N__29843\,
            I => \N__29832\
        );

    \I__6333\ : InMux
    port map (
            O => \N__29842\,
            I => \N__29828\
        );

    \I__6332\ : InMux
    port map (
            O => \N__29839\,
            I => \N__29823\
        );

    \I__6331\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29823\
        );

    \I__6330\ : Span4Mux_v
    port map (
            O => \N__29835\,
            I => \N__29818\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__29832\,
            I => \N__29818\
        );

    \I__6328\ : InMux
    port map (
            O => \N__29831\,
            I => \N__29815\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__29828\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__29823\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__6325\ : Odrv4
    port map (
            O => \N__29818\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__29815\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__6323\ : CascadeMux
    port map (
            O => \N__29806\,
            I => \this_vga_signals.mult1_un47_sum_3_3_cascade_\
        );

    \I__6322\ : InMux
    port map (
            O => \N__29803\,
            I => \N__29800\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__29800\,
            I => \N__29797\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__29797\,
            I => \N__29794\
        );

    \I__6319\ : Odrv4
    port map (
            O => \N__29794\,
            I => \this_vga_signals.mult1_un54_sum_2_0_3\
        );

    \I__6318\ : InMux
    port map (
            O => \N__29791\,
            I => \N__29788\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__29788\,
            I => \N__29785\
        );

    \I__6316\ : Span12Mux_v
    port map (
            O => \N__29785\,
            I => \N__29782\
        );

    \I__6315\ : Span12Mux_h
    port map (
            O => \N__29782\,
            I => \N__29779\
        );

    \I__6314\ : Odrv12
    port map (
            O => \N__29779\,
            I => \this_ppu.m18_i_o2_0\
        );

    \I__6313\ : CascadeMux
    port map (
            O => \N__29776\,
            I => \N__29773\
        );

    \I__6312\ : InMux
    port map (
            O => \N__29773\,
            I => \N__29770\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__29770\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_0\
        );

    \I__6310\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29761\
        );

    \I__6309\ : CascadeMux
    port map (
            O => \N__29766\,
            I => \N__29757\
        );

    \I__6308\ : InMux
    port map (
            O => \N__29765\,
            I => \N__29750\
        );

    \I__6307\ : InMux
    port map (
            O => \N__29764\,
            I => \N__29747\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__29761\,
            I => \N__29744\
        );

    \I__6305\ : InMux
    port map (
            O => \N__29760\,
            I => \N__29737\
        );

    \I__6304\ : InMux
    port map (
            O => \N__29757\,
            I => \N__29737\
        );

    \I__6303\ : InMux
    port map (
            O => \N__29756\,
            I => \N__29737\
        );

    \I__6302\ : InMux
    port map (
            O => \N__29755\,
            I => \N__29730\
        );

    \I__6301\ : InMux
    port map (
            O => \N__29754\,
            I => \N__29730\
        );

    \I__6300\ : InMux
    port map (
            O => \N__29753\,
            I => \N__29730\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__29750\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__29747\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__6297\ : Odrv4
    port map (
            O => \N__29744\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__29737\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__29730\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__6294\ : InMux
    port map (
            O => \N__29719\,
            I => \N__29711\
        );

    \I__6293\ : CascadeMux
    port map (
            O => \N__29718\,
            I => \N__29708\
        );

    \I__6292\ : InMux
    port map (
            O => \N__29717\,
            I => \N__29698\
        );

    \I__6291\ : InMux
    port map (
            O => \N__29716\,
            I => \N__29698\
        );

    \I__6290\ : InMux
    port map (
            O => \N__29715\,
            I => \N__29693\
        );

    \I__6289\ : InMux
    port map (
            O => \N__29714\,
            I => \N__29693\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__29711\,
            I => \N__29690\
        );

    \I__6287\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29683\
        );

    \I__6286\ : InMux
    port map (
            O => \N__29707\,
            I => \N__29683\
        );

    \I__6285\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29683\
        );

    \I__6284\ : InMux
    port map (
            O => \N__29705\,
            I => \N__29676\
        );

    \I__6283\ : InMux
    port map (
            O => \N__29704\,
            I => \N__29676\
        );

    \I__6282\ : InMux
    port map (
            O => \N__29703\,
            I => \N__29676\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__29698\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__29693\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__29690\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__29683\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__29676\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__6276\ : InMux
    port map (
            O => \N__29665\,
            I => \N__29662\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__29662\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_3_0_0\
        );

    \I__6274\ : InMux
    port map (
            O => \N__29659\,
            I => \N__29655\
        );

    \I__6273\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29652\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__29655\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__29652\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0\
        );

    \I__6270\ : CascadeMux
    port map (
            O => \N__29647\,
            I => \N_814_0_cascade_\
        );

    \I__6269\ : CascadeMux
    port map (
            O => \N__29644\,
            I => \N__29639\
        );

    \I__6268\ : CascadeMux
    port map (
            O => \N__29643\,
            I => \N__29636\
        );

    \I__6267\ : InMux
    port map (
            O => \N__29642\,
            I => \N__29632\
        );

    \I__6266\ : InMux
    port map (
            O => \N__29639\,
            I => \N__29627\
        );

    \I__6265\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29627\
        );

    \I__6264\ : InMux
    port map (
            O => \N__29635\,
            I => \N__29623\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__29632\,
            I => \N__29613\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__29627\,
            I => \N__29613\
        );

    \I__6261\ : InMux
    port map (
            O => \N__29626\,
            I => \N__29610\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__29623\,
            I => \N__29607\
        );

    \I__6259\ : InMux
    port map (
            O => \N__29622\,
            I => \N__29602\
        );

    \I__6258\ : InMux
    port map (
            O => \N__29621\,
            I => \N__29602\
        );

    \I__6257\ : InMux
    port map (
            O => \N__29620\,
            I => \N__29599\
        );

    \I__6256\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29594\
        );

    \I__6255\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29594\
        );

    \I__6254\ : Span4Mux_h
    port map (
            O => \N__29613\,
            I => \N__29591\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__29610\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__6252\ : Odrv12
    port map (
            O => \N__29607\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__29602\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__29599\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__29594\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__6248\ : Odrv4
    port map (
            O => \N__29591\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__6247\ : CascadeMux
    port map (
            O => \N__29578\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_2_1_cascade_\
        );

    \I__6246\ : CascadeMux
    port map (
            O => \N__29575\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_2_2_cascade_\
        );

    \I__6245\ : InMux
    port map (
            O => \N__29572\,
            I => \N__29566\
        );

    \I__6244\ : InMux
    port map (
            O => \N__29571\,
            I => \N__29559\
        );

    \I__6243\ : InMux
    port map (
            O => \N__29570\,
            I => \N__29559\
        );

    \I__6242\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29559\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__29566\,
            I => \N__29554\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__29559\,
            I => \N__29551\
        );

    \I__6239\ : InMux
    port map (
            O => \N__29558\,
            I => \N__29546\
        );

    \I__6238\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29546\
        );

    \I__6237\ : Span4Mux_v
    port map (
            O => \N__29554\,
            I => \N__29539\
        );

    \I__6236\ : Span4Mux_v
    port map (
            O => \N__29551\,
            I => \N__29539\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__29546\,
            I => \N__29539\
        );

    \I__6234\ : Odrv4
    port map (
            O => \N__29539\,
            I => \this_vga_signals.mult1_un47_sum_c3_0\
        );

    \I__6233\ : InMux
    port map (
            O => \N__29536\,
            I => \N__29533\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__29533\,
            I => \N__29528\
        );

    \I__6231\ : CascadeMux
    port map (
            O => \N__29532\,
            I => \N__29524\
        );

    \I__6230\ : InMux
    port map (
            O => \N__29531\,
            I => \N__29519\
        );

    \I__6229\ : Span4Mux_h
    port map (
            O => \N__29528\,
            I => \N__29516\
        );

    \I__6228\ : InMux
    port map (
            O => \N__29527\,
            I => \N__29509\
        );

    \I__6227\ : InMux
    port map (
            O => \N__29524\,
            I => \N__29509\
        );

    \I__6226\ : InMux
    port map (
            O => \N__29523\,
            I => \N__29509\
        );

    \I__6225\ : InMux
    port map (
            O => \N__29522\,
            I => \N__29506\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__29519\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_2_2\
        );

    \I__6223\ : Odrv4
    port map (
            O => \N__29516\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_2_2\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__29509\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_2_2\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__29506\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_2_2\
        );

    \I__6220\ : CascadeMux
    port map (
            O => \N__29497\,
            I => \N__29494\
        );

    \I__6219\ : InMux
    port map (
            O => \N__29494\,
            I => \N__29491\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__29491\,
            I => \N__29485\
        );

    \I__6217\ : CascadeMux
    port map (
            O => \N__29490\,
            I => \N__29482\
        );

    \I__6216\ : CascadeMux
    port map (
            O => \N__29489\,
            I => \N__29477\
        );

    \I__6215\ : InMux
    port map (
            O => \N__29488\,
            I => \N__29473\
        );

    \I__6214\ : Span4Mux_h
    port map (
            O => \N__29485\,
            I => \N__29470\
        );

    \I__6213\ : InMux
    port map (
            O => \N__29482\,
            I => \N__29463\
        );

    \I__6212\ : InMux
    port map (
            O => \N__29481\,
            I => \N__29463\
        );

    \I__6211\ : InMux
    port map (
            O => \N__29480\,
            I => \N__29463\
        );

    \I__6210\ : InMux
    port map (
            O => \N__29477\,
            I => \N__29458\
        );

    \I__6209\ : InMux
    port map (
            O => \N__29476\,
            I => \N__29458\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__29473\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_2_0\
        );

    \I__6207\ : Odrv4
    port map (
            O => \N__29470\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_2_0\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__29463\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_2_0\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__29458\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_2_0\
        );

    \I__6204\ : CascadeMux
    port map (
            O => \N__29449\,
            I => \N__29446\
        );

    \I__6203\ : InMux
    port map (
            O => \N__29446\,
            I => \N__29442\
        );

    \I__6202\ : CascadeMux
    port map (
            O => \N__29445\,
            I => \N__29439\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__29442\,
            I => \N__29436\
        );

    \I__6200\ : InMux
    port map (
            O => \N__29439\,
            I => \N__29433\
        );

    \I__6199\ : Odrv4
    port map (
            O => \N__29436\,
            I => \this_ppu.N_1341\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__29433\,
            I => \this_ppu.N_1341\
        );

    \I__6197\ : InMux
    port map (
            O => \N__29428\,
            I => \N__29424\
        );

    \I__6196\ : InMux
    port map (
            O => \N__29427\,
            I => \N__29419\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__29424\,
            I => \N__29415\
        );

    \I__6194\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29412\
        );

    \I__6193\ : InMux
    port map (
            O => \N__29422\,
            I => \N__29408\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__29419\,
            I => \N__29404\
        );

    \I__6191\ : InMux
    port map (
            O => \N__29418\,
            I => \N__29401\
        );

    \I__6190\ : Span4Mux_v
    port map (
            O => \N__29415\,
            I => \N__29396\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__29412\,
            I => \N__29396\
        );

    \I__6188\ : InMux
    port map (
            O => \N__29411\,
            I => \N__29393\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__29408\,
            I => \N__29390\
        );

    \I__6186\ : InMux
    port map (
            O => \N__29407\,
            I => \N__29387\
        );

    \I__6185\ : Span4Mux_h
    port map (
            O => \N__29404\,
            I => \N__29384\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__29401\,
            I => \N__29381\
        );

    \I__6183\ : Span4Mux_v
    port map (
            O => \N__29396\,
            I => \N__29376\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__29393\,
            I => \N__29376\
        );

    \I__6181\ : Span12Mux_s4_v
    port map (
            O => \N__29390\,
            I => \N__29370\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__29387\,
            I => \N__29370\
        );

    \I__6179\ : Span4Mux_v
    port map (
            O => \N__29384\,
            I => \N__29365\
        );

    \I__6178\ : Span4Mux_h
    port map (
            O => \N__29381\,
            I => \N__29365\
        );

    \I__6177\ : Sp12to4
    port map (
            O => \N__29376\,
            I => \N__29362\
        );

    \I__6176\ : InMux
    port map (
            O => \N__29375\,
            I => \N__29359\
        );

    \I__6175\ : Span12Mux_h
    port map (
            O => \N__29370\,
            I => \N__29356\
        );

    \I__6174\ : Span4Mux_h
    port map (
            O => \N__29365\,
            I => \N__29353\
        );

    \I__6173\ : Span12Mux_v
    port map (
            O => \N__29362\,
            I => \N__29348\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__29359\,
            I => \N__29348\
        );

    \I__6171\ : Odrv12
    port map (
            O => \N__29356\,
            I => \M_this_spr_ram_write_data_2\
        );

    \I__6170\ : Odrv4
    port map (
            O => \N__29353\,
            I => \M_this_spr_ram_write_data_2\
        );

    \I__6169\ : Odrv12
    port map (
            O => \N__29348\,
            I => \M_this_spr_ram_write_data_2\
        );

    \I__6168\ : InMux
    port map (
            O => \N__29341\,
            I => \N__29338\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__29338\,
            I => \N__29335\
        );

    \I__6166\ : Span4Mux_h
    port map (
            O => \N__29335\,
            I => \N__29332\
        );

    \I__6165\ : Span4Mux_h
    port map (
            O => \N__29332\,
            I => \N__29329\
        );

    \I__6164\ : Span4Mux_h
    port map (
            O => \N__29329\,
            I => \N__29326\
        );

    \I__6163\ : Span4Mux_h
    port map (
            O => \N__29326\,
            I => \N__29323\
        );

    \I__6162\ : Odrv4
    port map (
            O => \N__29323\,
            I => \this_ppu.oam_cache.mem_5\
        );

    \I__6161\ : InMux
    port map (
            O => \N__29320\,
            I => \N__29317\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__29317\,
            I => \N__29314\
        );

    \I__6159\ : Span4Mux_h
    port map (
            O => \N__29314\,
            I => \N__29311\
        );

    \I__6158\ : Odrv4
    port map (
            O => \N__29311\,
            I => \this_vga_signals.mult1_un54_sum_1_3\
        );

    \I__6157\ : CascadeMux
    port map (
            O => \N__29308\,
            I => \this_vga_signals.mult1_un47_sum_0_3_cascade_\
        );

    \I__6156\ : InMux
    port map (
            O => \N__29305\,
            I => \N__29302\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__29302\,
            I => \this_vga_signals.N_7\
        );

    \I__6154\ : CascadeMux
    port map (
            O => \N__29299\,
            I => \N__29296\
        );

    \I__6153\ : InMux
    port map (
            O => \N__29296\,
            I => \N__29293\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__29293\,
            I => \this_vga_signals.mult1_un47_sum_2_3\
        );

    \I__6151\ : InMux
    port map (
            O => \N__29290\,
            I => \N__29286\
        );

    \I__6150\ : InMux
    port map (
            O => \N__29289\,
            I => \N__29282\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__29286\,
            I => \N__29278\
        );

    \I__6148\ : InMux
    port map (
            O => \N__29285\,
            I => \N__29275\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__29282\,
            I => \N__29272\
        );

    \I__6146\ : InMux
    port map (
            O => \N__29281\,
            I => \N__29268\
        );

    \I__6145\ : Span12Mux_v
    port map (
            O => \N__29278\,
            I => \N__29263\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__29275\,
            I => \N__29263\
        );

    \I__6143\ : Span4Mux_v
    port map (
            O => \N__29272\,
            I => \N__29260\
        );

    \I__6142\ : InMux
    port map (
            O => \N__29271\,
            I => \N__29257\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__29268\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__6140\ : Odrv12
    port map (
            O => \N__29263\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__6139\ : Odrv4
    port map (
            O => \N__29260\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__29257\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__6137\ : InMux
    port map (
            O => \N__29248\,
            I => \N__29245\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__29245\,
            I => \N__29241\
        );

    \I__6135\ : CascadeMux
    port map (
            O => \N__29244\,
            I => \N__29237\
        );

    \I__6134\ : Span4Mux_v
    port map (
            O => \N__29241\,
            I => \N__29234\
        );

    \I__6133\ : InMux
    port map (
            O => \N__29240\,
            I => \N__29231\
        );

    \I__6132\ : InMux
    port map (
            O => \N__29237\,
            I => \N__29228\
        );

    \I__6131\ : Span4Mux_h
    port map (
            O => \N__29234\,
            I => \N__29223\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__29231\,
            I => \N__29223\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__29228\,
            I => \N__29216\
        );

    \I__6128\ : Span4Mux_h
    port map (
            O => \N__29223\,
            I => \N__29216\
        );

    \I__6127\ : InMux
    port map (
            O => \N__29222\,
            I => \N__29211\
        );

    \I__6126\ : InMux
    port map (
            O => \N__29221\,
            I => \N__29211\
        );

    \I__6125\ : Odrv4
    port map (
            O => \N__29216\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__29211\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__6123\ : CascadeMux
    port map (
            O => \N__29206\,
            I => \N__29202\
        );

    \I__6122\ : InMux
    port map (
            O => \N__29205\,
            I => \N__29198\
        );

    \I__6121\ : InMux
    port map (
            O => \N__29202\,
            I => \N__29195\
        );

    \I__6120\ : InMux
    port map (
            O => \N__29201\,
            I => \N__29191\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__29198\,
            I => \N__29185\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__29195\,
            I => \N__29185\
        );

    \I__6117\ : InMux
    port map (
            O => \N__29194\,
            I => \N__29182\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__29191\,
            I => \N__29179\
        );

    \I__6115\ : InMux
    port map (
            O => \N__29190\,
            I => \N__29176\
        );

    \I__6114\ : Span4Mux_v
    port map (
            O => \N__29185\,
            I => \N__29171\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__29182\,
            I => \N__29171\
        );

    \I__6112\ : Span4Mux_h
    port map (
            O => \N__29179\,
            I => \N__29168\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__29176\,
            I => \this_ppu.N_1301\
        );

    \I__6110\ : Odrv4
    port map (
            O => \N__29171\,
            I => \this_ppu.N_1301\
        );

    \I__6109\ : Odrv4
    port map (
            O => \N__29168\,
            I => \this_ppu.N_1301\
        );

    \I__6108\ : InMux
    port map (
            O => \N__29161\,
            I => \N__29158\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__29158\,
            I => \this_ppu.M_this_state_q_srsts_i_i_0_0Z0Z_15\
        );

    \I__6106\ : CascadeMux
    port map (
            O => \N__29155\,
            I => \N__29152\
        );

    \I__6105\ : InMux
    port map (
            O => \N__29152\,
            I => \N__29148\
        );

    \I__6104\ : CascadeMux
    port map (
            O => \N__29151\,
            I => \N__29145\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__29148\,
            I => \N__29139\
        );

    \I__6102\ : InMux
    port map (
            O => \N__29145\,
            I => \N__29136\
        );

    \I__6101\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29133\
        );

    \I__6100\ : InMux
    port map (
            O => \N__29143\,
            I => \N__29128\
        );

    \I__6099\ : InMux
    port map (
            O => \N__29142\,
            I => \N__29128\
        );

    \I__6098\ : Span4Mux_v
    port map (
            O => \N__29139\,
            I => \N__29121\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__29136\,
            I => \N__29121\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__29133\,
            I => \N__29121\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__29128\,
            I => \M_this_state_qZ0Z_15\
        );

    \I__6094\ : Odrv4
    port map (
            O => \N__29121\,
            I => \M_this_state_qZ0Z_15\
        );

    \I__6093\ : CascadeMux
    port map (
            O => \N__29116\,
            I => \N__29113\
        );

    \I__6092\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29110\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__29110\,
            I => \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_7\
        );

    \I__6090\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29104\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__29104\,
            I => \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_11\
        );

    \I__6088\ : CascadeMux
    port map (
            O => \N__29101\,
            I => \N__29098\
        );

    \I__6087\ : InMux
    port map (
            O => \N__29098\,
            I => \N__29095\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__29095\,
            I => \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_8\
        );

    \I__6085\ : CascadeMux
    port map (
            O => \N__29092\,
            I => \this_ppu.N_807_0_cascade_\
        );

    \I__6084\ : InMux
    port map (
            O => \N__29089\,
            I => \N__29086\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__29086\,
            I => \N__29083\
        );

    \I__6082\ : Span4Mux_v
    port map (
            O => \N__29083\,
            I => \N__29077\
        );

    \I__6081\ : InMux
    port map (
            O => \N__29082\,
            I => \N__29074\
        );

    \I__6080\ : InMux
    port map (
            O => \N__29081\,
            I => \N__29069\
        );

    \I__6079\ : InMux
    port map (
            O => \N__29080\,
            I => \N__29069\
        );

    \I__6078\ : Odrv4
    port map (
            O => \N__29077\,
            I => \this_ppu.N_1002_0\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__29074\,
            I => \this_ppu.N_1002_0\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__29069\,
            I => \this_ppu.N_1002_0\
        );

    \I__6075\ : InMux
    port map (
            O => \N__29062\,
            I => \N__29059\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__29059\,
            I => \this_ppu.N_235_2_0\
        );

    \I__6073\ : CascadeMux
    port map (
            O => \N__29056\,
            I => \this_ppu.N_235_2_0_cascade_\
        );

    \I__6072\ : InMux
    port map (
            O => \N__29053\,
            I => \N__29047\
        );

    \I__6071\ : InMux
    port map (
            O => \N__29052\,
            I => \N__29047\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__29047\,
            I => \N__29043\
        );

    \I__6069\ : InMux
    port map (
            O => \N__29046\,
            I => \N__29038\
        );

    \I__6068\ : Span4Mux_h
    port map (
            O => \N__29043\,
            I => \N__29035\
        );

    \I__6067\ : InMux
    port map (
            O => \N__29042\,
            I => \N__29032\
        );

    \I__6066\ : InMux
    port map (
            O => \N__29041\,
            I => \N__29029\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__29038\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__6064\ : Odrv4
    port map (
            O => \N__29035\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__29032\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__29029\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__6061\ : InMux
    port map (
            O => \N__29020\,
            I => \N__29017\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__29017\,
            I => \this_ppu.N_1162\
        );

    \I__6059\ : InMux
    port map (
            O => \N__29014\,
            I => \N__29011\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__29011\,
            I => \this_vga_signals.g0_5\
        );

    \I__6057\ : CascadeMux
    port map (
            O => \N__29008\,
            I => \N__29004\
        );

    \I__6056\ : InMux
    port map (
            O => \N__29007\,
            I => \N__28999\
        );

    \I__6055\ : InMux
    port map (
            O => \N__29004\,
            I => \N__28992\
        );

    \I__6054\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28992\
        );

    \I__6053\ : InMux
    port map (
            O => \N__29002\,
            I => \N__28992\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__28999\,
            I => \this_vga_signals.mult1_un61_sum_axb1_0\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__28992\,
            I => \this_vga_signals.mult1_un61_sum_axb1_0\
        );

    \I__6050\ : CascadeMux
    port map (
            O => \N__28987\,
            I => \N__28983\
        );

    \I__6049\ : CascadeMux
    port map (
            O => \N__28986\,
            I => \N__28978\
        );

    \I__6048\ : InMux
    port map (
            O => \N__28983\,
            I => \N__28972\
        );

    \I__6047\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28972\
        );

    \I__6046\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28969\
        );

    \I__6045\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28964\
        );

    \I__6044\ : InMux
    port map (
            O => \N__28977\,
            I => \N__28964\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__28972\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__28969\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__28964\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__6040\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28954\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__28954\,
            I => \N__28951\
        );

    \I__6038\ : Odrv4
    port map (
            O => \N__28951\,
            I => \this_vga_signals.g0_1_0\
        );

    \I__6037\ : InMux
    port map (
            O => \N__28948\,
            I => \N__28944\
        );

    \I__6036\ : CascadeMux
    port map (
            O => \N__28947\,
            I => \N__28941\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__28944\,
            I => \N__28938\
        );

    \I__6034\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28932\
        );

    \I__6033\ : Span4Mux_h
    port map (
            O => \N__28938\,
            I => \N__28925\
        );

    \I__6032\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28918\
        );

    \I__6031\ : InMux
    port map (
            O => \N__28936\,
            I => \N__28918\
        );

    \I__6030\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28918\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__28932\,
            I => \N__28915\
        );

    \I__6028\ : InMux
    port map (
            O => \N__28931\,
            I => \N__28910\
        );

    \I__6027\ : InMux
    port map (
            O => \N__28930\,
            I => \N__28910\
        );

    \I__6026\ : CascadeMux
    port map (
            O => \N__28929\,
            I => \N__28906\
        );

    \I__6025\ : InMux
    port map (
            O => \N__28928\,
            I => \N__28900\
        );

    \I__6024\ : Span4Mux_h
    port map (
            O => \N__28925\,
            I => \N__28897\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__28918\,
            I => \N__28894\
        );

    \I__6022\ : Span4Mux_v
    port map (
            O => \N__28915\,
            I => \N__28891\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__28910\,
            I => \N__28888\
        );

    \I__6020\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28885\
        );

    \I__6019\ : InMux
    port map (
            O => \N__28906\,
            I => \N__28880\
        );

    \I__6018\ : InMux
    port map (
            O => \N__28905\,
            I => \N__28880\
        );

    \I__6017\ : InMux
    port map (
            O => \N__28904\,
            I => \N__28875\
        );

    \I__6016\ : InMux
    port map (
            O => \N__28903\,
            I => \N__28875\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__28900\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__6014\ : Odrv4
    port map (
            O => \N__28897\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__6013\ : Odrv4
    port map (
            O => \N__28894\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__6012\ : Odrv4
    port map (
            O => \N__28891\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__6011\ : Odrv4
    port map (
            O => \N__28888\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__28885\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__28880\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__28875\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__6007\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28852\
        );

    \I__6006\ : InMux
    port map (
            O => \N__28857\,
            I => \N__28849\
        );

    \I__6005\ : InMux
    port map (
            O => \N__28856\,
            I => \N__28844\
        );

    \I__6004\ : InMux
    port map (
            O => \N__28855\,
            I => \N__28844\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__28852\,
            I => \this_vga_signals.mult1_un61_sum_c3_0\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__28849\,
            I => \this_vga_signals.mult1_un61_sum_c3_0\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__28844\,
            I => \this_vga_signals.mult1_un61_sum_c3_0\
        );

    \I__6000\ : CascadeMux
    port map (
            O => \N__28837\,
            I => \this_vga_signals.mult1_un68_sum_c2_0_cascade_\
        );

    \I__5999\ : InMux
    port map (
            O => \N__28834\,
            I => \N__28831\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__28831\,
            I => \this_vga_signals.g0_0_3_1\
        );

    \I__5997\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28825\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__28825\,
            I => \this_vga_signals.g0_0_3\
        );

    \I__5995\ : InMux
    port map (
            O => \N__28822\,
            I => \N__28819\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__28819\,
            I => \N__28816\
        );

    \I__5993\ : Odrv4
    port map (
            O => \N__28816\,
            I => \this_vga_signals.g1_1\
        );

    \I__5992\ : CascadeMux
    port map (
            O => \N__28813\,
            I => \N__28810\
        );

    \I__5991\ : InMux
    port map (
            O => \N__28810\,
            I => \N__28807\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__28807\,
            I => \N__28804\
        );

    \I__5989\ : Span4Mux_v
    port map (
            O => \N__28804\,
            I => \N__28801\
        );

    \I__5988\ : Odrv4
    port map (
            O => \N__28801\,
            I => \this_vga_signals.mult1_un54_sum_0_1\
        );

    \I__5987\ : InMux
    port map (
            O => \N__28798\,
            I => \N__28795\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__28795\,
            I => \this_vga_signals.g0_2_0\
        );

    \I__5985\ : InMux
    port map (
            O => \N__28792\,
            I => \N__28789\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__28789\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_0\
        );

    \I__5983\ : InMux
    port map (
            O => \N__28786\,
            I => \N__28781\
        );

    \I__5982\ : InMux
    port map (
            O => \N__28785\,
            I => \N__28776\
        );

    \I__5981\ : InMux
    port map (
            O => \N__28784\,
            I => \N__28776\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__28781\,
            I => \this_vga_signals.vaddress_9\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__28776\,
            I => \this_vga_signals.vaddress_9\
        );

    \I__5978\ : InMux
    port map (
            O => \N__28771\,
            I => \N__28761\
        );

    \I__5977\ : InMux
    port map (
            O => \N__28770\,
            I => \N__28761\
        );

    \I__5976\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28758\
        );

    \I__5975\ : InMux
    port map (
            O => \N__28768\,
            I => \N__28755\
        );

    \I__5974\ : InMux
    port map (
            O => \N__28767\,
            I => \N__28750\
        );

    \I__5973\ : InMux
    port map (
            O => \N__28766\,
            I => \N__28750\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__28761\,
            I => \N__28745\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__28758\,
            I => \N__28742\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__28755\,
            I => \N__28737\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__28750\,
            I => \N__28737\
        );

    \I__5968\ : InMux
    port map (
            O => \N__28749\,
            I => \N__28732\
        );

    \I__5967\ : InMux
    port map (
            O => \N__28748\,
            I => \N__28732\
        );

    \I__5966\ : Span4Mux_v
    port map (
            O => \N__28745\,
            I => \N__28729\
        );

    \I__5965\ : Span4Mux_h
    port map (
            O => \N__28742\,
            I => \N__28726\
        );

    \I__5964\ : Odrv12
    port map (
            O => \N__28737\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_1\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__28732\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_1\
        );

    \I__5962\ : Odrv4
    port map (
            O => \N__28729\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_1\
        );

    \I__5961\ : Odrv4
    port map (
            O => \N__28726\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_1\
        );

    \I__5960\ : CascadeMux
    port map (
            O => \N__28717\,
            I => \N__28714\
        );

    \I__5959\ : InMux
    port map (
            O => \N__28714\,
            I => \N__28706\
        );

    \I__5958\ : InMux
    port map (
            O => \N__28713\,
            I => \N__28706\
        );

    \I__5957\ : InMux
    port map (
            O => \N__28712\,
            I => \N__28697\
        );

    \I__5956\ : InMux
    port map (
            O => \N__28711\,
            I => \N__28697\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__28706\,
            I => \N__28694\
        );

    \I__5954\ : InMux
    port map (
            O => \N__28705\,
            I => \N__28690\
        );

    \I__5953\ : InMux
    port map (
            O => \N__28704\,
            I => \N__28683\
        );

    \I__5952\ : InMux
    port map (
            O => \N__28703\,
            I => \N__28683\
        );

    \I__5951\ : InMux
    port map (
            O => \N__28702\,
            I => \N__28683\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__28697\,
            I => \N__28678\
        );

    \I__5949\ : Span4Mux_h
    port map (
            O => \N__28694\,
            I => \N__28678\
        );

    \I__5948\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28675\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__28690\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__28683\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__5945\ : Odrv4
    port map (
            O => \N__28678\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__28675\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__5943\ : InMux
    port map (
            O => \N__28666\,
            I => \N__28661\
        );

    \I__5942\ : InMux
    port map (
            O => \N__28665\,
            I => \N__28658\
        );

    \I__5941\ : InMux
    port map (
            O => \N__28664\,
            I => \N__28655\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__28661\,
            I => \N__28652\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__28658\,
            I => \N__28645\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__28655\,
            I => \N__28642\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__28652\,
            I => \N__28639\
        );

    \I__5936\ : InMux
    port map (
            O => \N__28651\,
            I => \N__28634\
        );

    \I__5935\ : InMux
    port map (
            O => \N__28650\,
            I => \N__28634\
        );

    \I__5934\ : InMux
    port map (
            O => \N__28649\,
            I => \N__28629\
        );

    \I__5933\ : InMux
    port map (
            O => \N__28648\,
            I => \N__28629\
        );

    \I__5932\ : Odrv4
    port map (
            O => \N__28645\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__5931\ : Odrv12
    port map (
            O => \N__28642\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__5930\ : Odrv4
    port map (
            O => \N__28639\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__28634\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__28629\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__5927\ : CascadeMux
    port map (
            O => \N__28618\,
            I => \N__28615\
        );

    \I__5926\ : InMux
    port map (
            O => \N__28615\,
            I => \N__28612\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__28612\,
            I => \N__28609\
        );

    \I__5924\ : Span4Mux_h
    port map (
            O => \N__28609\,
            I => \N__28606\
        );

    \I__5923\ : Odrv4
    port map (
            O => \N__28606\,
            I => \this_vga_signals.g0_0_x2\
        );

    \I__5922\ : InMux
    port map (
            O => \N__28603\,
            I => \N__28600\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__28600\,
            I => \this_vga_signals.if_m5_i_0_0_0\
        );

    \I__5920\ : InMux
    port map (
            O => \N__28597\,
            I => \N__28594\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__28594\,
            I => \this_vga_signals.mult1_un54_sum_c3_x0\
        );

    \I__5918\ : CascadeMux
    port map (
            O => \N__28591\,
            I => \this_vga_signals.if_N_7_0_cascade_\
        );

    \I__5917\ : InMux
    port map (
            O => \N__28588\,
            I => \N__28585\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__28585\,
            I => \N__28581\
        );

    \I__5915\ : InMux
    port map (
            O => \N__28584\,
            I => \N__28578\
        );

    \I__5914\ : Span4Mux_v
    port map (
            O => \N__28581\,
            I => \N__28575\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__28578\,
            I => \N__28572\
        );

    \I__5912\ : Span4Mux_v
    port map (
            O => \N__28575\,
            I => \N__28569\
        );

    \I__5911\ : Odrv12
    port map (
            O => \N__28572\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__5910\ : Odrv4
    port map (
            O => \N__28569\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__5909\ : CascadeMux
    port map (
            O => \N__28564\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_d_cascade_\
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__28561\,
            I => \N__28558\
        );

    \I__5907\ : InMux
    port map (
            O => \N__28558\,
            I => \N__28555\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__28555\,
            I => \N__28552\
        );

    \I__5905\ : Odrv4
    port map (
            O => \N__28552\,
            I => \this_vga_signals.mult1_un47_sum_1_3\
        );

    \I__5904\ : InMux
    port map (
            O => \N__28549\,
            I => \N__28546\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__28546\,
            I => \N__28543\
        );

    \I__5902\ : Odrv4
    port map (
            O => \N__28543\,
            I => \this_vga_signals.mult1_un54_sum_1_1\
        );

    \I__5901\ : InMux
    port map (
            O => \N__28540\,
            I => \N__28536\
        );

    \I__5900\ : InMux
    port map (
            O => \N__28539\,
            I => \N__28533\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__28536\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__28533\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c\
        );

    \I__5897\ : CascadeMux
    port map (
            O => \N__28528\,
            I => \this_vga_signals.mult1_un54_sum_0_3_cascade_\
        );

    \I__5896\ : InMux
    port map (
            O => \N__28525\,
            I => \N__28521\
        );

    \I__5895\ : InMux
    port map (
            O => \N__28524\,
            I => \N__28518\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__28521\,
            I => \N__28513\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__28518\,
            I => \N__28510\
        );

    \I__5892\ : InMux
    port map (
            O => \N__28517\,
            I => \N__28507\
        );

    \I__5891\ : InMux
    port map (
            O => \N__28516\,
            I => \N__28504\
        );

    \I__5890\ : Span4Mux_h
    port map (
            O => \N__28513\,
            I => \N__28501\
        );

    \I__5889\ : Odrv4
    port map (
            O => \N__28510\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_d\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__28507\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_d\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__28504\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_d\
        );

    \I__5886\ : Odrv4
    port map (
            O => \N__28501\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_d\
        );

    \I__5885\ : CascadeMux
    port map (
            O => \N__28492\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_1_cascade_\
        );

    \I__5884\ : InMux
    port map (
            O => \N__28489\,
            I => \N__28486\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__28486\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0\
        );

    \I__5882\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28480\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__28480\,
            I => \N__28477\
        );

    \I__5880\ : Odrv12
    port map (
            O => \N__28477\,
            I => \this_vga_signals.N_3_1_0_1\
        );

    \I__5879\ : CascadeMux
    port map (
            O => \N__28474\,
            I => \N__28471\
        );

    \I__5878\ : InMux
    port map (
            O => \N__28471\,
            I => \N__28468\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__28468\,
            I => \N__28465\
        );

    \I__5876\ : Span4Mux_h
    port map (
            O => \N__28465\,
            I => \N__28462\
        );

    \I__5875\ : Odrv4
    port map (
            O => \N__28462\,
            I => \this_vga_signals.g0_2_1\
        );

    \I__5874\ : CascadeMux
    port map (
            O => \N__28459\,
            I => \this_vga_signals.mult1_un54_sum_c2_0_cascade_\
        );

    \I__5873\ : InMux
    port map (
            O => \N__28456\,
            I => \N__28453\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__28453\,
            I => \N__28450\
        );

    \I__5871\ : Odrv4
    port map (
            O => \N__28450\,
            I => \this_vga_signals.g0_4\
        );

    \I__5870\ : CascadeMux
    port map (
            O => \N__28447\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\
        );

    \I__5869\ : InMux
    port map (
            O => \N__28444\,
            I => \N__28441\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__28441\,
            I => \this_vga_signals.mult1_un47_sum_4_3\
        );

    \I__5867\ : CascadeMux
    port map (
            O => \N__28438\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1_cascade_\
        );

    \I__5866\ : CascadeMux
    port map (
            O => \N__28435\,
            I => \N__28432\
        );

    \I__5865\ : InMux
    port map (
            O => \N__28432\,
            I => \N__28429\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__28429\,
            I => \this_vga_signals.mult1_un54_sum_c3_x1\
        );

    \I__5863\ : InMux
    port map (
            O => \N__28426\,
            I => \N__28420\
        );

    \I__5862\ : InMux
    port map (
            O => \N__28425\,
            I => \N__28417\
        );

    \I__5861\ : InMux
    port map (
            O => \N__28424\,
            I => \N__28414\
        );

    \I__5860\ : InMux
    port map (
            O => \N__28423\,
            I => \N__28411\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__28420\,
            I => \N__28408\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__28417\,
            I => \N__28403\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__28414\,
            I => \N__28403\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__28411\,
            I => \N__28400\
        );

    \I__5855\ : Span4Mux_h
    port map (
            O => \N__28408\,
            I => \N__28397\
        );

    \I__5854\ : Span4Mux_v
    port map (
            O => \N__28403\,
            I => \N__28392\
        );

    \I__5853\ : Span4Mux_h
    port map (
            O => \N__28400\,
            I => \N__28392\
        );

    \I__5852\ : Odrv4
    port map (
            O => \N__28397\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_3\
        );

    \I__5851\ : Odrv4
    port map (
            O => \N__28392\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_3\
        );

    \I__5850\ : InMux
    port map (
            O => \N__28387\,
            I => \N__28384\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__28384\,
            I => \N__28380\
        );

    \I__5848\ : InMux
    port map (
            O => \N__28383\,
            I => \N__28377\
        );

    \I__5847\ : Span4Mux_h
    port map (
            O => \N__28380\,
            I => \N__28374\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__28377\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1\
        );

    \I__5845\ : Odrv4
    port map (
            O => \N__28374\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1\
        );

    \I__5844\ : InMux
    port map (
            O => \N__28369\,
            I => \N__28366\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__28366\,
            I => \this_vga_signals.N_27_0\
        );

    \I__5842\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28360\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__28360\,
            I => \N__28356\
        );

    \I__5840\ : InMux
    port map (
            O => \N__28359\,
            I => \N__28353\
        );

    \I__5839\ : Span4Mux_v
    port map (
            O => \N__28356\,
            I => \N__28350\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__28353\,
            I => \N__28347\
        );

    \I__5837\ : Span4Mux_h
    port map (
            O => \N__28350\,
            I => \N__28344\
        );

    \I__5836\ : Span4Mux_v
    port map (
            O => \N__28347\,
            I => \N__28341\
        );

    \I__5835\ : Odrv4
    port map (
            O => \N__28344\,
            I => \this_vga_signals.N_1247\
        );

    \I__5834\ : Odrv4
    port map (
            O => \N__28341\,
            I => \this_vga_signals.N_1247\
        );

    \I__5833\ : CascadeMux
    port map (
            O => \N__28336\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0_cascade_\
        );

    \I__5832\ : InMux
    port map (
            O => \N__28333\,
            I => \N__28329\
        );

    \I__5831\ : InMux
    port map (
            O => \N__28332\,
            I => \N__28326\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__28329\,
            I => \N__28322\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__28326\,
            I => \N__28319\
        );

    \I__5828\ : InMux
    port map (
            O => \N__28325\,
            I => \N__28316\
        );

    \I__5827\ : Span12Mux_v
    port map (
            O => \N__28322\,
            I => \N__28313\
        );

    \I__5826\ : Span4Mux_v
    port map (
            O => \N__28319\,
            I => \N__28310\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__28316\,
            I => \N__28307\
        );

    \I__5824\ : Odrv12
    port map (
            O => \N__28313\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__28310\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__5822\ : Odrv12
    port map (
            O => \N__28307\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__5821\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28297\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__28297\,
            I => \N__28294\
        );

    \I__5819\ : Span4Mux_v
    port map (
            O => \N__28294\,
            I => \N__28289\
        );

    \I__5818\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28286\
        );

    \I__5817\ : InMux
    port map (
            O => \N__28292\,
            I => \N__28283\
        );

    \I__5816\ : Span4Mux_v
    port map (
            O => \N__28289\,
            I => \N__28280\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__28286\,
            I => \N__28275\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__28283\,
            I => \N__28275\
        );

    \I__5813\ : Odrv4
    port map (
            O => \N__28280\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\
        );

    \I__5812\ : Odrv12
    port map (
            O => \N__28275\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\
        );

    \I__5811\ : InMux
    port map (
            O => \N__28270\,
            I => \N__28264\
        );

    \I__5810\ : InMux
    port map (
            O => \N__28269\,
            I => \N__28264\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__28264\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__5808\ : InMux
    port map (
            O => \N__28261\,
            I => \N__28257\
        );

    \I__5807\ : CascadeMux
    port map (
            O => \N__28260\,
            I => \N__28254\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__28257\,
            I => \N__28250\
        );

    \I__5805\ : InMux
    port map (
            O => \N__28254\,
            I => \N__28247\
        );

    \I__5804\ : InMux
    port map (
            O => \N__28253\,
            I => \N__28244\
        );

    \I__5803\ : Odrv4
    port map (
            O => \N__28250\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__28247\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__28244\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__5800\ : InMux
    port map (
            O => \N__28237\,
            I => \N__28234\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__28234\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_1_1_1\
        );

    \I__5798\ : InMux
    port map (
            O => \N__28231\,
            I => \N__28224\
        );

    \I__5797\ : InMux
    port map (
            O => \N__28230\,
            I => \N__28224\
        );

    \I__5796\ : InMux
    port map (
            O => \N__28229\,
            I => \N__28221\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__28224\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__28221\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__5793\ : CascadeMux
    port map (
            O => \N__28216\,
            I => \N__28212\
        );

    \I__5792\ : InMux
    port map (
            O => \N__28215\,
            I => \N__28209\
        );

    \I__5791\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28206\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__28209\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__28206\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__5788\ : InMux
    port map (
            O => \N__28201\,
            I => \N__28197\
        );

    \I__5787\ : InMux
    port map (
            O => \N__28200\,
            I => \N__28191\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__28197\,
            I => \N__28188\
        );

    \I__5785\ : InMux
    port map (
            O => \N__28196\,
            I => \N__28185\
        );

    \I__5784\ : InMux
    port map (
            O => \N__28195\,
            I => \N__28180\
        );

    \I__5783\ : InMux
    port map (
            O => \N__28194\,
            I => \N__28180\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__28191\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__28188\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__28185\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__28180\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__5778\ : CascadeMux
    port map (
            O => \N__28171\,
            I => \this_vga_signals.mult1_un54_sum_axb1_cascade_\
        );

    \I__5777\ : InMux
    port map (
            O => \N__28168\,
            I => \N__28157\
        );

    \I__5776\ : InMux
    port map (
            O => \N__28167\,
            I => \N__28157\
        );

    \I__5775\ : InMux
    port map (
            O => \N__28166\,
            I => \N__28150\
        );

    \I__5774\ : InMux
    port map (
            O => \N__28165\,
            I => \N__28150\
        );

    \I__5773\ : InMux
    port map (
            O => \N__28164\,
            I => \N__28150\
        );

    \I__5772\ : InMux
    port map (
            O => \N__28163\,
            I => \N__28145\
        );

    \I__5771\ : InMux
    port map (
            O => \N__28162\,
            I => \N__28145\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__28157\,
            I => \M_this_state_qZ0Z_18\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__28150\,
            I => \M_this_state_qZ0Z_18\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__28145\,
            I => \M_this_state_qZ0Z_18\
        );

    \I__5767\ : InMux
    port map (
            O => \N__28138\,
            I => \N__28135\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__28135\,
            I => \N__28132\
        );

    \I__5765\ : Odrv12
    port map (
            O => \N__28132\,
            I => \this_ppu_M_this_map_address_d_4_sqmuxa_0_a3_i_o3_i_a3_0\
        );

    \I__5764\ : CascadeMux
    port map (
            O => \N__28129\,
            I => \this_ppu.N_1322_cascade_\
        );

    \I__5763\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28123\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__28123\,
            I => \N__28119\
        );

    \I__5761\ : InMux
    port map (
            O => \N__28122\,
            I => \N__28116\
        );

    \I__5760\ : Span4Mux_v
    port map (
            O => \N__28119\,
            I => \N__28109\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__28116\,
            I => \N__28109\
        );

    \I__5758\ : InMux
    port map (
            O => \N__28115\,
            I => \N__28106\
        );

    \I__5757\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28102\
        );

    \I__5756\ : Span4Mux_v
    port map (
            O => \N__28109\,
            I => \N__28097\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__28106\,
            I => \N__28097\
        );

    \I__5754\ : InMux
    port map (
            O => \N__28105\,
            I => \N__28094\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__28102\,
            I => \N__28090\
        );

    \I__5752\ : Span4Mux_v
    port map (
            O => \N__28097\,
            I => \N__28085\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__28094\,
            I => \N__28085\
        );

    \I__5750\ : InMux
    port map (
            O => \N__28093\,
            I => \N__28082\
        );

    \I__5749\ : Span4Mux_h
    port map (
            O => \N__28090\,
            I => \N__28077\
        );

    \I__5748\ : Span4Mux_v
    port map (
            O => \N__28085\,
            I => \N__28072\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__28082\,
            I => \N__28072\
        );

    \I__5746\ : InMux
    port map (
            O => \N__28081\,
            I => \N__28069\
        );

    \I__5745\ : InMux
    port map (
            O => \N__28080\,
            I => \N__28066\
        );

    \I__5744\ : Span4Mux_h
    port map (
            O => \N__28077\,
            I => \N__28063\
        );

    \I__5743\ : Span4Mux_v
    port map (
            O => \N__28072\,
            I => \N__28058\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__28069\,
            I => \N__28058\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__28066\,
            I => \N__28055\
        );

    \I__5740\ : Span4Mux_h
    port map (
            O => \N__28063\,
            I => \N__28052\
        );

    \I__5739\ : Span4Mux_v
    port map (
            O => \N__28058\,
            I => \N__28047\
        );

    \I__5738\ : Span4Mux_v
    port map (
            O => \N__28055\,
            I => \N__28047\
        );

    \I__5737\ : Span4Mux_v
    port map (
            O => \N__28052\,
            I => \N__28042\
        );

    \I__5736\ : Span4Mux_h
    port map (
            O => \N__28047\,
            I => \N__28042\
        );

    \I__5735\ : Odrv4
    port map (
            O => \N__28042\,
            I => \M_this_spr_ram_write_data_0\
        );

    \I__5734\ : InMux
    port map (
            O => \N__28039\,
            I => \N__28035\
        );

    \I__5733\ : InMux
    port map (
            O => \N__28038\,
            I => \N__28032\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__28035\,
            I => \N__28026\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__28032\,
            I => \N__28023\
        );

    \I__5730\ : CascadeMux
    port map (
            O => \N__28031\,
            I => \N__28020\
        );

    \I__5729\ : InMux
    port map (
            O => \N__28030\,
            I => \N__28015\
        );

    \I__5728\ : InMux
    port map (
            O => \N__28029\,
            I => \N__28015\
        );

    \I__5727\ : Span4Mux_h
    port map (
            O => \N__28026\,
            I => \N__28012\
        );

    \I__5726\ : Span4Mux_h
    port map (
            O => \N__28023\,
            I => \N__28009\
        );

    \I__5725\ : InMux
    port map (
            O => \N__28020\,
            I => \N__28006\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__28015\,
            I => \N__28003\
        );

    \I__5723\ : Odrv4
    port map (
            O => \N__28012\,
            I => \this_vga_signals_CO0_0_i_i\
        );

    \I__5722\ : Odrv4
    port map (
            O => \N__28009\,
            I => \this_vga_signals_CO0_0_i_i\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__28006\,
            I => \this_vga_signals_CO0_0_i_i\
        );

    \I__5720\ : Odrv4
    port map (
            O => \N__28003\,
            I => \this_vga_signals_CO0_0_i_i\
        );

    \I__5719\ : CascadeMux
    port map (
            O => \N__27994\,
            I => \this_vga_signals_CO0_0_i_i_cascade_\
        );

    \I__5718\ : InMux
    port map (
            O => \N__27991\,
            I => \N__27986\
        );

    \I__5717\ : CascadeMux
    port map (
            O => \N__27990\,
            I => \N__27983\
        );

    \I__5716\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27979\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__27986\,
            I => \N__27976\
        );

    \I__5714\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27971\
        );

    \I__5713\ : InMux
    port map (
            O => \N__27982\,
            I => \N__27971\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__27979\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__5711\ : Odrv4
    port map (
            O => \N__27976\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__27971\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__5709\ : InMux
    port map (
            O => \N__27964\,
            I => \N__27961\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__27961\,
            I => \this_vga_signals.g1\
        );

    \I__5707\ : InMux
    port map (
            O => \N__27958\,
            I => \N__27953\
        );

    \I__5706\ : InMux
    port map (
            O => \N__27957\,
            I => \N__27950\
        );

    \I__5705\ : InMux
    port map (
            O => \N__27956\,
            I => \N__27946\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__27953\,
            I => \N__27940\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__27950\,
            I => \N__27940\
        );

    \I__5702\ : InMux
    port map (
            O => \N__27949\,
            I => \N__27937\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__27946\,
            I => \N__27934\
        );

    \I__5700\ : InMux
    port map (
            O => \N__27945\,
            I => \N__27931\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__27940\,
            I => \N__27922\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__27937\,
            I => \N__27922\
        );

    \I__5697\ : Span4Mux_h
    port map (
            O => \N__27934\,
            I => \N__27922\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__27931\,
            I => \N__27922\
        );

    \I__5695\ : Odrv4
    port map (
            O => \N__27922\,
            I => \this_vga_signals.N_39_0\
        );

    \I__5694\ : CascadeMux
    port map (
            O => \N__27919\,
            I => \N__27916\
        );

    \I__5693\ : InMux
    port map (
            O => \N__27916\,
            I => \N__27911\
        );

    \I__5692\ : InMux
    port map (
            O => \N__27915\,
            I => \N__27906\
        );

    \I__5691\ : InMux
    port map (
            O => \N__27914\,
            I => \N__27903\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__27911\,
            I => \N__27900\
        );

    \I__5689\ : InMux
    port map (
            O => \N__27910\,
            I => \N__27897\
        );

    \I__5688\ : InMux
    port map (
            O => \N__27909\,
            I => \N__27894\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__27906\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__27903\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__5685\ : Odrv4
    port map (
            O => \N__27900\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__27897\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__27894\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__5682\ : InMux
    port map (
            O => \N__27883\,
            I => \N__27880\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__27880\,
            I => \this_vga_signals.N_38_i_0_a2_0_4Z0Z_1\
        );

    \I__5680\ : CascadeMux
    port map (
            O => \N__27877\,
            I => \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_17_cascade_\
        );

    \I__5679\ : InMux
    port map (
            O => \N__27874\,
            I => \N__27868\
        );

    \I__5678\ : InMux
    port map (
            O => \N__27873\,
            I => \N__27865\
        );

    \I__5677\ : InMux
    port map (
            O => \N__27872\,
            I => \N__27860\
        );

    \I__5676\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27860\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__27868\,
            I => \M_this_state_qZ0Z_17\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__27865\,
            I => \M_this_state_qZ0Z_17\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__27860\,
            I => \M_this_state_qZ0Z_17\
        );

    \I__5672\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27850\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__27850\,
            I => \N__27847\
        );

    \I__5670\ : Odrv12
    port map (
            O => \N__27847\,
            I => \this_vga_signals.vsync_1_0_a3_0_a3_0\
        );

    \I__5669\ : InMux
    port map (
            O => \N__27844\,
            I => \N__27841\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__27841\,
            I => \this_vga_signals.N_2840_0_0\
        );

    \I__5667\ : InMux
    port map (
            O => \N__27838\,
            I => \N__27835\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__27835\,
            I => \this_vga_signals.N_27_0_0\
        );

    \I__5665\ : CascadeMux
    port map (
            O => \N__27832\,
            I => \this_vga_signals.vaddress_7_cascade_\
        );

    \I__5664\ : InMux
    port map (
            O => \N__27829\,
            I => \N__27825\
        );

    \I__5663\ : InMux
    port map (
            O => \N__27828\,
            I => \N__27822\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__27825\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__27822\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__5660\ : InMux
    port map (
            O => \N__27817\,
            I => \N__27813\
        );

    \I__5659\ : CascadeMux
    port map (
            O => \N__27816\,
            I => \N__27810\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__27813\,
            I => \N__27807\
        );

    \I__5657\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27804\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__27807\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__27804\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__5654\ : CascadeMux
    port map (
            O => \N__27799\,
            I => \this_vga_signals.g1_2_0_cascade_\
        );

    \I__5653\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27793\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__27793\,
            I => \N__27790\
        );

    \I__5651\ : Odrv4
    port map (
            O => \N__27790\,
            I => \this_vga_signals.if_m6_i_x2_3\
        );

    \I__5650\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27784\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__27784\,
            I => \this_vga_signals.g1_3\
        );

    \I__5648\ : CascadeMux
    port map (
            O => \N__27781\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0_ns_1_cascade_\
        );

    \I__5647\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27775\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__27775\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1\
        );

    \I__5645\ : InMux
    port map (
            O => \N__27772\,
            I => \N__27769\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__27769\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_1_0\
        );

    \I__5643\ : CascadeMux
    port map (
            O => \N__27766\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0_cascade_\
        );

    \I__5642\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27759\
        );

    \I__5641\ : InMux
    port map (
            O => \N__27762\,
            I => \N__27756\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__27759\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_1_1\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__27756\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_1_1\
        );

    \I__5638\ : CascadeMux
    port map (
            O => \N__27751\,
            I => \this_vga_signals.if_m5_s_cascade_\
        );

    \I__5637\ : CascadeMux
    port map (
            O => \N__27748\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_1_0_cascade_\
        );

    \I__5636\ : CascadeMux
    port map (
            O => \N__27745\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\
        );

    \I__5635\ : InMux
    port map (
            O => \N__27742\,
            I => \N__27739\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__27739\,
            I => \this_vga_signals.if_m5_d\
        );

    \I__5633\ : CascadeMux
    port map (
            O => \N__27736\,
            I => \this_vga_signals.if_m5_d_cascade_\
        );

    \I__5632\ : InMux
    port map (
            O => \N__27733\,
            I => \N__27730\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__27730\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_1\
        );

    \I__5630\ : CascadeMux
    port map (
            O => \N__27727\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_1_cascade_\
        );

    \I__5629\ : CascadeMux
    port map (
            O => \N__27724\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_x0_cascade_\
        );

    \I__5628\ : InMux
    port map (
            O => \N__27721\,
            I => \N__27718\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__27718\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_x1\
        );

    \I__5626\ : InMux
    port map (
            O => \N__27715\,
            I => \N__27712\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__27712\,
            I => \N__27709\
        );

    \I__5624\ : Span4Mux_v
    port map (
            O => \N__27709\,
            I => \N__27705\
        );

    \I__5623\ : InMux
    port map (
            O => \N__27708\,
            I => \N__27702\
        );

    \I__5622\ : Span4Mux_h
    port map (
            O => \N__27705\,
            I => \N__27699\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__27702\,
            I => \N__27696\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__27699\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__5619\ : Odrv12
    port map (
            O => \N__27696\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__5618\ : CascadeMux
    port map (
            O => \N__27691\,
            I => \this_vga_signals.N_38_i_0_a2_3_cascade_\
        );

    \I__5617\ : InMux
    port map (
            O => \N__27688\,
            I => \N__27685\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__27685\,
            I => \this_vga_signals.N_38_i_0_a2_0_3\
        );

    \I__5615\ : CascadeMux
    port map (
            O => \N__27682\,
            I => \N__27676\
        );

    \I__5614\ : CascadeMux
    port map (
            O => \N__27681\,
            I => \N__27672\
        );

    \I__5613\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27667\
        );

    \I__5612\ : InMux
    port map (
            O => \N__27679\,
            I => \N__27667\
        );

    \I__5611\ : InMux
    port map (
            O => \N__27676\,
            I => \N__27664\
        );

    \I__5610\ : InMux
    port map (
            O => \N__27675\,
            I => \N__27661\
        );

    \I__5609\ : InMux
    port map (
            O => \N__27672\,
            I => \N__27658\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__27667\,
            I => \N__27655\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__27664\,
            I => \N__27652\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__27661\,
            I => \N__27647\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__27658\,
            I => \N__27647\
        );

    \I__5604\ : Span4Mux_v
    port map (
            O => \N__27655\,
            I => \N__27642\
        );

    \I__5603\ : Span4Mux_v
    port map (
            O => \N__27652\,
            I => \N__27642\
        );

    \I__5602\ : Span4Mux_v
    port map (
            O => \N__27647\,
            I => \N__27639\
        );

    \I__5601\ : Span4Mux_v
    port map (
            O => \N__27642\,
            I => \N__27636\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__27639\,
            I => \N__27633\
        );

    \I__5599\ : Span4Mux_h
    port map (
            O => \N__27636\,
            I => \N__27630\
        );

    \I__5598\ : Span4Mux_v
    port map (
            O => \N__27633\,
            I => \N__27627\
        );

    \I__5597\ : Sp12to4
    port map (
            O => \N__27630\,
            I => \N__27622\
        );

    \I__5596\ : Sp12to4
    port map (
            O => \N__27627\,
            I => \N__27622\
        );

    \I__5595\ : Span12Mux_h
    port map (
            O => \N__27622\,
            I => \N__27619\
        );

    \I__5594\ : Odrv12
    port map (
            O => \N__27619\,
            I => port_enb_c
        );

    \I__5593\ : InMux
    port map (
            O => \N__27616\,
            I => \N__27610\
        );

    \I__5592\ : InMux
    port map (
            O => \N__27615\,
            I => \N__27607\
        );

    \I__5591\ : InMux
    port map (
            O => \N__27614\,
            I => \N__27604\
        );

    \I__5590\ : InMux
    port map (
            O => \N__27613\,
            I => \N__27601\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__27610\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__27607\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__27604\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__27601\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__5585\ : InMux
    port map (
            O => \N__27592\,
            I => \N__27589\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__27589\,
            I => \N__27582\
        );

    \I__5583\ : InMux
    port map (
            O => \N__27588\,
            I => \N__27577\
        );

    \I__5582\ : InMux
    port map (
            O => \N__27587\,
            I => \N__27577\
        );

    \I__5581\ : InMux
    port map (
            O => \N__27586\,
            I => \N__27572\
        );

    \I__5580\ : InMux
    port map (
            O => \N__27585\,
            I => \N__27572\
        );

    \I__5579\ : Odrv4
    port map (
            O => \N__27582\,
            I => \M_this_delay_clk_out_0\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__27577\,
            I => \M_this_delay_clk_out_0\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__27572\,
            I => \M_this_delay_clk_out_0\
        );

    \I__5576\ : CascadeMux
    port map (
            O => \N__27565\,
            I => \N_765_0_cascade_\
        );

    \I__5575\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27559\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__27559\,
            I => \N__27556\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__27556\,
            I => \this_ppu.N_229_1_0\
        );

    \I__5572\ : CascadeMux
    port map (
            O => \N__27553\,
            I => \this_ppu.N_229_1_0_cascade_\
        );

    \I__5571\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27532\
        );

    \I__5570\ : InMux
    port map (
            O => \N__27549\,
            I => \N__27532\
        );

    \I__5569\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27521\
        );

    \I__5568\ : InMux
    port map (
            O => \N__27547\,
            I => \N__27521\
        );

    \I__5567\ : InMux
    port map (
            O => \N__27546\,
            I => \N__27521\
        );

    \I__5566\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27521\
        );

    \I__5565\ : InMux
    port map (
            O => \N__27544\,
            I => \N__27521\
        );

    \I__5564\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27506\
        );

    \I__5563\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27506\
        );

    \I__5562\ : InMux
    port map (
            O => \N__27541\,
            I => \N__27506\
        );

    \I__5561\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27506\
        );

    \I__5560\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27506\
        );

    \I__5559\ : InMux
    port map (
            O => \N__27538\,
            I => \N__27506\
        );

    \I__5558\ : InMux
    port map (
            O => \N__27537\,
            I => \N__27506\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__27532\,
            I => \N__27501\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__27521\,
            I => \N__27501\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__27506\,
            I => \N__27498\
        );

    \I__5554\ : Span4Mux_h
    port map (
            O => \N__27501\,
            I => \N__27495\
        );

    \I__5553\ : Odrv4
    port map (
            O => \N__27498\,
            I => \N_229\
        );

    \I__5552\ : Odrv4
    port map (
            O => \N__27495\,
            I => \N_229\
        );

    \I__5551\ : CascadeMux
    port map (
            O => \N__27490\,
            I => \N__27486\
        );

    \I__5550\ : InMux
    port map (
            O => \N__27489\,
            I => \N__27483\
        );

    \I__5549\ : InMux
    port map (
            O => \N__27486\,
            I => \N__27477\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__27483\,
            I => \N__27474\
        );

    \I__5547\ : InMux
    port map (
            O => \N__27482\,
            I => \N__27467\
        );

    \I__5546\ : InMux
    port map (
            O => \N__27481\,
            I => \N__27467\
        );

    \I__5545\ : InMux
    port map (
            O => \N__27480\,
            I => \N__27467\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__27477\,
            I => \N__27460\
        );

    \I__5543\ : Span4Mux_h
    port map (
            O => \N__27474\,
            I => \N__27457\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__27467\,
            I => \N__27454\
        );

    \I__5541\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27445\
        );

    \I__5540\ : InMux
    port map (
            O => \N__27465\,
            I => \N__27445\
        );

    \I__5539\ : InMux
    port map (
            O => \N__27464\,
            I => \N__27445\
        );

    \I__5538\ : InMux
    port map (
            O => \N__27463\,
            I => \N__27445\
        );

    \I__5537\ : Odrv12
    port map (
            O => \N__27460\,
            I => \N_1423\
        );

    \I__5536\ : Odrv4
    port map (
            O => \N__27457\,
            I => \N_1423\
        );

    \I__5535\ : Odrv4
    port map (
            O => \N__27454\,
            I => \N_1423\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__27445\,
            I => \N_1423\
        );

    \I__5533\ : CascadeMux
    port map (
            O => \N__27436\,
            I => \this_vga_signals.SUM_2_i_i_1_0_3_cascade_\
        );

    \I__5532\ : InMux
    port map (
            O => \N__27433\,
            I => \N__27428\
        );

    \I__5531\ : InMux
    port map (
            O => \N__27432\,
            I => \N__27422\
        );

    \I__5530\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27419\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__27428\,
            I => \N__27416\
        );

    \I__5528\ : InMux
    port map (
            O => \N__27427\,
            I => \N__27411\
        );

    \I__5527\ : InMux
    port map (
            O => \N__27426\,
            I => \N__27411\
        );

    \I__5526\ : InMux
    port map (
            O => \N__27425\,
            I => \N__27408\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__27422\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__27419\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__5523\ : Odrv4
    port map (
            O => \N__27416\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__27411\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__27408\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__5520\ : InMux
    port map (
            O => \N__27397\,
            I => \N__27394\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__27394\,
            I => \N__27391\
        );

    \I__5518\ : Span4Mux_v
    port map (
            O => \N__27391\,
            I => \N__27388\
        );

    \I__5517\ : Odrv4
    port map (
            O => \N__27388\,
            I => \this_vga_signals.vsync_1_0_a3_0_a3_5\
        );

    \I__5516\ : InMux
    port map (
            O => \N__27385\,
            I => \N__27379\
        );

    \I__5515\ : InMux
    port map (
            O => \N__27384\,
            I => \N__27376\
        );

    \I__5514\ : InMux
    port map (
            O => \N__27383\,
            I => \N__27371\
        );

    \I__5513\ : InMux
    port map (
            O => \N__27382\,
            I => \N__27371\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__27379\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__27376\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__27371\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__5509\ : CascadeMux
    port map (
            O => \N__27364\,
            I => \this_ppu.N_430_1_0_cascade_\
        );

    \I__5508\ : InMux
    port map (
            O => \N__27361\,
            I => \N__27355\
        );

    \I__5507\ : InMux
    port map (
            O => \N__27360\,
            I => \N__27355\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__27355\,
            I => \M_this_state_q_fastZ0Z_13\
        );

    \I__5505\ : CascadeMux
    port map (
            O => \N__27352\,
            I => \this_vga_signals.N_38_i_0_a2_3Z0Z_0_cascade_\
        );

    \I__5504\ : CascadeMux
    port map (
            O => \N__27349\,
            I => \this_vga_signals.N_38_i_0_a2_3_xZ0Z1_cascade_\
        );

    \I__5503\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27336\
        );

    \I__5502\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27336\
        );

    \I__5501\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27336\
        );

    \I__5500\ : InMux
    port map (
            O => \N__27343\,
            I => \N__27330\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__27336\,
            I => \N__27323\
        );

    \I__5498\ : CEMux
    port map (
            O => \N__27335\,
            I => \N__27320\
        );

    \I__5497\ : InMux
    port map (
            O => \N__27334\,
            I => \N__27317\
        );

    \I__5496\ : InMux
    port map (
            O => \N__27333\,
            I => \N__27314\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__27330\,
            I => \N__27309\
        );

    \I__5494\ : InMux
    port map (
            O => \N__27329\,
            I => \N__27304\
        );

    \I__5493\ : InMux
    port map (
            O => \N__27328\,
            I => \N__27304\
        );

    \I__5492\ : InMux
    port map (
            O => \N__27327\,
            I => \N__27299\
        );

    \I__5491\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27299\
        );

    \I__5490\ : Span4Mux_v
    port map (
            O => \N__27323\,
            I => \N__27286\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__27320\,
            I => \N__27286\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__27317\,
            I => \N__27281\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__27314\,
            I => \N__27281\
        );

    \I__5486\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27274\
        );

    \I__5485\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27274\
        );

    \I__5484\ : Span12Mux_v
    port map (
            O => \N__27309\,
            I => \N__27271\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__27304\,
            I => \N__27266\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__27299\,
            I => \N__27266\
        );

    \I__5481\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27263\
        );

    \I__5480\ : InMux
    port map (
            O => \N__27297\,
            I => \N__27260\
        );

    \I__5479\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27255\
        );

    \I__5478\ : InMux
    port map (
            O => \N__27295\,
            I => \N__27255\
        );

    \I__5477\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27246\
        );

    \I__5476\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27246\
        );

    \I__5475\ : InMux
    port map (
            O => \N__27292\,
            I => \N__27246\
        );

    \I__5474\ : InMux
    port map (
            O => \N__27291\,
            I => \N__27246\
        );

    \I__5473\ : Span4Mux_v
    port map (
            O => \N__27286\,
            I => \N__27243\
        );

    \I__5472\ : Span4Mux_v
    port map (
            O => \N__27281\,
            I => \N__27240\
        );

    \I__5471\ : InMux
    port map (
            O => \N__27280\,
            I => \N__27235\
        );

    \I__5470\ : InMux
    port map (
            O => \N__27279\,
            I => \N__27235\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__27274\,
            I => \N__27230\
        );

    \I__5468\ : Span12Mux_h
    port map (
            O => \N__27271\,
            I => \N__27230\
        );

    \I__5467\ : Span12Mux_v
    port map (
            O => \N__27266\,
            I => \N__27225\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__27263\,
            I => \N__27225\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__27260\,
            I => \G_535\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__27255\,
            I => \G_535\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__27246\,
            I => \G_535\
        );

    \I__5462\ : Odrv4
    port map (
            O => \N__27243\,
            I => \G_535\
        );

    \I__5461\ : Odrv4
    port map (
            O => \N__27240\,
            I => \G_535\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__27235\,
            I => \G_535\
        );

    \I__5459\ : Odrv12
    port map (
            O => \N__27230\,
            I => \G_535\
        );

    \I__5458\ : Odrv12
    port map (
            O => \N__27225\,
            I => \G_535\
        );

    \I__5457\ : InMux
    port map (
            O => \N__27208\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_2\
        );

    \I__5456\ : InMux
    port map (
            O => \N__27205\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3\
        );

    \I__5455\ : InMux
    port map (
            O => \N__27202\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4\
        );

    \I__5454\ : InMux
    port map (
            O => \N__27199\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5\
        );

    \I__5453\ : InMux
    port map (
            O => \N__27196\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6\
        );

    \I__5452\ : InMux
    port map (
            O => \N__27193\,
            I => \bfn_18_22_0_\
        );

    \I__5451\ : InMux
    port map (
            O => \N__27190\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__27187\,
            I => \N__27184\
        );

    \I__5449\ : InMux
    port map (
            O => \N__27184\,
            I => \N__27181\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__27181\,
            I => \N__27178\
        );

    \I__5447\ : Span4Mux_v
    port map (
            O => \N__27178\,
            I => \N__27175\
        );

    \I__5446\ : Odrv4
    port map (
            O => \N__27175\,
            I => \this_vga_signals.g0_0_0\
        );

    \I__5445\ : InMux
    port map (
            O => \N__27172\,
            I => \N__27169\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__27169\,
            I => \N__27166\
        );

    \I__5443\ : Odrv12
    port map (
            O => \N__27166\,
            I => \this_vga_signals.IO_port_data_write_0_a2_i_o2_2Z0Z_1\
        );

    \I__5442\ : CascadeMux
    port map (
            O => \N__27163\,
            I => \N__27160\
        );

    \I__5441\ : InMux
    port map (
            O => \N__27160\,
            I => \N__27157\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__27157\,
            I => \N__27154\
        );

    \I__5439\ : Odrv4
    port map (
            O => \N__27154\,
            I => \this_vga_signals.mult1_un54_sum_2_1\
        );

    \I__5438\ : InMux
    port map (
            O => \N__27151\,
            I => \N__27148\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__27148\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0\
        );

    \I__5436\ : InMux
    port map (
            O => \N__27145\,
            I => \N__27142\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__27142\,
            I => \this_ppu.N_1115\
        );

    \I__5434\ : CascadeMux
    port map (
            O => \N__27139\,
            I => \N__27136\
        );

    \I__5433\ : InMux
    port map (
            O => \N__27136\,
            I => \N__27133\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__27133\,
            I => \this_vga_signals.g0_33_N_3L4\
        );

    \I__5431\ : InMux
    port map (
            O => \N__27130\,
            I => \N__27127\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__27127\,
            I => \this_vga_signals.g0_33_N_4L6\
        );

    \I__5429\ : InMux
    port map (
            O => \N__27124\,
            I => \N__27121\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__27121\,
            I => \this_vga_signals.g0_33_N_5L8\
        );

    \I__5427\ : CascadeMux
    port map (
            O => \N__27118\,
            I => \N__27113\
        );

    \I__5426\ : InMux
    port map (
            O => \N__27117\,
            I => \N__27110\
        );

    \I__5425\ : InMux
    port map (
            O => \N__27116\,
            I => \N__27107\
        );

    \I__5424\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27104\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__27110\,
            I => \N__27098\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__27107\,
            I => \N__27095\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__27104\,
            I => \N__27092\
        );

    \I__5420\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27089\
        );

    \I__5419\ : InMux
    port map (
            O => \N__27102\,
            I => \N__27086\
        );

    \I__5418\ : InMux
    port map (
            O => \N__27101\,
            I => \N__27083\
        );

    \I__5417\ : Span4Mux_v
    port map (
            O => \N__27098\,
            I => \N__27075\
        );

    \I__5416\ : Span4Mux_h
    port map (
            O => \N__27095\,
            I => \N__27075\
        );

    \I__5415\ : Span4Mux_v
    port map (
            O => \N__27092\,
            I => \N__27075\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__27089\,
            I => \N__27069\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__27086\,
            I => \N__27069\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__27083\,
            I => \N__27066\
        );

    \I__5411\ : InMux
    port map (
            O => \N__27082\,
            I => \N__27063\
        );

    \I__5410\ : Span4Mux_v
    port map (
            O => \N__27075\,
            I => \N__27058\
        );

    \I__5409\ : InMux
    port map (
            O => \N__27074\,
            I => \N__27055\
        );

    \I__5408\ : Span4Mux_h
    port map (
            O => \N__27069\,
            I => \N__27052\
        );

    \I__5407\ : Span4Mux_v
    port map (
            O => \N__27066\,
            I => \N__27047\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__27063\,
            I => \N__27047\
        );

    \I__5405\ : InMux
    port map (
            O => \N__27062\,
            I => \N__27042\
        );

    \I__5404\ : InMux
    port map (
            O => \N__27061\,
            I => \N__27042\
        );

    \I__5403\ : Sp12to4
    port map (
            O => \N__27058\,
            I => \N__27037\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__27055\,
            I => \N__27037\
        );

    \I__5401\ : Odrv4
    port map (
            O => \N__27052\,
            I => \this_vga_signals.M_hcounter_d7_0_i_0_0\
        );

    \I__5400\ : Odrv4
    port map (
            O => \N__27047\,
            I => \this_vga_signals.M_hcounter_d7_0_i_0_0\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__27042\,
            I => \this_vga_signals.M_hcounter_d7_0_i_0_0\
        );

    \I__5398\ : Odrv12
    port map (
            O => \N__27037\,
            I => \this_vga_signals.M_hcounter_d7_0_i_0_0\
        );

    \I__5397\ : InMux
    port map (
            O => \N__27028\,
            I => \N__27023\
        );

    \I__5396\ : InMux
    port map (
            O => \N__27027\,
            I => \N__27020\
        );

    \I__5395\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27017\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__27023\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__27020\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__27017\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__5391\ : InMux
    port map (
            O => \N__27010\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_0\
        );

    \I__5390\ : InMux
    port map (
            O => \N__27007\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_1\
        );

    \I__5389\ : InMux
    port map (
            O => \N__27004\,
            I => \N__27001\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__27001\,
            I => \this_vga_signals.mult1_un61_sum_axb2_i\
        );

    \I__5387\ : CascadeMux
    port map (
            O => \N__26998\,
            I => \N__26995\
        );

    \I__5386\ : CascadeBuf
    port map (
            O => \N__26995\,
            I => \N__26992\
        );

    \I__5385\ : CascadeMux
    port map (
            O => \N__26992\,
            I => \N__26989\
        );

    \I__5384\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26985\
        );

    \I__5383\ : InMux
    port map (
            O => \N__26988\,
            I => \N__26982\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__26985\,
            I => \N__26978\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__26982\,
            I => \N__26974\
        );

    \I__5380\ : CascadeMux
    port map (
            O => \N__26981\,
            I => \N__26971\
        );

    \I__5379\ : Span4Mux_v
    port map (
            O => \N__26978\,
            I => \N__26967\
        );

    \I__5378\ : InMux
    port map (
            O => \N__26977\,
            I => \N__26964\
        );

    \I__5377\ : Span4Mux_h
    port map (
            O => \N__26974\,
            I => \N__26961\
        );

    \I__5376\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26956\
        );

    \I__5375\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26956\
        );

    \I__5374\ : Sp12to4
    port map (
            O => \N__26967\,
            I => \N__26953\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__26964\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__5372\ : Odrv4
    port map (
            O => \N__26961\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__26956\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__5370\ : Odrv12
    port map (
            O => \N__26953\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__5369\ : InMux
    port map (
            O => \N__26944\,
            I => \N__26940\
        );

    \I__5368\ : InMux
    port map (
            O => \N__26943\,
            I => \N__26937\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__26940\,
            I => \un1_M_this_oam_address_q_c3\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__26937\,
            I => \un1_M_this_oam_address_q_c3\
        );

    \I__5365\ : CascadeMux
    port map (
            O => \N__26932\,
            I => \N__26929\
        );

    \I__5364\ : CascadeBuf
    port map (
            O => \N__26929\,
            I => \N__26926\
        );

    \I__5363\ : CascadeMux
    port map (
            O => \N__26926\,
            I => \N__26920\
        );

    \I__5362\ : CascadeMux
    port map (
            O => \N__26925\,
            I => \N__26917\
        );

    \I__5361\ : CascadeMux
    port map (
            O => \N__26924\,
            I => \N__26914\
        );

    \I__5360\ : InMux
    port map (
            O => \N__26923\,
            I => \N__26911\
        );

    \I__5359\ : InMux
    port map (
            O => \N__26920\,
            I => \N__26908\
        );

    \I__5358\ : InMux
    port map (
            O => \N__26917\,
            I => \N__26905\
        );

    \I__5357\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26902\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__26911\,
            I => \N__26897\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__26908\,
            I => \N__26897\
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__26905\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__26902\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__5352\ : Odrv12
    port map (
            O => \N__26897\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__5351\ : CascadeMux
    port map (
            O => \N__26890\,
            I => \N__26884\
        );

    \I__5350\ : CascadeMux
    port map (
            O => \N__26889\,
            I => \N__26881\
        );

    \I__5349\ : CascadeMux
    port map (
            O => \N__26888\,
            I => \N__26877\
        );

    \I__5348\ : InMux
    port map (
            O => \N__26887\,
            I => \N__26870\
        );

    \I__5347\ : InMux
    port map (
            O => \N__26884\,
            I => \N__26870\
        );

    \I__5346\ : InMux
    port map (
            O => \N__26881\,
            I => \N__26867\
        );

    \I__5345\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26860\
        );

    \I__5344\ : InMux
    port map (
            O => \N__26877\,
            I => \N__26860\
        );

    \I__5343\ : InMux
    port map (
            O => \N__26876\,
            I => \N__26860\
        );

    \I__5342\ : InMux
    port map (
            O => \N__26875\,
            I => \N__26857\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__26870\,
            I => \N__26854\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__26867\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__26860\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__26857\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__26854\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__5336\ : InMux
    port map (
            O => \N__26845\,
            I => \N__26835\
        );

    \I__5335\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26830\
        );

    \I__5334\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26830\
        );

    \I__5333\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26827\
        );

    \I__5332\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26824\
        );

    \I__5331\ : InMux
    port map (
            O => \N__26840\,
            I => \N__26819\
        );

    \I__5330\ : InMux
    port map (
            O => \N__26839\,
            I => \N__26819\
        );

    \I__5329\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26816\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__26835\,
            I => \N__26813\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__26830\,
            I => \N__26810\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__26827\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__26824\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__26819\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__26816\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__5322\ : Odrv4
    port map (
            O => \N__26813\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__5321\ : Odrv4
    port map (
            O => \N__26810\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__5320\ : CascadeMux
    port map (
            O => \N__26797\,
            I => \N__26793\
        );

    \I__5319\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26786\
        );

    \I__5318\ : InMux
    port map (
            O => \N__26793\,
            I => \N__26779\
        );

    \I__5317\ : InMux
    port map (
            O => \N__26792\,
            I => \N__26779\
        );

    \I__5316\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26779\
        );

    \I__5315\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26776\
        );

    \I__5314\ : InMux
    port map (
            O => \N__26789\,
            I => \N__26773\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__26786\,
            I => \N__26766\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__26779\,
            I => \N__26766\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__26776\,
            I => \N__26766\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__26773\,
            I => \N_778_0\
        );

    \I__5309\ : Odrv4
    port map (
            O => \N__26766\,
            I => \N_778_0\
        );

    \I__5308\ : InMux
    port map (
            O => \N__26761\,
            I => \N__26754\
        );

    \I__5307\ : InMux
    port map (
            O => \N__26760\,
            I => \N__26749\
        );

    \I__5306\ : InMux
    port map (
            O => \N__26759\,
            I => \N__26749\
        );

    \I__5305\ : CEMux
    port map (
            O => \N__26758\,
            I => \N__26744\
        );

    \I__5304\ : CEMux
    port map (
            O => \N__26757\,
            I => \N__26741\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__26754\,
            I => \N__26713\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__26749\,
            I => \N__26713\
        );

    \I__5301\ : InMux
    port map (
            O => \N__26748\,
            I => \N__26708\
        );

    \I__5300\ : InMux
    port map (
            O => \N__26747\,
            I => \N__26708\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__26744\,
            I => \N__26703\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__26741\,
            I => \N__26703\
        );

    \I__5297\ : InMux
    port map (
            O => \N__26740\,
            I => \N__26698\
        );

    \I__5296\ : InMux
    port map (
            O => \N__26739\,
            I => \N__26698\
        );

    \I__5295\ : InMux
    port map (
            O => \N__26738\,
            I => \N__26689\
        );

    \I__5294\ : InMux
    port map (
            O => \N__26737\,
            I => \N__26689\
        );

    \I__5293\ : InMux
    port map (
            O => \N__26736\,
            I => \N__26689\
        );

    \I__5292\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26689\
        );

    \I__5291\ : InMux
    port map (
            O => \N__26734\,
            I => \N__26680\
        );

    \I__5290\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26680\
        );

    \I__5289\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26680\
        );

    \I__5288\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26680\
        );

    \I__5287\ : InMux
    port map (
            O => \N__26730\,
            I => \N__26675\
        );

    \I__5286\ : InMux
    port map (
            O => \N__26729\,
            I => \N__26675\
        );

    \I__5285\ : InMux
    port map (
            O => \N__26728\,
            I => \N__26667\
        );

    \I__5284\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26667\
        );

    \I__5283\ : InMux
    port map (
            O => \N__26726\,
            I => \N__26667\
        );

    \I__5282\ : InMux
    port map (
            O => \N__26725\,
            I => \N__26658\
        );

    \I__5281\ : InMux
    port map (
            O => \N__26724\,
            I => \N__26658\
        );

    \I__5280\ : InMux
    port map (
            O => \N__26723\,
            I => \N__26658\
        );

    \I__5279\ : InMux
    port map (
            O => \N__26722\,
            I => \N__26658\
        );

    \I__5278\ : InMux
    port map (
            O => \N__26721\,
            I => \N__26649\
        );

    \I__5277\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26649\
        );

    \I__5276\ : InMux
    port map (
            O => \N__26719\,
            I => \N__26649\
        );

    \I__5275\ : InMux
    port map (
            O => \N__26718\,
            I => \N__26649\
        );

    \I__5274\ : Span4Mux_h
    port map (
            O => \N__26713\,
            I => \N__26644\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__26708\,
            I => \N__26644\
        );

    \I__5272\ : Span4Mux_v
    port map (
            O => \N__26703\,
            I => \N__26638\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__26698\,
            I => \N__26633\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__26689\,
            I => \N__26633\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__26680\,
            I => \N__26628\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__26675\,
            I => \N__26628\
        );

    \I__5267\ : InMux
    port map (
            O => \N__26674\,
            I => \N__26625\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__26667\,
            I => \N__26618\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__26658\,
            I => \N__26618\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__26649\,
            I => \N__26618\
        );

    \I__5263\ : Span4Mux_v
    port map (
            O => \N__26644\,
            I => \N__26615\
        );

    \I__5262\ : InMux
    port map (
            O => \N__26643\,
            I => \N__26612\
        );

    \I__5261\ : InMux
    port map (
            O => \N__26642\,
            I => \N__26609\
        );

    \I__5260\ : InMux
    port map (
            O => \N__26641\,
            I => \N__26606\
        );

    \I__5259\ : Span4Mux_h
    port map (
            O => \N__26638\,
            I => \N__26599\
        );

    \I__5258\ : Span4Mux_v
    port map (
            O => \N__26633\,
            I => \N__26599\
        );

    \I__5257\ : Span4Mux_h
    port map (
            O => \N__26628\,
            I => \N__26599\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__26625\,
            I => \N__26594\
        );

    \I__5255\ : Span4Mux_h
    port map (
            O => \N__26618\,
            I => \N__26594\
        );

    \I__5254\ : Sp12to4
    port map (
            O => \N__26615\,
            I => \N__26585\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__26612\,
            I => \N__26585\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__26609\,
            I => \N__26585\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__26606\,
            I => \N__26585\
        );

    \I__5250\ : Span4Mux_h
    port map (
            O => \N__26599\,
            I => \N__26582\
        );

    \I__5249\ : Span4Mux_h
    port map (
            O => \N__26594\,
            I => \N__26579\
        );

    \I__5248\ : Odrv12
    port map (
            O => \N__26585\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__26582\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__5246\ : Odrv4
    port map (
            O => \N__26579\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__5245\ : CascadeMux
    port map (
            O => \N__26572\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1_cascade_\
        );

    \I__5244\ : CascadeMux
    port map (
            O => \N__26569\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_1_cascade_\
        );

    \I__5243\ : CascadeMux
    port map (
            O => \N__26566\,
            I => \N_778_0_cascade_\
        );

    \I__5242\ : CEMux
    port map (
            O => \N__26563\,
            I => \N__26560\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__26560\,
            I => \N__26555\
        );

    \I__5240\ : CEMux
    port map (
            O => \N__26559\,
            I => \N__26552\
        );

    \I__5239\ : CEMux
    port map (
            O => \N__26558\,
            I => \N__26549\
        );

    \I__5238\ : Span4Mux_h
    port map (
            O => \N__26555\,
            I => \N__26544\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__26552\,
            I => \N__26544\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__26549\,
            I => \N__26541\
        );

    \I__5235\ : Span4Mux_h
    port map (
            O => \N__26544\,
            I => \N__26538\
        );

    \I__5234\ : Span4Mux_h
    port map (
            O => \N__26541\,
            I => \N__26535\
        );

    \I__5233\ : Span4Mux_v
    port map (
            O => \N__26538\,
            I => \N__26532\
        );

    \I__5232\ : Odrv4
    port map (
            O => \N__26535\,
            I => \N_1701_0\
        );

    \I__5231\ : Odrv4
    port map (
            O => \N__26532\,
            I => \N_1701_0\
        );

    \I__5230\ : InMux
    port map (
            O => \N__26527\,
            I => \N__26524\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__26524\,
            I => \un1_M_this_oam_address_q_c5\
        );

    \I__5228\ : CascadeMux
    port map (
            O => \N__26521\,
            I => \N__26518\
        );

    \I__5227\ : CascadeBuf
    port map (
            O => \N__26518\,
            I => \N__26515\
        );

    \I__5226\ : CascadeMux
    port map (
            O => \N__26515\,
            I => \N__26511\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__26514\,
            I => \N__26508\
        );

    \I__5224\ : InMux
    port map (
            O => \N__26511\,
            I => \N__26505\
        );

    \I__5223\ : InMux
    port map (
            O => \N__26508\,
            I => \N__26502\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__26505\,
            I => \N__26499\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__26502\,
            I => \N__26494\
        );

    \I__5220\ : Sp12to4
    port map (
            O => \N__26499\,
            I => \N__26491\
        );

    \I__5219\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26486\
        );

    \I__5218\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26486\
        );

    \I__5217\ : Span4Mux_v
    port map (
            O => \N__26494\,
            I => \N__26483\
        );

    \I__5216\ : Span12Mux_s7_v
    port map (
            O => \N__26491\,
            I => \N__26480\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__26486\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__5214\ : Odrv4
    port map (
            O => \N__26483\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__5213\ : Odrv12
    port map (
            O => \N__26480\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__26473\,
            I => \un1_M_this_oam_address_q_c5_cascade_\
        );

    \I__5211\ : CascadeMux
    port map (
            O => \N__26470\,
            I => \N__26467\
        );

    \I__5210\ : CascadeBuf
    port map (
            O => \N__26467\,
            I => \N__26464\
        );

    \I__5209\ : CascadeMux
    port map (
            O => \N__26464\,
            I => \N__26461\
        );

    \I__5208\ : InMux
    port map (
            O => \N__26461\,
            I => \N__26458\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__26458\,
            I => \N__26454\
        );

    \I__5206\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26451\
        );

    \I__5205\ : Span4Mux_h
    port map (
            O => \N__26454\,
            I => \N__26448\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__26451\,
            I => \N__26442\
        );

    \I__5203\ : Span4Mux_h
    port map (
            O => \N__26448\,
            I => \N__26442\
        );

    \I__5202\ : InMux
    port map (
            O => \N__26447\,
            I => \N__26439\
        );

    \I__5201\ : Span4Mux_h
    port map (
            O => \N__26442\,
            I => \N__26436\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__26439\,
            I => \M_this_oam_address_qZ0Z_6\
        );

    \I__5199\ : Odrv4
    port map (
            O => \N__26436\,
            I => \M_this_oam_address_qZ0Z_6\
        );

    \I__5198\ : InMux
    port map (
            O => \N__26431\,
            I => \N__26428\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__26428\,
            I => \N__26423\
        );

    \I__5196\ : InMux
    port map (
            O => \N__26427\,
            I => \N__26418\
        );

    \I__5195\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26418\
        );

    \I__5194\ : Odrv4
    port map (
            O => \N__26423\,
            I => \un1_M_this_oam_address_q_c2\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__26418\,
            I => \un1_M_this_oam_address_q_c2\
        );

    \I__5192\ : CascadeMux
    port map (
            O => \N__26413\,
            I => \N__26410\
        );

    \I__5191\ : CascadeBuf
    port map (
            O => \N__26410\,
            I => \N__26407\
        );

    \I__5190\ : CascadeMux
    port map (
            O => \N__26407\,
            I => \N__26404\
        );

    \I__5189\ : InMux
    port map (
            O => \N__26404\,
            I => \N__26400\
        );

    \I__5188\ : CascadeMux
    port map (
            O => \N__26403\,
            I => \N__26394\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__26400\,
            I => \N__26391\
        );

    \I__5186\ : InMux
    port map (
            O => \N__26399\,
            I => \N__26388\
        );

    \I__5185\ : InMux
    port map (
            O => \N__26398\,
            I => \N__26383\
        );

    \I__5184\ : InMux
    port map (
            O => \N__26397\,
            I => \N__26383\
        );

    \I__5183\ : InMux
    port map (
            O => \N__26394\,
            I => \N__26380\
        );

    \I__5182\ : Span12Mux_s8_h
    port map (
            O => \N__26391\,
            I => \N__26377\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__26388\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__26383\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__26380\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__5178\ : Odrv12
    port map (
            O => \N__26377\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__5177\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26364\
        );

    \I__5176\ : InMux
    port map (
            O => \N__26367\,
            I => \N__26361\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__26364\,
            I => \N__26358\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__26361\,
            I => \N__26354\
        );

    \I__5173\ : Span4Mux_h
    port map (
            O => \N__26358\,
            I => \N__26351\
        );

    \I__5172\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26348\
        );

    \I__5171\ : Odrv12
    port map (
            O => \N__26354\,
            I => \N_782_0\
        );

    \I__5170\ : Odrv4
    port map (
            O => \N__26351\,
            I => \N_782_0\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__26348\,
            I => \N_782_0\
        );

    \I__5168\ : CEMux
    port map (
            O => \N__26341\,
            I => \N__26338\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__26338\,
            I => \N__26335\
        );

    \I__5166\ : Span4Mux_h
    port map (
            O => \N__26335\,
            I => \N__26332\
        );

    \I__5165\ : Span4Mux_h
    port map (
            O => \N__26332\,
            I => \N__26329\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__26329\,
            I => \N_1725_0\
        );

    \I__5163\ : CEMux
    port map (
            O => \N__26326\,
            I => \N__26323\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__26323\,
            I => \N__26320\
        );

    \I__5161\ : Span4Mux_v
    port map (
            O => \N__26320\,
            I => \N__26317\
        );

    \I__5160\ : Odrv4
    port map (
            O => \N__26317\,
            I => \N_1717_0\
        );

    \I__5159\ : InMux
    port map (
            O => \N__26314\,
            I => \N__26311\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__26311\,
            I => \N__26308\
        );

    \I__5157\ : Odrv4
    port map (
            O => \N__26308\,
            I => \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_12\
        );

    \I__5156\ : InMux
    port map (
            O => \N__26305\,
            I => \N__26302\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__26302\,
            I => \N__26299\
        );

    \I__5154\ : Span4Mux_h
    port map (
            O => \N__26299\,
            I => \N__26296\
        );

    \I__5153\ : Span4Mux_h
    port map (
            O => \N__26296\,
            I => \N__26293\
        );

    \I__5152\ : Odrv4
    port map (
            O => \N__26293\,
            I => \this_delay_clk.M_pipe_qZ0Z_3\
        );

    \I__5151\ : InMux
    port map (
            O => \N__26290\,
            I => \N__26287\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__26287\,
            I => \N__26284\
        );

    \I__5149\ : Span4Mux_h
    port map (
            O => \N__26284\,
            I => \N__26280\
        );

    \I__5148\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26277\
        );

    \I__5147\ : Odrv4
    port map (
            O => \N__26280\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_16\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__26277\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_16\
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__26272\,
            I => \N__26269\
        );

    \I__5144\ : InMux
    port map (
            O => \N__26269\,
            I => \N__26266\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__26266\,
            I => \N__26262\
        );

    \I__5142\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26259\
        );

    \I__5141\ : Odrv4
    port map (
            O => \N__26262\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_16\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__26259\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_16\
        );

    \I__5139\ : InMux
    port map (
            O => \N__26254\,
            I => \N__26250\
        );

    \I__5138\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26247\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__26250\,
            I => \N__26244\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__26247\,
            I => \N__26241\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__26244\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_10Z0Z_16\
        );

    \I__5134\ : Odrv4
    port map (
            O => \N__26241\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_10Z0Z_16\
        );

    \I__5133\ : CascadeMux
    port map (
            O => \N__26236\,
            I => \N__26232\
        );

    \I__5132\ : CascadeMux
    port map (
            O => \N__26235\,
            I => \N__26229\
        );

    \I__5131\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26225\
        );

    \I__5130\ : InMux
    port map (
            O => \N__26229\,
            I => \N__26222\
        );

    \I__5129\ : CascadeMux
    port map (
            O => \N__26228\,
            I => \N__26219\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__26225\,
            I => \N__26216\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__26222\,
            I => \N__26213\
        );

    \I__5126\ : InMux
    port map (
            O => \N__26219\,
            I => \N__26210\
        );

    \I__5125\ : Odrv12
    port map (
            O => \N__26216\,
            I => \N_771_0\
        );

    \I__5124\ : Odrv12
    port map (
            O => \N__26213\,
            I => \N_771_0\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__26210\,
            I => \N_771_0\
        );

    \I__5122\ : CascadeMux
    port map (
            O => \N__26203\,
            I => \N_771_0_cascade_\
        );

    \I__5121\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26196\
        );

    \I__5120\ : InMux
    port map (
            O => \N__26199\,
            I => \N__26193\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__26196\,
            I => \N__26190\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__26193\,
            I => \N__26187\
        );

    \I__5117\ : Span4Mux_h
    port map (
            O => \N__26190\,
            I => \N__26184\
        );

    \I__5116\ : Span4Mux_v
    port map (
            O => \N__26187\,
            I => \N__26181\
        );

    \I__5115\ : Span4Mux_h
    port map (
            O => \N__26184\,
            I => \N__26178\
        );

    \I__5114\ : Odrv4
    port map (
            O => \N__26181\,
            I => \this_ppu.N_774_0\
        );

    \I__5113\ : Odrv4
    port map (
            O => \N__26178\,
            I => \this_ppu.N_774_0\
        );

    \I__5112\ : CascadeMux
    port map (
            O => \N__26173\,
            I => \this_vga_signals.g1_0_0_cascade_\
        );

    \I__5111\ : InMux
    port map (
            O => \N__26170\,
            I => \N__26167\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__26167\,
            I => \this_vga_signals.if_N_6_0_0_0\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__26164\,
            I => \N__26161\
        );

    \I__5108\ : InMux
    port map (
            O => \N__26161\,
            I => \N__26158\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__26158\,
            I => \this_vga_signals.g1_0_0\
        );

    \I__5106\ : CascadeMux
    port map (
            O => \N__26155\,
            I => \this_vga_signals.N_27_0_1_0_cascade_\
        );

    \I__5105\ : InMux
    port map (
            O => \N__26152\,
            I => \N__26149\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__26149\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0\
        );

    \I__5103\ : CascadeMux
    port map (
            O => \N__26146\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_1_0_cascade_\
        );

    \I__5102\ : CascadeMux
    port map (
            O => \N__26143\,
            I => \N__26138\
        );

    \I__5101\ : CascadeMux
    port map (
            O => \N__26142\,
            I => \N__26132\
        );

    \I__5100\ : CascadeMux
    port map (
            O => \N__26141\,
            I => \N__26125\
        );

    \I__5099\ : InMux
    port map (
            O => \N__26138\,
            I => \N__26122\
        );

    \I__5098\ : InMux
    port map (
            O => \N__26137\,
            I => \N__26119\
        );

    \I__5097\ : InMux
    port map (
            O => \N__26136\,
            I => \N__26112\
        );

    \I__5096\ : InMux
    port map (
            O => \N__26135\,
            I => \N__26109\
        );

    \I__5095\ : InMux
    port map (
            O => \N__26132\,
            I => \N__26106\
        );

    \I__5094\ : InMux
    port map (
            O => \N__26131\,
            I => \N__26103\
        );

    \I__5093\ : InMux
    port map (
            O => \N__26130\,
            I => \N__26098\
        );

    \I__5092\ : InMux
    port map (
            O => \N__26129\,
            I => \N__26098\
        );

    \I__5091\ : InMux
    port map (
            O => \N__26128\,
            I => \N__26093\
        );

    \I__5090\ : InMux
    port map (
            O => \N__26125\,
            I => \N__26093\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__26122\,
            I => \N__26090\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__26119\,
            I => \N__26087\
        );

    \I__5087\ : InMux
    port map (
            O => \N__26118\,
            I => \N__26081\
        );

    \I__5086\ : InMux
    port map (
            O => \N__26117\,
            I => \N__26081\
        );

    \I__5085\ : IoInMux
    port map (
            O => \N__26116\,
            I => \N__26078\
        );

    \I__5084\ : InMux
    port map (
            O => \N__26115\,
            I => \N__26070\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__26112\,
            I => \N__26067\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__26109\,
            I => \N__26064\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__26106\,
            I => \N__26051\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__26103\,
            I => \N__26051\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__26098\,
            I => \N__26051\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__26093\,
            I => \N__26051\
        );

    \I__5077\ : Span4Mux_h
    port map (
            O => \N__26090\,
            I => \N__26051\
        );

    \I__5076\ : Span4Mux_v
    port map (
            O => \N__26087\,
            I => \N__26051\
        );

    \I__5075\ : InMux
    port map (
            O => \N__26086\,
            I => \N__26048\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__26081\,
            I => \N__26045\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__26078\,
            I => \N__26042\
        );

    \I__5072\ : InMux
    port map (
            O => \N__26077\,
            I => \N__26039\
        );

    \I__5071\ : InMux
    port map (
            O => \N__26076\,
            I => \N__26036\
        );

    \I__5070\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26033\
        );

    \I__5069\ : InMux
    port map (
            O => \N__26074\,
            I => \N__26028\
        );

    \I__5068\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26028\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__26070\,
            I => \N__26025\
        );

    \I__5066\ : Span4Mux_v
    port map (
            O => \N__26067\,
            I => \N__26018\
        );

    \I__5065\ : Span4Mux_v
    port map (
            O => \N__26064\,
            I => \N__26018\
        );

    \I__5064\ : Span4Mux_v
    port map (
            O => \N__26051\,
            I => \N__26018\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__26048\,
            I => \N__26013\
        );

    \I__5062\ : Span4Mux_h
    port map (
            O => \N__26045\,
            I => \N__26013\
        );

    \I__5061\ : Span12Mux_s6_h
    port map (
            O => \N__26042\,
            I => \N__26010\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__26039\,
            I => \M_this_reset_cond_out_0\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__26036\,
            I => \M_this_reset_cond_out_0\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__26033\,
            I => \M_this_reset_cond_out_0\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__26028\,
            I => \M_this_reset_cond_out_0\
        );

    \I__5056\ : Odrv4
    port map (
            O => \N__26025\,
            I => \M_this_reset_cond_out_0\
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__26018\,
            I => \M_this_reset_cond_out_0\
        );

    \I__5054\ : Odrv4
    port map (
            O => \N__26013\,
            I => \M_this_reset_cond_out_0\
        );

    \I__5053\ : Odrv12
    port map (
            O => \N__26010\,
            I => \M_this_reset_cond_out_0\
        );

    \I__5052\ : CascadeMux
    port map (
            O => \N__25993\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_2_cascade_\
        );

    \I__5051\ : CascadeMux
    port map (
            O => \N__25990\,
            I => \N__25987\
        );

    \I__5050\ : InMux
    port map (
            O => \N__25987\,
            I => \N__25984\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__25984\,
            I => \this_vga_signals.N_4_0\
        );

    \I__5048\ : InMux
    port map (
            O => \N__25981\,
            I => \N__25978\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__25978\,
            I => \this_vga_signals.if_m1_0_x2_1\
        );

    \I__5046\ : InMux
    port map (
            O => \N__25975\,
            I => \N__25972\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__25972\,
            I => \this_vga_signals.r_N_2_i_0\
        );

    \I__5044\ : CascadeMux
    port map (
            O => \N__25969\,
            I => \N__25965\
        );

    \I__5043\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25962\
        );

    \I__5042\ : InMux
    port map (
            O => \N__25965\,
            I => \N__25958\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__25962\,
            I => \N__25955\
        );

    \I__5040\ : InMux
    port map (
            O => \N__25961\,
            I => \N__25952\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__25958\,
            I => \N__25949\
        );

    \I__5038\ : Odrv4
    port map (
            O => \N__25955\,
            I => \this_vga_signals.N_836_0\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__25952\,
            I => \this_vga_signals.N_836_0\
        );

    \I__5036\ : Odrv12
    port map (
            O => \N__25949\,
            I => \this_vga_signals.N_836_0\
        );

    \I__5035\ : CascadeMux
    port map (
            O => \N__25942\,
            I => \this_vga_signals.N_1043_cascade_\
        );

    \I__5034\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25933\
        );

    \I__5033\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25933\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__25933\,
            I => \N__25928\
        );

    \I__5031\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25923\
        );

    \I__5030\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25923\
        );

    \I__5029\ : Odrv4
    port map (
            O => \N__25928\,
            I => \this_vga_signals_M_lcounter_q_0\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__25923\,
            I => \this_vga_signals_M_lcounter_q_0\
        );

    \I__5027\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25913\
        );

    \I__5026\ : InMux
    port map (
            O => \N__25917\,
            I => \N__25910\
        );

    \I__5025\ : InMux
    port map (
            O => \N__25916\,
            I => \N__25907\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__25913\,
            I => \N__25899\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__25910\,
            I => \N__25899\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__25907\,
            I => \N__25899\
        );

    \I__5021\ : InMux
    port map (
            O => \N__25906\,
            I => \N__25896\
        );

    \I__5020\ : Odrv12
    port map (
            O => \N__25899\,
            I => \N_792_0\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__25896\,
            I => \N_792_0\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__25891\,
            I => \N__25888\
        );

    \I__5017\ : InMux
    port map (
            O => \N__25888\,
            I => \N__25880\
        );

    \I__5016\ : InMux
    port map (
            O => \N__25887\,
            I => \N__25880\
        );

    \I__5015\ : CascadeMux
    port map (
            O => \N__25886\,
            I => \N__25876\
        );

    \I__5014\ : CascadeMux
    port map (
            O => \N__25885\,
            I => \N__25873\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__25880\,
            I => \N__25870\
        );

    \I__5012\ : InMux
    port map (
            O => \N__25879\,
            I => \N__25863\
        );

    \I__5011\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25863\
        );

    \I__5010\ : InMux
    port map (
            O => \N__25873\,
            I => \N__25863\
        );

    \I__5009\ : Span4Mux_v
    port map (
            O => \N__25870\,
            I => \N__25860\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__25863\,
            I => \this_vga_signals_M_lcounter_q_1\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__25860\,
            I => \this_vga_signals_M_lcounter_q_1\
        );

    \I__5006\ : InMux
    port map (
            O => \N__25855\,
            I => \N__25852\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__25852\,
            I => \N__25849\
        );

    \I__5004\ : Odrv4
    port map (
            O => \N__25849\,
            I => \this_ppu.M_last_q_0\
        );

    \I__5003\ : InMux
    port map (
            O => \N__25846\,
            I => \N__25843\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__25843\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_4_1_0_x1\
        );

    \I__5001\ : CascadeMux
    port map (
            O => \N__25840\,
            I => \N__25837\
        );

    \I__5000\ : InMux
    port map (
            O => \N__25837\,
            I => \N__25834\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__25834\,
            I => \M_this_scroll_qZ0Z_10\
        );

    \I__4998\ : InMux
    port map (
            O => \N__25831\,
            I => \N__25828\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__25828\,
            I => \N__25825\
        );

    \I__4996\ : Odrv12
    port map (
            O => \N__25825\,
            I => \M_this_scroll_qZ0Z_11\
        );

    \I__4995\ : CascadeMux
    port map (
            O => \N__25822\,
            I => \N__25819\
        );

    \I__4994\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25816\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__25816\,
            I => \N__25813\
        );

    \I__4992\ : Span4Mux_v
    port map (
            O => \N__25813\,
            I => \N__25810\
        );

    \I__4991\ : Span4Mux_h
    port map (
            O => \N__25810\,
            I => \N__25807\
        );

    \I__4990\ : Odrv4
    port map (
            O => \N__25807\,
            I => \M_this_scroll_qZ0Z_12\
        );

    \I__4989\ : InMux
    port map (
            O => \N__25804\,
            I => \N__25801\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__25801\,
            I => \N__25798\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__25798\,
            I => \M_this_scroll_qZ0Z_13\
        );

    \I__4986\ : CascadeMux
    port map (
            O => \N__25795\,
            I => \N__25792\
        );

    \I__4985\ : InMux
    port map (
            O => \N__25792\,
            I => \N__25789\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__25789\,
            I => \N__25786\
        );

    \I__4983\ : Span4Mux_h
    port map (
            O => \N__25786\,
            I => \N__25783\
        );

    \I__4982\ : Odrv4
    port map (
            O => \N__25783\,
            I => \M_this_scroll_qZ0Z_14\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__25780\,
            I => \N__25777\
        );

    \I__4980\ : InMux
    port map (
            O => \N__25777\,
            I => \N__25774\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__25774\,
            I => \N__25771\
        );

    \I__4978\ : Span4Mux_h
    port map (
            O => \N__25771\,
            I => \N__25768\
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__25768\,
            I => \M_this_scroll_qZ0Z_15\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__25765\,
            I => \N__25762\
        );

    \I__4975\ : InMux
    port map (
            O => \N__25762\,
            I => \N__25759\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__25759\,
            I => \N__25756\
        );

    \I__4973\ : Odrv4
    port map (
            O => \N__25756\,
            I => \M_this_scroll_qZ0Z_8\
        );

    \I__4972\ : InMux
    port map (
            O => \N__25753\,
            I => \N__25750\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__25750\,
            I => \N__25747\
        );

    \I__4970\ : Span4Mux_h
    port map (
            O => \N__25747\,
            I => \N__25744\
        );

    \I__4969\ : Odrv4
    port map (
            O => \N__25744\,
            I => \M_this_scroll_qZ0Z_9\
        );

    \I__4968\ : InMux
    port map (
            O => \N__25741\,
            I => \N__25738\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__25738\,
            I => \N__25734\
        );

    \I__4966\ : InMux
    port map (
            O => \N__25737\,
            I => \N__25730\
        );

    \I__4965\ : Span4Mux_v
    port map (
            O => \N__25734\,
            I => \N__25727\
        );

    \I__4964\ : InMux
    port map (
            O => \N__25733\,
            I => \N__25724\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__25730\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__4962\ : Odrv4
    port map (
            O => \N__25727\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__25724\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__4960\ : CascadeMux
    port map (
            O => \N__25717\,
            I => \N__25712\
        );

    \I__4959\ : InMux
    port map (
            O => \N__25716\,
            I => \N__25709\
        );

    \I__4958\ : InMux
    port map (
            O => \N__25715\,
            I => \N__25706\
        );

    \I__4957\ : InMux
    port map (
            O => \N__25712\,
            I => \N__25703\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__25709\,
            I => \N__25700\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__25706\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__25703\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__4953\ : Odrv4
    port map (
            O => \N__25700\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__4952\ : InMux
    port map (
            O => \N__25693\,
            I => \N__25690\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__25690\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_16\
        );

    \I__4950\ : CEMux
    port map (
            O => \N__25687\,
            I => \N__25682\
        );

    \I__4949\ : CEMux
    port map (
            O => \N__25686\,
            I => \N__25678\
        );

    \I__4948\ : CEMux
    port map (
            O => \N__25685\,
            I => \N__25675\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__25682\,
            I => \N__25672\
        );

    \I__4946\ : CEMux
    port map (
            O => \N__25681\,
            I => \N__25669\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__25678\,
            I => \N__25665\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__25675\,
            I => \N__25662\
        );

    \I__4943\ : Span4Mux_v
    port map (
            O => \N__25672\,
            I => \N__25657\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__25669\,
            I => \N__25657\
        );

    \I__4941\ : CEMux
    port map (
            O => \N__25668\,
            I => \N__25654\
        );

    \I__4940\ : Span4Mux_v
    port map (
            O => \N__25665\,
            I => \N__25651\
        );

    \I__4939\ : Span4Mux_v
    port map (
            O => \N__25662\,
            I => \N__25644\
        );

    \I__4938\ : Span4Mux_v
    port map (
            O => \N__25657\,
            I => \N__25644\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__25654\,
            I => \N__25644\
        );

    \I__4936\ : Span4Mux_h
    port map (
            O => \N__25651\,
            I => \N__25641\
        );

    \I__4935\ : Span4Mux_h
    port map (
            O => \N__25644\,
            I => \N__25638\
        );

    \I__4934\ : Odrv4
    port map (
            O => \N__25641\,
            I => \N_1709_0\
        );

    \I__4933\ : Odrv4
    port map (
            O => \N__25638\,
            I => \N_1709_0\
        );

    \I__4932\ : CEMux
    port map (
            O => \N__25633\,
            I => \N__25628\
        );

    \I__4931\ : CEMux
    port map (
            O => \N__25632\,
            I => \N__25625\
        );

    \I__4930\ : CEMux
    port map (
            O => \N__25631\,
            I => \N__25622\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__25628\,
            I => \N__25619\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__25625\,
            I => \N__25616\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__25622\,
            I => \N__25613\
        );

    \I__4926\ : Span4Mux_h
    port map (
            O => \N__25619\,
            I => \N__25610\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__25616\,
            I => \N__25605\
        );

    \I__4924\ : Span4Mux_h
    port map (
            O => \N__25613\,
            I => \N__25605\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__25610\,
            I => \N_1693_0\
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__25605\,
            I => \N_1693_0\
        );

    \I__4921\ : IoInMux
    port map (
            O => \N__25600\,
            I => \N__25597\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__25597\,
            I => \N__25594\
        );

    \I__4919\ : Span12Mux_s5_v
    port map (
            O => \N__25594\,
            I => \N__25591\
        );

    \I__4918\ : Odrv12
    port map (
            O => \N__25591\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI01JU6Z0Z_9\
        );

    \I__4917\ : CascadeMux
    port map (
            O => \N__25588\,
            I => \this_ppu.N_1269_cascade_\
        );

    \I__4916\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25582\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__25582\,
            I => \N__25579\
        );

    \I__4914\ : Span4Mux_v
    port map (
            O => \N__25579\,
            I => \N__25576\
        );

    \I__4913\ : Odrv4
    port map (
            O => \N__25576\,
            I => \this_ppu.N_1006_0\
        );

    \I__4912\ : CascadeMux
    port map (
            O => \N__25573\,
            I => \this_vga_signals.N_1264_cascade_\
        );

    \I__4911\ : InMux
    port map (
            O => \N__25570\,
            I => \N__25567\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__25567\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_4_1_0_x0\
        );

    \I__4909\ : CascadeMux
    port map (
            O => \N__25564\,
            I => \this_ppu.N_1301_cascade_\
        );

    \I__4908\ : InMux
    port map (
            O => \N__25561\,
            I => \N__25558\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__25558\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1_THRU_CO\
        );

    \I__4906\ : CascadeMux
    port map (
            O => \N__25555\,
            I => \N__25552\
        );

    \I__4905\ : InMux
    port map (
            O => \N__25552\,
            I => \N__25547\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__25551\,
            I => \N__25544\
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__25550\,
            I => \N__25541\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__25547\,
            I => \N__25538\
        );

    \I__4901\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25533\
        );

    \I__4900\ : InMux
    port map (
            O => \N__25541\,
            I => \N__25533\
        );

    \I__4899\ : Odrv4
    port map (
            O => \N__25538\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_6\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__25533\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_6\
        );

    \I__4897\ : InMux
    port map (
            O => \N__25528\,
            I => \N__25520\
        );

    \I__4896\ : InMux
    port map (
            O => \N__25527\,
            I => \N__25509\
        );

    \I__4895\ : InMux
    port map (
            O => \N__25526\,
            I => \N__25509\
        );

    \I__4894\ : InMux
    port map (
            O => \N__25525\,
            I => \N__25509\
        );

    \I__4893\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25509\
        );

    \I__4892\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25509\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__25520\,
            I => \N__25505\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__25509\,
            I => \N__25502\
        );

    \I__4889\ : InMux
    port map (
            O => \N__25508\,
            I => \N__25499\
        );

    \I__4888\ : Odrv4
    port map (
            O => \N__25505\,
            I => \this_ppu.N_1730_0\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__25502\,
            I => \this_ppu.N_1730_0\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__25499\,
            I => \this_ppu.N_1730_0\
        );

    \I__4885\ : InMux
    port map (
            O => \N__25492\,
            I => \N__25489\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__25489\,
            I => \N__25486\
        );

    \I__4883\ : Odrv4
    port map (
            O => \N__25486\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1_THRU_CO\
        );

    \I__4882\ : InMux
    port map (
            O => \N__25483\,
            I => \N__25475\
        );

    \I__4881\ : InMux
    port map (
            O => \N__25482\,
            I => \N__25464\
        );

    \I__4880\ : InMux
    port map (
            O => \N__25481\,
            I => \N__25464\
        );

    \I__4879\ : InMux
    port map (
            O => \N__25480\,
            I => \N__25464\
        );

    \I__4878\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25464\
        );

    \I__4877\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25464\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__25475\,
            I => \N__25459\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__25464\,
            I => \N__25456\
        );

    \I__4874\ : InMux
    port map (
            O => \N__25463\,
            I => \N__25453\
        );

    \I__4873\ : InMux
    port map (
            O => \N__25462\,
            I => \N__25450\
        );

    \I__4872\ : Odrv12
    port map (
            O => \N__25459\,
            I => \this_ppu.N_677_0\
        );

    \I__4871\ : Odrv4
    port map (
            O => \N__25456\,
            I => \this_ppu.N_677_0\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__25453\,
            I => \this_ppu.N_677_0\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__25450\,
            I => \this_ppu.N_677_0\
        );

    \I__4868\ : CascadeMux
    port map (
            O => \N__25441\,
            I => \N__25436\
        );

    \I__4867\ : CascadeMux
    port map (
            O => \N__25440\,
            I => \N__25433\
        );

    \I__4866\ : CascadeMux
    port map (
            O => \N__25439\,
            I => \N__25430\
        );

    \I__4865\ : InMux
    port map (
            O => \N__25436\,
            I => \N__25427\
        );

    \I__4864\ : InMux
    port map (
            O => \N__25433\,
            I => \N__25424\
        );

    \I__4863\ : InMux
    port map (
            O => \N__25430\,
            I => \N__25421\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__25427\,
            I => \N__25418\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__25424\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_4\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__25421\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_4\
        );

    \I__4859\ : Odrv12
    port map (
            O => \N__25418\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_4\
        );

    \I__4858\ : InMux
    port map (
            O => \N__25411\,
            I => \N__25408\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__25408\,
            I => \N__25405\
        );

    \I__4856\ : Span4Mux_v
    port map (
            O => \N__25405\,
            I => \N__25402\
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__25402\,
            I => \M_this_data_count_q_cry_6_THRU_CO\
        );

    \I__4854\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25396\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__25396\,
            I => \N__25393\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__25393\,
            I => \M_this_data_count_q_cry_8_THRU_CO\
        );

    \I__4851\ : InMux
    port map (
            O => \N__25390\,
            I => \N__25385\
        );

    \I__4850\ : CascadeMux
    port map (
            O => \N__25389\,
            I => \N__25382\
        );

    \I__4849\ : InMux
    port map (
            O => \N__25388\,
            I => \N__25379\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__25385\,
            I => \N__25376\
        );

    \I__4847\ : InMux
    port map (
            O => \N__25382\,
            I => \N__25373\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__25379\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__4845\ : Odrv4
    port map (
            O => \N__25376\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__25373\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__4843\ : CEMux
    port map (
            O => \N__25366\,
            I => \N__25362\
        );

    \I__4842\ : CEMux
    port map (
            O => \N__25365\,
            I => \N__25359\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__25362\,
            I => \N__25353\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__25359\,
            I => \N__25353\
        );

    \I__4839\ : CEMux
    port map (
            O => \N__25358\,
            I => \N__25350\
        );

    \I__4838\ : Span4Mux_v
    port map (
            O => \N__25353\,
            I => \N__25347\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__25350\,
            I => \N__25344\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__25347\,
            I => \N_231\
        );

    \I__4835\ : Odrv4
    port map (
            O => \N__25344\,
            I => \N_231\
        );

    \I__4834\ : InMux
    port map (
            O => \N__25339\,
            I => \N__25336\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__25336\,
            I => \N__25333\
        );

    \I__4832\ : Span4Mux_h
    port map (
            O => \N__25333\,
            I => \N__25330\
        );

    \I__4831\ : Odrv4
    port map (
            O => \N__25330\,
            I => \M_this_data_tmp_qZ0Z_2\
        );

    \I__4830\ : InMux
    port map (
            O => \N__25327\,
            I => \N__25324\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__25324\,
            I => \N__25321\
        );

    \I__4828\ : Span4Mux_h
    port map (
            O => \N__25321\,
            I => \N__25318\
        );

    \I__4827\ : Span4Mux_h
    port map (
            O => \N__25318\,
            I => \N__25315\
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__25315\,
            I => \M_this_oam_ram_write_data_2\
        );

    \I__4825\ : InMux
    port map (
            O => \N__25312\,
            I => \N__25307\
        );

    \I__4824\ : InMux
    port map (
            O => \N__25311\,
            I => \N__25304\
        );

    \I__4823\ : InMux
    port map (
            O => \N__25310\,
            I => \N__25301\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__25307\,
            I => \N__25298\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__25304\,
            I => \N__25295\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__25301\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_3\
        );

    \I__4819\ : Odrv12
    port map (
            O => \N__25298\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_3\
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__25295\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_3\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__25288\,
            I => \N__25285\
        );

    \I__4816\ : InMux
    port map (
            O => \N__25285\,
            I => \N__25282\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__25282\,
            I => \N__25279\
        );

    \I__4814\ : Span4Mux_v
    port map (
            O => \N__25279\,
            I => \N__25276\
        );

    \I__4813\ : Odrv4
    port map (
            O => \N__25276\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1_THRU_CO\
        );

    \I__4812\ : InMux
    port map (
            O => \N__25273\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1\
        );

    \I__4811\ : InMux
    port map (
            O => \N__25270\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1\
        );

    \I__4810\ : InMux
    port map (
            O => \N__25267\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1\
        );

    \I__4809\ : SRMux
    port map (
            O => \N__25264\,
            I => \N__25256\
        );

    \I__4808\ : SRMux
    port map (
            O => \N__25263\,
            I => \N__25252\
        );

    \I__4807\ : SRMux
    port map (
            O => \N__25262\,
            I => \N__25248\
        );

    \I__4806\ : SRMux
    port map (
            O => \N__25261\,
            I => \N__25244\
        );

    \I__4805\ : IoInMux
    port map (
            O => \N__25260\,
            I => \N__25240\
        );

    \I__4804\ : SRMux
    port map (
            O => \N__25259\,
            I => \N__25237\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__25256\,
            I => \N__25232\
        );

    \I__4802\ : SRMux
    port map (
            O => \N__25255\,
            I => \N__25229\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__25252\,
            I => \N__25224\
        );

    \I__4800\ : SRMux
    port map (
            O => \N__25251\,
            I => \N__25221\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__25248\,
            I => \N__25216\
        );

    \I__4798\ : SRMux
    port map (
            O => \N__25247\,
            I => \N__25213\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__25244\,
            I => \N__25210\
        );

    \I__4796\ : SRMux
    port map (
            O => \N__25243\,
            I => \N__25207\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__25240\,
            I => \N__25200\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__25237\,
            I => \N__25196\
        );

    \I__4793\ : SRMux
    port map (
            O => \N__25236\,
            I => \N__25193\
        );

    \I__4792\ : SRMux
    port map (
            O => \N__25235\,
            I => \N__25190\
        );

    \I__4791\ : Span4Mux_s3_v
    port map (
            O => \N__25232\,
            I => \N__25187\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__25229\,
            I => \N__25184\
        );

    \I__4789\ : SRMux
    port map (
            O => \N__25228\,
            I => \N__25181\
        );

    \I__4788\ : SRMux
    port map (
            O => \N__25227\,
            I => \N__25178\
        );

    \I__4787\ : Span4Mux_v
    port map (
            O => \N__25224\,
            I => \N__25171\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__25221\,
            I => \N__25171\
        );

    \I__4785\ : SRMux
    port map (
            O => \N__25220\,
            I => \N__25168\
        );

    \I__4784\ : SRMux
    port map (
            O => \N__25219\,
            I => \N__25165\
        );

    \I__4783\ : Span4Mux_v
    port map (
            O => \N__25216\,
            I => \N__25155\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__25213\,
            I => \N__25155\
        );

    \I__4781\ : Span4Mux_h
    port map (
            O => \N__25210\,
            I => \N__25155\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__25207\,
            I => \N__25155\
        );

    \I__4779\ : SRMux
    port map (
            O => \N__25206\,
            I => \N__25152\
        );

    \I__4778\ : SRMux
    port map (
            O => \N__25205\,
            I => \N__25149\
        );

    \I__4777\ : SRMux
    port map (
            O => \N__25204\,
            I => \N__25146\
        );

    \I__4776\ : SRMux
    port map (
            O => \N__25203\,
            I => \N__25143\
        );

    \I__4775\ : IoSpan4Mux
    port map (
            O => \N__25200\,
            I => \N__25139\
        );

    \I__4774\ : SRMux
    port map (
            O => \N__25199\,
            I => \N__25135\
        );

    \I__4773\ : Span4Mux_s3_v
    port map (
            O => \N__25196\,
            I => \N__25126\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__25193\,
            I => \N__25126\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__25190\,
            I => \N__25126\
        );

    \I__4770\ : Span4Mux_h
    port map (
            O => \N__25187\,
            I => \N__25117\
        );

    \I__4769\ : Span4Mux_s3_v
    port map (
            O => \N__25184\,
            I => \N__25117\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__25181\,
            I => \N__25117\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__25178\,
            I => \N__25117\
        );

    \I__4766\ : SRMux
    port map (
            O => \N__25177\,
            I => \N__25114\
        );

    \I__4765\ : SRMux
    port map (
            O => \N__25176\,
            I => \N__25111\
        );

    \I__4764\ : Span4Mux_v
    port map (
            O => \N__25171\,
            I => \N__25103\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__25168\,
            I => \N__25103\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__25165\,
            I => \N__25103\
        );

    \I__4761\ : SRMux
    port map (
            O => \N__25164\,
            I => \N__25100\
        );

    \I__4760\ : Span4Mux_v
    port map (
            O => \N__25155\,
            I => \N__25093\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__25152\,
            I => \N__25093\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__25149\,
            I => \N__25093\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__25146\,
            I => \N__25088\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__25143\,
            I => \N__25088\
        );

    \I__4755\ : SRMux
    port map (
            O => \N__25142\,
            I => \N__25085\
        );

    \I__4754\ : Span4Mux_s0_h
    port map (
            O => \N__25139\,
            I => \N__25080\
        );

    \I__4753\ : SRMux
    port map (
            O => \N__25138\,
            I => \N__25077\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__25135\,
            I => \N__25068\
        );

    \I__4751\ : SRMux
    port map (
            O => \N__25134\,
            I => \N__25065\
        );

    \I__4750\ : SRMux
    port map (
            O => \N__25133\,
            I => \N__25062\
        );

    \I__4749\ : Span4Mux_v
    port map (
            O => \N__25126\,
            I => \N__25050\
        );

    \I__4748\ : Span4Mux_v
    port map (
            O => \N__25117\,
            I => \N__25050\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__25114\,
            I => \N__25050\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__25111\,
            I => \N__25050\
        );

    \I__4745\ : SRMux
    port map (
            O => \N__25110\,
            I => \N__25047\
        );

    \I__4744\ : Span4Mux_v
    port map (
            O => \N__25103\,
            I => \N__25036\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__25100\,
            I => \N__25036\
        );

    \I__4742\ : Span4Mux_v
    port map (
            O => \N__25093\,
            I => \N__25036\
        );

    \I__4741\ : Span4Mux_v
    port map (
            O => \N__25088\,
            I => \N__25036\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__25085\,
            I => \N__25036\
        );

    \I__4739\ : SRMux
    port map (
            O => \N__25084\,
            I => \N__25033\
        );

    \I__4738\ : SRMux
    port map (
            O => \N__25083\,
            I => \N__25030\
        );

    \I__4737\ : Span4Mux_h
    port map (
            O => \N__25080\,
            I => \N__25025\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__25077\,
            I => \N__25025\
        );

    \I__4735\ : SRMux
    port map (
            O => \N__25076\,
            I => \N__25022\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__25075\,
            I => \N__25014\
        );

    \I__4733\ : CascadeMux
    port map (
            O => \N__25074\,
            I => \N__25010\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__25073\,
            I => \N__25006\
        );

    \I__4731\ : SRMux
    port map (
            O => \N__25072\,
            I => \N__25003\
        );

    \I__4730\ : SRMux
    port map (
            O => \N__25071\,
            I => \N__25000\
        );

    \I__4729\ : Span4Mux_s3_v
    port map (
            O => \N__25068\,
            I => \N__24992\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__25065\,
            I => \N__24992\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__25062\,
            I => \N__24992\
        );

    \I__4726\ : SRMux
    port map (
            O => \N__25061\,
            I => \N__24988\
        );

    \I__4725\ : SRMux
    port map (
            O => \N__25060\,
            I => \N__24983\
        );

    \I__4724\ : SRMux
    port map (
            O => \N__25059\,
            I => \N__24980\
        );

    \I__4723\ : Span4Mux_v
    port map (
            O => \N__25050\,
            I => \N__24971\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__25047\,
            I => \N__24971\
        );

    \I__4721\ : Span4Mux_v
    port map (
            O => \N__25036\,
            I => \N__24971\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__25033\,
            I => \N__24971\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__25030\,
            I => \N__24968\
        );

    \I__4718\ : Span4Mux_h
    port map (
            O => \N__25025\,
            I => \N__24965\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__25022\,
            I => \N__24962\
        );

    \I__4716\ : CascadeMux
    port map (
            O => \N__25021\,
            I => \N__24959\
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__25020\,
            I => \N__24955\
        );

    \I__4714\ : CascadeMux
    port map (
            O => \N__25019\,
            I => \N__24951\
        );

    \I__4713\ : CascadeMux
    port map (
            O => \N__25018\,
            I => \N__24947\
        );

    \I__4712\ : InMux
    port map (
            O => \N__25017\,
            I => \N__24934\
        );

    \I__4711\ : InMux
    port map (
            O => \N__25014\,
            I => \N__24934\
        );

    \I__4710\ : InMux
    port map (
            O => \N__25013\,
            I => \N__24934\
        );

    \I__4709\ : InMux
    port map (
            O => \N__25010\,
            I => \N__24934\
        );

    \I__4708\ : InMux
    port map (
            O => \N__25009\,
            I => \N__24934\
        );

    \I__4707\ : InMux
    port map (
            O => \N__25006\,
            I => \N__24934\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__25003\,
            I => \N__24930\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__25000\,
            I => \N__24927\
        );

    \I__4704\ : SRMux
    port map (
            O => \N__24999\,
            I => \N__24924\
        );

    \I__4703\ : Span4Mux_v
    port map (
            O => \N__24992\,
            I => \N__24920\
        );

    \I__4702\ : SRMux
    port map (
            O => \N__24991\,
            I => \N__24917\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__24988\,
            I => \N__24914\
        );

    \I__4700\ : SRMux
    port map (
            O => \N__24987\,
            I => \N__24911\
        );

    \I__4699\ : SRMux
    port map (
            O => \N__24986\,
            I => \N__24908\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__24983\,
            I => \N__24899\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__24980\,
            I => \N__24899\
        );

    \I__4696\ : Span4Mux_v
    port map (
            O => \N__24971\,
            I => \N__24899\
        );

    \I__4695\ : Span4Mux_h
    port map (
            O => \N__24968\,
            I => \N__24896\
        );

    \I__4694\ : Span4Mux_v
    port map (
            O => \N__24965\,
            I => \N__24891\
        );

    \I__4693\ : Span4Mux_h
    port map (
            O => \N__24962\,
            I => \N__24891\
        );

    \I__4692\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24871\
        );

    \I__4691\ : InMux
    port map (
            O => \N__24958\,
            I => \N__24871\
        );

    \I__4690\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24871\
        );

    \I__4689\ : InMux
    port map (
            O => \N__24954\,
            I => \N__24871\
        );

    \I__4688\ : InMux
    port map (
            O => \N__24951\,
            I => \N__24871\
        );

    \I__4687\ : InMux
    port map (
            O => \N__24950\,
            I => \N__24871\
        );

    \I__4686\ : InMux
    port map (
            O => \N__24947\,
            I => \N__24871\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__24934\,
            I => \N__24866\
        );

    \I__4684\ : InMux
    port map (
            O => \N__24933\,
            I => \N__24863\
        );

    \I__4683\ : Span4Mux_v
    port map (
            O => \N__24930\,
            I => \N__24856\
        );

    \I__4682\ : Span4Mux_v
    port map (
            O => \N__24927\,
            I => \N__24856\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__24924\,
            I => \N__24856\
        );

    \I__4680\ : SRMux
    port map (
            O => \N__24923\,
            I => \N__24853\
        );

    \I__4679\ : Span4Mux_h
    port map (
            O => \N__24920\,
            I => \N__24847\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__24917\,
            I => \N__24847\
        );

    \I__4677\ : Span4Mux_v
    port map (
            O => \N__24914\,
            I => \N__24840\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__24911\,
            I => \N__24840\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__24908\,
            I => \N__24840\
        );

    \I__4674\ : SRMux
    port map (
            O => \N__24907\,
            I => \N__24837\
        );

    \I__4673\ : SRMux
    port map (
            O => \N__24906\,
            I => \N__24834\
        );

    \I__4672\ : Span4Mux_v
    port map (
            O => \N__24899\,
            I => \N__24830\
        );

    \I__4671\ : Sp12to4
    port map (
            O => \N__24896\,
            I => \N__24825\
        );

    \I__4670\ : Sp12to4
    port map (
            O => \N__24891\,
            I => \N__24825\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__24890\,
            I => \N__24822\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__24889\,
            I => \N__24819\
        );

    \I__4667\ : CascadeMux
    port map (
            O => \N__24888\,
            I => \N__24816\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__24887\,
            I => \N__24813\
        );

    \I__4665\ : CascadeMux
    port map (
            O => \N__24886\,
            I => \N__24810\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__24871\,
            I => \N__24807\
        );

    \I__4663\ : SRMux
    port map (
            O => \N__24870\,
            I => \N__24804\
        );

    \I__4662\ : IoInMux
    port map (
            O => \N__24869\,
            I => \N__24801\
        );

    \I__4661\ : Span4Mux_v
    port map (
            O => \N__24866\,
            I => \N__24796\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__24863\,
            I => \N__24796\
        );

    \I__4659\ : Span4Mux_v
    port map (
            O => \N__24856\,
            I => \N__24791\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__24853\,
            I => \N__24791\
        );

    \I__4657\ : SRMux
    port map (
            O => \N__24852\,
            I => \N__24788\
        );

    \I__4656\ : Span4Mux_v
    port map (
            O => \N__24847\,
            I => \N__24779\
        );

    \I__4655\ : Span4Mux_v
    port map (
            O => \N__24840\,
            I => \N__24779\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__24837\,
            I => \N__24779\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__24834\,
            I => \N__24779\
        );

    \I__4652\ : SRMux
    port map (
            O => \N__24833\,
            I => \N__24776\
        );

    \I__4651\ : Sp12to4
    port map (
            O => \N__24830\,
            I => \N__24771\
        );

    \I__4650\ : Span12Mux_v
    port map (
            O => \N__24825\,
            I => \N__24771\
        );

    \I__4649\ : InMux
    port map (
            O => \N__24822\,
            I => \N__24766\
        );

    \I__4648\ : InMux
    port map (
            O => \N__24819\,
            I => \N__24766\
        );

    \I__4647\ : InMux
    port map (
            O => \N__24816\,
            I => \N__24759\
        );

    \I__4646\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24759\
        );

    \I__4645\ : InMux
    port map (
            O => \N__24810\,
            I => \N__24759\
        );

    \I__4644\ : Span4Mux_v
    port map (
            O => \N__24807\,
            I => \N__24756\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__24804\,
            I => \N__24753\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__24801\,
            I => \N__24750\
        );

    \I__4641\ : Span4Mux_h
    port map (
            O => \N__24796\,
            I => \N__24743\
        );

    \I__4640\ : Span4Mux_v
    port map (
            O => \N__24791\,
            I => \N__24743\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__24788\,
            I => \N__24743\
        );

    \I__4638\ : Span4Mux_v
    port map (
            O => \N__24779\,
            I => \N__24738\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__24776\,
            I => \N__24738\
        );

    \I__4636\ : Span12Mux_h
    port map (
            O => \N__24771\,
            I => \N__24729\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__24766\,
            I => \N__24729\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__24759\,
            I => \N__24729\
        );

    \I__4633\ : Sp12to4
    port map (
            O => \N__24756\,
            I => \N__24729\
        );

    \I__4632\ : Span4Mux_v
    port map (
            O => \N__24753\,
            I => \N__24726\
        );

    \I__4631\ : IoSpan4Mux
    port map (
            O => \N__24750\,
            I => \N__24723\
        );

    \I__4630\ : Span4Mux_h
    port map (
            O => \N__24743\,
            I => \N__24720\
        );

    \I__4629\ : Span4Mux_v
    port map (
            O => \N__24738\,
            I => \N__24717\
        );

    \I__4628\ : Span12Mux_h
    port map (
            O => \N__24729\,
            I => \N__24714\
        );

    \I__4627\ : Span4Mux_h
    port map (
            O => \N__24726\,
            I => \N__24707\
        );

    \I__4626\ : Span4Mux_s3_h
    port map (
            O => \N__24723\,
            I => \N__24707\
        );

    \I__4625\ : Span4Mux_h
    port map (
            O => \N__24720\,
            I => \N__24707\
        );

    \I__4624\ : Span4Mux_h
    port map (
            O => \N__24717\,
            I => \N__24704\
        );

    \I__4623\ : Odrv12
    port map (
            O => \N__24714\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4622\ : Odrv4
    port map (
            O => \N__24707\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4621\ : Odrv4
    port map (
            O => \N__24704\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4620\ : InMux
    port map (
            O => \N__24697\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1\
        );

    \I__4619\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24690\
        );

    \I__4618\ : InMux
    port map (
            O => \N__24693\,
            I => \N__24687\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__24690\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_7\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__24687\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_7\
        );

    \I__4615\ : CascadeMux
    port map (
            O => \N__24682\,
            I => \N__24671\
        );

    \I__4614\ : InMux
    port map (
            O => \N__24681\,
            I => \N__24661\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__24680\,
            I => \N__24658\
        );

    \I__4612\ : CascadeMux
    port map (
            O => \N__24679\,
            I => \N__24655\
        );

    \I__4611\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24652\
        );

    \I__4610\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24649\
        );

    \I__4609\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24644\
        );

    \I__4608\ : InMux
    port map (
            O => \N__24675\,
            I => \N__24644\
        );

    \I__4607\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24631\
        );

    \I__4606\ : InMux
    port map (
            O => \N__24671\,
            I => \N__24631\
        );

    \I__4605\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24631\
        );

    \I__4604\ : InMux
    port map (
            O => \N__24669\,
            I => \N__24631\
        );

    \I__4603\ : InMux
    port map (
            O => \N__24668\,
            I => \N__24631\
        );

    \I__4602\ : InMux
    port map (
            O => \N__24667\,
            I => \N__24631\
        );

    \I__4601\ : InMux
    port map (
            O => \N__24666\,
            I => \N__24628\
        );

    \I__4600\ : InMux
    port map (
            O => \N__24665\,
            I => \N__24625\
        );

    \I__4599\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24622\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__24661\,
            I => \N__24619\
        );

    \I__4597\ : InMux
    port map (
            O => \N__24658\,
            I => \N__24616\
        );

    \I__4596\ : InMux
    port map (
            O => \N__24655\,
            I => \N__24611\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__24652\,
            I => \N__24608\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__24649\,
            I => \N__24605\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__24644\,
            I => \N__24600\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__24631\,
            I => \N__24600\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__24628\,
            I => \N__24597\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__24625\,
            I => \N__24588\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__24622\,
            I => \N__24588\
        );

    \I__4588\ : Span4Mux_v
    port map (
            O => \N__24619\,
            I => \N__24588\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__24616\,
            I => \N__24588\
        );

    \I__4586\ : InMux
    port map (
            O => \N__24615\,
            I => \N__24583\
        );

    \I__4585\ : InMux
    port map (
            O => \N__24614\,
            I => \N__24583\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__24611\,
            I => \N__24577\
        );

    \I__4583\ : Span4Mux_v
    port map (
            O => \N__24608\,
            I => \N__24570\
        );

    \I__4582\ : Span4Mux_h
    port map (
            O => \N__24605\,
            I => \N__24570\
        );

    \I__4581\ : Span4Mux_h
    port map (
            O => \N__24600\,
            I => \N__24570\
        );

    \I__4580\ : Span4Mux_v
    port map (
            O => \N__24597\,
            I => \N__24562\
        );

    \I__4579\ : Span4Mux_v
    port map (
            O => \N__24588\,
            I => \N__24562\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__24583\,
            I => \N__24562\
        );

    \I__4577\ : InMux
    port map (
            O => \N__24582\,
            I => \N__24557\
        );

    \I__4576\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24557\
        );

    \I__4575\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24554\
        );

    \I__4574\ : Span4Mux_h
    port map (
            O => \N__24577\,
            I => \N__24551\
        );

    \I__4573\ : Span4Mux_h
    port map (
            O => \N__24570\,
            I => \N__24548\
        );

    \I__4572\ : InMux
    port map (
            O => \N__24569\,
            I => \N__24545\
        );

    \I__4571\ : Span4Mux_h
    port map (
            O => \N__24562\,
            I => \N__24542\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__24557\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__24554\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0\
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__24551\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0\
        );

    \I__4567\ : Odrv4
    port map (
            O => \N__24548\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__24545\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0\
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__24542\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0\
        );

    \I__4564\ : InMux
    port map (
            O => \N__24529\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_6_s1\
        );

    \I__4563\ : InMux
    port map (
            O => \N__24526\,
            I => \N__24523\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__24523\,
            I => \this_ppu.N_1205\
        );

    \I__4561\ : InMux
    port map (
            O => \N__24520\,
            I => \N__24517\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__24517\,
            I => \N__24514\
        );

    \I__4559\ : Odrv4
    port map (
            O => \N__24514\,
            I => \this_ppu.M_state_d30_i_i_o2_4\
        );

    \I__4558\ : InMux
    port map (
            O => \N__24511\,
            I => \N__24508\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__24508\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_THRU_CO\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__24505\,
            I => \N__24501\
        );

    \I__4555\ : InMux
    port map (
            O => \N__24504\,
            I => \N__24497\
        );

    \I__4554\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24492\
        );

    \I__4553\ : InMux
    port map (
            O => \N__24500\,
            I => \N__24492\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__24497\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_1\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__24492\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_1\
        );

    \I__4550\ : CascadeMux
    port map (
            O => \N__24487\,
            I => \N__24484\
        );

    \I__4549\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24481\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__24481\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1_THRU_CO\
        );

    \I__4547\ : CascadeMux
    port map (
            O => \N__24478\,
            I => \N__24475\
        );

    \I__4546\ : InMux
    port map (
            O => \N__24475\,
            I => \N__24470\
        );

    \I__4545\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24465\
        );

    \I__4544\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24465\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__24470\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_2\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__24465\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_2\
        );

    \I__4541\ : CascadeMux
    port map (
            O => \N__24460\,
            I => \N__24457\
        );

    \I__4540\ : InMux
    port map (
            O => \N__24457\,
            I => \N__24454\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__24454\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1_THRU_CO\
        );

    \I__4538\ : InMux
    port map (
            O => \N__24451\,
            I => \N__24446\
        );

    \I__4537\ : InMux
    port map (
            O => \N__24450\,
            I => \N__24441\
        );

    \I__4536\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24441\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__24446\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_5\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__24441\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_5\
        );

    \I__4533\ : InMux
    port map (
            O => \N__24436\,
            I => \N__24433\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__24433\,
            I => \this_ppu.M_state_d30_i_i_o2_3\
        );

    \I__4531\ : InMux
    port map (
            O => \N__24430\,
            I => \N__24425\
        );

    \I__4530\ : InMux
    port map (
            O => \N__24429\,
            I => \N__24417\
        );

    \I__4529\ : InMux
    port map (
            O => \N__24428\,
            I => \N__24417\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__24425\,
            I => \N__24414\
        );

    \I__4527\ : InMux
    port map (
            O => \N__24424\,
            I => \N__24411\
        );

    \I__4526\ : InMux
    port map (
            O => \N__24423\,
            I => \N__24408\
        );

    \I__4525\ : InMux
    port map (
            O => \N__24422\,
            I => \N__24405\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__24417\,
            I => \N__24402\
        );

    \I__4523\ : Span4Mux_v
    port map (
            O => \N__24414\,
            I => \N__24398\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__24411\,
            I => \N__24393\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__24408\,
            I => \N__24393\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__24405\,
            I => \N__24388\
        );

    \I__4519\ : Span4Mux_h
    port map (
            O => \N__24402\,
            I => \N__24388\
        );

    \I__4518\ : InMux
    port map (
            O => \N__24401\,
            I => \N__24385\
        );

    \I__4517\ : Span4Mux_v
    port map (
            O => \N__24398\,
            I => \N__24382\
        );

    \I__4516\ : Span4Mux_v
    port map (
            O => \N__24393\,
            I => \N__24377\
        );

    \I__4515\ : Span4Mux_h
    port map (
            O => \N__24388\,
            I => \N__24377\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__24385\,
            I => \N__24374\
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__24382\,
            I => \this_ppu.N_79_0\
        );

    \I__4512\ : Odrv4
    port map (
            O => \N__24377\,
            I => \this_ppu.N_79_0\
        );

    \I__4511\ : Odrv4
    port map (
            O => \N__24374\,
            I => \this_ppu.N_79_0\
        );

    \I__4510\ : CascadeMux
    port map (
            O => \N__24367\,
            I => \this_ppu.N_79_0_cascade_\
        );

    \I__4509\ : InMux
    port map (
            O => \N__24364\,
            I => \N__24361\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__24361\,
            I => \N__24358\
        );

    \I__4507\ : Odrv4
    port map (
            O => \N__24358\,
            I => \this_ppu.M_pixel_cnt_q_600_1\
        );

    \I__4506\ : CascadeMux
    port map (
            O => \N__24355\,
            I => \N__24352\
        );

    \I__4505\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24349\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__24349\,
            I => \N__24346\
        );

    \I__4503\ : Odrv4
    port map (
            O => \N__24346\,
            I => \this_ppu.un1_M_pixel_cnt_d_1_sqmuxa_0_i_0_0\
        );

    \I__4502\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24336\
        );

    \I__4501\ : InMux
    port map (
            O => \N__24342\,
            I => \N__24336\
        );

    \I__4500\ : InMux
    port map (
            O => \N__24341\,
            I => \N__24333\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__24336\,
            I => \N__24330\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__24333\,
            I => \N__24327\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__24330\,
            I => \N__24324\
        );

    \I__4496\ : Odrv4
    port map (
            O => \N__24327\,
            I => \this_ppu.N_999_0\
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__24324\,
            I => \this_ppu.N_999_0\
        );

    \I__4494\ : InMux
    port map (
            O => \N__24319\,
            I => \N__24315\
        );

    \I__4493\ : InMux
    port map (
            O => \N__24318\,
            I => \N__24312\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__24315\,
            I => \N__24308\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__24312\,
            I => \N__24305\
        );

    \I__4490\ : InMux
    port map (
            O => \N__24311\,
            I => \N__24302\
        );

    \I__4489\ : Span4Mux_v
    port map (
            O => \N__24308\,
            I => \N__24298\
        );

    \I__4488\ : Span4Mux_v
    port map (
            O => \N__24305\,
            I => \N__24295\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__24302\,
            I => \N__24292\
        );

    \I__4486\ : InMux
    port map (
            O => \N__24301\,
            I => \N__24289\
        );

    \I__4485\ : Span4Mux_h
    port map (
            O => \N__24298\,
            I => \N__24286\
        );

    \I__4484\ : Span4Mux_h
    port map (
            O => \N__24295\,
            I => \N__24283\
        );

    \I__4483\ : Sp12to4
    port map (
            O => \N__24292\,
            I => \N__24278\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__24289\,
            I => \N__24278\
        );

    \I__4481\ : Odrv4
    port map (
            O => \N__24286\,
            I => \this_ppu.N_838_0\
        );

    \I__4480\ : Odrv4
    port map (
            O => \N__24283\,
            I => \this_ppu.N_838_0\
        );

    \I__4479\ : Odrv12
    port map (
            O => \N__24278\,
            I => \this_ppu.N_838_0\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__24271\,
            I => \N__24267\
        );

    \I__4477\ : InMux
    port map (
            O => \N__24270\,
            I => \N__24264\
        );

    \I__4476\ : InMux
    port map (
            O => \N__24267\,
            I => \N__24260\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__24264\,
            I => \N__24257\
        );

    \I__4474\ : CascadeMux
    port map (
            O => \N__24263\,
            I => \N__24254\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__24260\,
            I => \N__24251\
        );

    \I__4472\ : Span4Mux_v
    port map (
            O => \N__24257\,
            I => \N__24247\
        );

    \I__4471\ : InMux
    port map (
            O => \N__24254\,
            I => \N__24244\
        );

    \I__4470\ : Span4Mux_h
    port map (
            O => \N__24251\,
            I => \N__24241\
        );

    \I__4469\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24238\
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__24247\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__24244\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__24241\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__24238\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__4464\ : InMux
    port map (
            O => \N__24229\,
            I => \N__24226\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__24226\,
            I => \this_ppu.N_1042_0\
        );

    \I__4462\ : CascadeMux
    port map (
            O => \N__24223\,
            I => \N__24215\
        );

    \I__4461\ : InMux
    port map (
            O => \N__24222\,
            I => \N__24212\
        );

    \I__4460\ : InMux
    port map (
            O => \N__24221\,
            I => \N__24209\
        );

    \I__4459\ : InMux
    port map (
            O => \N__24220\,
            I => \N__24206\
        );

    \I__4458\ : InMux
    port map (
            O => \N__24219\,
            I => \N__24201\
        );

    \I__4457\ : InMux
    port map (
            O => \N__24218\,
            I => \N__24201\
        );

    \I__4456\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24198\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__24212\,
            I => \N__24193\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__24209\,
            I => \N__24193\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__24206\,
            I => \this_ppu.M_state_qZ0Z_11\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__24201\,
            I => \this_ppu.M_state_qZ0Z_11\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__24198\,
            I => \this_ppu.M_state_qZ0Z_11\
        );

    \I__4450\ : Odrv12
    port map (
            O => \N__24193\,
            I => \this_ppu.M_state_qZ0Z_11\
        );

    \I__4449\ : CEMux
    port map (
            O => \N__24184\,
            I => \N__24168\
        );

    \I__4448\ : CascadeMux
    port map (
            O => \N__24183\,
            I => \N__24165\
        );

    \I__4447\ : InMux
    port map (
            O => \N__24182\,
            I => \N__24160\
        );

    \I__4446\ : InMux
    port map (
            O => \N__24181\,
            I => \N__24157\
        );

    \I__4445\ : InMux
    port map (
            O => \N__24180\,
            I => \N__24154\
        );

    \I__4444\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24149\
        );

    \I__4443\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24149\
        );

    \I__4442\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24146\
        );

    \I__4441\ : CascadeMux
    port map (
            O => \N__24176\,
            I => \N__24143\
        );

    \I__4440\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24125\
        );

    \I__4439\ : InMux
    port map (
            O => \N__24174\,
            I => \N__24125\
        );

    \I__4438\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24125\
        );

    \I__4437\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24125\
        );

    \I__4436\ : InMux
    port map (
            O => \N__24171\,
            I => \N__24122\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__24168\,
            I => \N__24119\
        );

    \I__4434\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24116\
        );

    \I__4433\ : CascadeMux
    port map (
            O => \N__24164\,
            I => \N__24110\
        );

    \I__4432\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24107\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__24160\,
            I => \N__24102\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__24157\,
            I => \N__24102\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__24154\,
            I => \N__24097\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__24149\,
            I => \N__24097\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__24146\,
            I => \N__24091\
        );

    \I__4426\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24088\
        );

    \I__4425\ : InMux
    port map (
            O => \N__24142\,
            I => \N__24085\
        );

    \I__4424\ : CEMux
    port map (
            O => \N__24141\,
            I => \N__24082\
        );

    \I__4423\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24078\
        );

    \I__4422\ : InMux
    port map (
            O => \N__24139\,
            I => \N__24075\
        );

    \I__4421\ : InMux
    port map (
            O => \N__24138\,
            I => \N__24070\
        );

    \I__4420\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24070\
        );

    \I__4419\ : InMux
    port map (
            O => \N__24136\,
            I => \N__24067\
        );

    \I__4418\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24064\
        );

    \I__4417\ : InMux
    port map (
            O => \N__24134\,
            I => \N__24061\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__24125\,
            I => \N__24056\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__24122\,
            I => \N__24056\
        );

    \I__4414\ : Span4Mux_h
    port map (
            O => \N__24119\,
            I => \N__24051\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__24116\,
            I => \N__24051\
        );

    \I__4412\ : InMux
    port map (
            O => \N__24115\,
            I => \N__24044\
        );

    \I__4411\ : InMux
    port map (
            O => \N__24114\,
            I => \N__24044\
        );

    \I__4410\ : InMux
    port map (
            O => \N__24113\,
            I => \N__24044\
        );

    \I__4409\ : InMux
    port map (
            O => \N__24110\,
            I => \N__24041\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__24107\,
            I => \N__24034\
        );

    \I__4407\ : Span4Mux_v
    port map (
            O => \N__24102\,
            I => \N__24034\
        );

    \I__4406\ : Span4Mux_h
    port map (
            O => \N__24097\,
            I => \N__24034\
        );

    \I__4405\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24031\
        );

    \I__4404\ : InMux
    port map (
            O => \N__24095\,
            I => \N__24026\
        );

    \I__4403\ : InMux
    port map (
            O => \N__24094\,
            I => \N__24026\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__24091\,
            I => \N__24023\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__24088\,
            I => \N__24018\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__24085\,
            I => \N__24018\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__24082\,
            I => \N__24013\
        );

    \I__4398\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24004\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__24078\,
            I => \N__24001\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__24075\,
            I => \N__23994\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__24070\,
            I => \N__23994\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__24067\,
            I => \N__23994\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__24064\,
            I => \N__23986\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__24061\,
            I => \N__23986\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__24056\,
            I => \N__23986\
        );

    \I__4390\ : Span4Mux_h
    port map (
            O => \N__24051\,
            I => \N__23977\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__24044\,
            I => \N__23977\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__24041\,
            I => \N__23977\
        );

    \I__4387\ : Span4Mux_h
    port map (
            O => \N__24034\,
            I => \N__23977\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__24031\,
            I => \N__23968\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__24026\,
            I => \N__23968\
        );

    \I__4384\ : Span4Mux_v
    port map (
            O => \N__24023\,
            I => \N__23968\
        );

    \I__4383\ : Span4Mux_h
    port map (
            O => \N__24018\,
            I => \N__23968\
        );

    \I__4382\ : InMux
    port map (
            O => \N__24017\,
            I => \N__23963\
        );

    \I__4381\ : InMux
    port map (
            O => \N__24016\,
            I => \N__23963\
        );

    \I__4380\ : Span4Mux_v
    port map (
            O => \N__24013\,
            I => \N__23960\
        );

    \I__4379\ : InMux
    port map (
            O => \N__24012\,
            I => \N__23957\
        );

    \I__4378\ : InMux
    port map (
            O => \N__24011\,
            I => \N__23946\
        );

    \I__4377\ : InMux
    port map (
            O => \N__24010\,
            I => \N__23946\
        );

    \I__4376\ : InMux
    port map (
            O => \N__24009\,
            I => \N__23946\
        );

    \I__4375\ : InMux
    port map (
            O => \N__24008\,
            I => \N__23946\
        );

    \I__4374\ : InMux
    port map (
            O => \N__24007\,
            I => \N__23946\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__24004\,
            I => \N__23939\
        );

    \I__4372\ : Span4Mux_v
    port map (
            O => \N__24001\,
            I => \N__23939\
        );

    \I__4371\ : Span4Mux_v
    port map (
            O => \N__23994\,
            I => \N__23939\
        );

    \I__4370\ : InMux
    port map (
            O => \N__23993\,
            I => \N__23936\
        );

    \I__4369\ : Span4Mux_v
    port map (
            O => \N__23986\,
            I => \N__23933\
        );

    \I__4368\ : Span4Mux_v
    port map (
            O => \N__23977\,
            I => \N__23930\
        );

    \I__4367\ : Span4Mux_h
    port map (
            O => \N__23968\,
            I => \N__23927\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__23963\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__23960\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__23957\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__23946\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4362\ : Odrv4
    port map (
            O => \N__23939\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__23936\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4360\ : Odrv4
    port map (
            O => \N__23933\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4359\ : Odrv4
    port map (
            O => \N__23930\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__23927\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__23908\,
            I => \this_ppu.N_1042_0_cascade_\
        );

    \I__4356\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23902\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__23902\,
            I => \N__23899\
        );

    \I__4354\ : Span4Mux_h
    port map (
            O => \N__23899\,
            I => \N__23896\
        );

    \I__4353\ : Sp12to4
    port map (
            O => \N__23896\,
            I => \N__23893\
        );

    \I__4352\ : Odrv12
    port map (
            O => \N__23893\,
            I => \this_ppu.un30_0_a2_i_0\
        );

    \I__4351\ : InMux
    port map (
            O => \N__23890\,
            I => \N__23887\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__23887\,
            I => \N__23882\
        );

    \I__4349\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23877\
        );

    \I__4348\ : InMux
    port map (
            O => \N__23885\,
            I => \N__23877\
        );

    \I__4347\ : Odrv4
    port map (
            O => \N__23882\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_0\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__23877\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_0\
        );

    \I__4345\ : InMux
    port map (
            O => \N__23872\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1\
        );

    \I__4344\ : InMux
    port map (
            O => \N__23869\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1\
        );

    \I__4343\ : InMux
    port map (
            O => \N__23866\,
            I => \N__23863\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__23863\,
            I => \N__23860\
        );

    \I__4341\ : Odrv12
    port map (
            O => \N__23860\,
            I => \this_vga_signals.g0_2\
        );

    \I__4340\ : CascadeMux
    port map (
            O => \N__23857\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_cascade_\
        );

    \I__4339\ : CascadeMux
    port map (
            O => \N__23854\,
            I => \N__23851\
        );

    \I__4338\ : InMux
    port map (
            O => \N__23851\,
            I => \N__23848\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__23848\,
            I => \N__23845\
        );

    \I__4336\ : Span4Mux_h
    port map (
            O => \N__23845\,
            I => \N__23842\
        );

    \I__4335\ : Span4Mux_h
    port map (
            O => \N__23842\,
            I => \N__23839\
        );

    \I__4334\ : Odrv4
    port map (
            O => \N__23839\,
            I => \M_this_vga_signals_address_7\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__23836\,
            I => \N__23832\
        );

    \I__4332\ : InMux
    port map (
            O => \N__23835\,
            I => \N__23829\
        );

    \I__4331\ : InMux
    port map (
            O => \N__23832\,
            I => \N__23826\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__23829\,
            I => \N__23823\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__23826\,
            I => \N__23819\
        );

    \I__4328\ : Span4Mux_v
    port map (
            O => \N__23823\,
            I => \N__23815\
        );

    \I__4327\ : InMux
    port map (
            O => \N__23822\,
            I => \N__23812\
        );

    \I__4326\ : Span4Mux_h
    port map (
            O => \N__23819\,
            I => \N__23809\
        );

    \I__4325\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23806\
        );

    \I__4324\ : Odrv4
    port map (
            O => \N__23815\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__23812\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__23809\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__23806\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__4320\ : InMux
    port map (
            O => \N__23797\,
            I => \N__23794\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__23794\,
            I => \N__23790\
        );

    \I__4318\ : InMux
    port map (
            O => \N__23793\,
            I => \N__23787\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__23790\,
            I => \N__23781\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__23787\,
            I => \N__23781\
        );

    \I__4315\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23778\
        );

    \I__4314\ : Odrv4
    port map (
            O => \N__23781\,
            I => \this_ppu.N_82_0\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__23778\,
            I => \this_ppu.N_82_0\
        );

    \I__4312\ : InMux
    port map (
            O => \N__23773\,
            I => \N__23766\
        );

    \I__4311\ : InMux
    port map (
            O => \N__23772\,
            I => \N__23757\
        );

    \I__4310\ : InMux
    port map (
            O => \N__23771\,
            I => \N__23757\
        );

    \I__4309\ : InMux
    port map (
            O => \N__23770\,
            I => \N__23757\
        );

    \I__4308\ : InMux
    port map (
            O => \N__23769\,
            I => \N__23757\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__23766\,
            I => \this_ppu.N_1659_0\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__23757\,
            I => \this_ppu.N_1659_0\
        );

    \I__4305\ : InMux
    port map (
            O => \N__23752\,
            I => \N__23746\
        );

    \I__4304\ : InMux
    port map (
            O => \N__23751\,
            I => \N__23743\
        );

    \I__4303\ : InMux
    port map (
            O => \N__23750\,
            I => \N__23740\
        );

    \I__4302\ : InMux
    port map (
            O => \N__23749\,
            I => \N__23737\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__23746\,
            I => \N__23733\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__23743\,
            I => \N__23730\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__23740\,
            I => \N__23727\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__23737\,
            I => \N__23724\
        );

    \I__4297\ : InMux
    port map (
            O => \N__23736\,
            I => \N__23721\
        );

    \I__4296\ : Span4Mux_v
    port map (
            O => \N__23733\,
            I => \N__23718\
        );

    \I__4295\ : Span4Mux_h
    port map (
            O => \N__23730\,
            I => \N__23715\
        );

    \I__4294\ : Span4Mux_h
    port map (
            O => \N__23727\,
            I => \N__23712\
        );

    \I__4293\ : Span4Mux_h
    port map (
            O => \N__23724\,
            I => \N__23709\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__23721\,
            I => \this_ppu.M_screen_y_qZ0Z_3\
        );

    \I__4291\ : Odrv4
    port map (
            O => \N__23718\,
            I => \this_ppu.M_screen_y_qZ0Z_3\
        );

    \I__4290\ : Odrv4
    port map (
            O => \N__23715\,
            I => \this_ppu.M_screen_y_qZ0Z_3\
        );

    \I__4289\ : Odrv4
    port map (
            O => \N__23712\,
            I => \this_ppu.M_screen_y_qZ0Z_3\
        );

    \I__4288\ : Odrv4
    port map (
            O => \N__23709\,
            I => \this_ppu.M_screen_y_qZ0Z_3\
        );

    \I__4287\ : CascadeMux
    port map (
            O => \N__23698\,
            I => \N__23694\
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__23697\,
            I => \N__23691\
        );

    \I__4285\ : InMux
    port map (
            O => \N__23694\,
            I => \N__23688\
        );

    \I__4284\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23685\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__23688\,
            I => \M_this_scroll_qZ0Z_3\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__23685\,
            I => \M_this_scroll_qZ0Z_3\
        );

    \I__4281\ : InMux
    port map (
            O => \N__23680\,
            I => \N__23677\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__23677\,
            I => \N__23674\
        );

    \I__4279\ : Odrv4
    port map (
            O => \N__23674\,
            I => \this_ppu.M_screen_y_q_esr_RNIF77F7Z0Z_3\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__23671\,
            I => \N__23668\
        );

    \I__4277\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23662\
        );

    \I__4276\ : InMux
    port map (
            O => \N__23667\,
            I => \N__23659\
        );

    \I__4275\ : CascadeMux
    port map (
            O => \N__23666\,
            I => \N__23654\
        );

    \I__4274\ : InMux
    port map (
            O => \N__23665\,
            I => \N__23650\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__23662\,
            I => \N__23647\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__23659\,
            I => \N__23644\
        );

    \I__4271\ : InMux
    port map (
            O => \N__23658\,
            I => \N__23639\
        );

    \I__4270\ : InMux
    port map (
            O => \N__23657\,
            I => \N__23639\
        );

    \I__4269\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23636\
        );

    \I__4268\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23633\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__23650\,
            I => \N__23628\
        );

    \I__4266\ : Span4Mux_h
    port map (
            O => \N__23647\,
            I => \N__23628\
        );

    \I__4265\ : Span4Mux_v
    port map (
            O => \N__23644\,
            I => \N__23625\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__23639\,
            I => \this_ppu.M_state_qZ0Z_9\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__23636\,
            I => \this_ppu.M_state_qZ0Z_9\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__23633\,
            I => \this_ppu.M_state_qZ0Z_9\
        );

    \I__4261\ : Odrv4
    port map (
            O => \N__23628\,
            I => \this_ppu.M_state_qZ0Z_9\
        );

    \I__4260\ : Odrv4
    port map (
            O => \N__23625\,
            I => \this_ppu.M_state_qZ0Z_9\
        );

    \I__4259\ : InMux
    port map (
            O => \N__23614\,
            I => \N__23606\
        );

    \I__4258\ : CascadeMux
    port map (
            O => \N__23613\,
            I => \N__23603\
        );

    \I__4257\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23597\
        );

    \I__4256\ : InMux
    port map (
            O => \N__23611\,
            I => \N__23597\
        );

    \I__4255\ : InMux
    port map (
            O => \N__23610\,
            I => \N__23593\
        );

    \I__4254\ : InMux
    port map (
            O => \N__23609\,
            I => \N__23590\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__23606\,
            I => \N__23587\
        );

    \I__4252\ : InMux
    port map (
            O => \N__23603\,
            I => \N__23584\
        );

    \I__4251\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23581\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__23597\,
            I => \N__23578\
        );

    \I__4249\ : InMux
    port map (
            O => \N__23596\,
            I => \N__23575\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__23593\,
            I => \N__23572\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__23590\,
            I => \N__23567\
        );

    \I__4246\ : Span4Mux_h
    port map (
            O => \N__23587\,
            I => \N__23567\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__23584\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__23581\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__23578\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__23575\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__4241\ : Odrv4
    port map (
            O => \N__23572\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__23567\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__4239\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23548\
        );

    \I__4238\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23548\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__23548\,
            I => \this_ppu.N_61_0\
        );

    \I__4236\ : CascadeMux
    port map (
            O => \N__23545\,
            I => \N__23542\
        );

    \I__4235\ : InMux
    port map (
            O => \N__23542\,
            I => \N__23539\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__23539\,
            I => \N__23536\
        );

    \I__4233\ : Span4Mux_v
    port map (
            O => \N__23536\,
            I => \N__23532\
        );

    \I__4232\ : CascadeMux
    port map (
            O => \N__23535\,
            I => \N__23529\
        );

    \I__4231\ : Span4Mux_h
    port map (
            O => \N__23532\,
            I => \N__23525\
        );

    \I__4230\ : InMux
    port map (
            O => \N__23529\,
            I => \N__23520\
        );

    \I__4229\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23520\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__23525\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__23520\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__23515\,
            I => \this_ppu.N_61_0_cascade_\
        );

    \I__4225\ : CascadeMux
    port map (
            O => \N__23512\,
            I => \N__23509\
        );

    \I__4224\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23506\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__23506\,
            I => \N__23503\
        );

    \I__4222\ : Span4Mux_h
    port map (
            O => \N__23503\,
            I => \N__23500\
        );

    \I__4221\ : Span4Mux_h
    port map (
            O => \N__23500\,
            I => \N__23494\
        );

    \I__4220\ : InMux
    port map (
            O => \N__23499\,
            I => \N__23487\
        );

    \I__4219\ : InMux
    port map (
            O => \N__23498\,
            I => \N__23487\
        );

    \I__4218\ : InMux
    port map (
            O => \N__23497\,
            I => \N__23487\
        );

    \I__4217\ : Odrv4
    port map (
            O => \N__23494\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__23487\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__4215\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23470\
        );

    \I__4214\ : InMux
    port map (
            O => \N__23481\,
            I => \N__23470\
        );

    \I__4213\ : InMux
    port map (
            O => \N__23480\,
            I => \N__23470\
        );

    \I__4212\ : InMux
    port map (
            O => \N__23479\,
            I => \N__23470\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__23470\,
            I => \this_ppu.un1_M_screen_x_q_c2\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__23467\,
            I => \N__23462\
        );

    \I__4209\ : InMux
    port map (
            O => \N__23466\,
            I => \N__23456\
        );

    \I__4208\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23456\
        );

    \I__4207\ : InMux
    port map (
            O => \N__23462\,
            I => \N__23450\
        );

    \I__4206\ : InMux
    port map (
            O => \N__23461\,
            I => \N__23447\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__23456\,
            I => \N__23444\
        );

    \I__4204\ : InMux
    port map (
            O => \N__23455\,
            I => \N__23437\
        );

    \I__4203\ : InMux
    port map (
            O => \N__23454\,
            I => \N__23437\
        );

    \I__4202\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23437\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23434\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__23447\,
            I => \this_ppu.offset_x\
        );

    \I__4199\ : Odrv4
    port map (
            O => \N__23444\,
            I => \this_ppu.offset_x\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__23437\,
            I => \this_ppu.offset_x\
        );

    \I__4197\ : Odrv4
    port map (
            O => \N__23434\,
            I => \this_ppu.offset_x\
        );

    \I__4196\ : InMux
    port map (
            O => \N__23425\,
            I => \N__23422\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__23422\,
            I => \N__23419\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__23419\,
            I => \this_ppu.un1_M_surface_x_q_c1\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__23416\,
            I => \N__23413\
        );

    \I__4192\ : CascadeBuf
    port map (
            O => \N__23413\,
            I => \N__23410\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__23410\,
            I => \N__23407\
        );

    \I__4190\ : InMux
    port map (
            O => \N__23407\,
            I => \N__23404\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__23404\,
            I => \N__23401\
        );

    \I__4188\ : Sp12to4
    port map (
            O => \N__23401\,
            I => \N__23394\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__23400\,
            I => \N__23391\
        );

    \I__4186\ : InMux
    port map (
            O => \N__23399\,
            I => \N__23385\
        );

    \I__4185\ : InMux
    port map (
            O => \N__23398\,
            I => \N__23385\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__23397\,
            I => \N__23382\
        );

    \I__4183\ : Span12Mux_s7_v
    port map (
            O => \N__23394\,
            I => \N__23379\
        );

    \I__4182\ : InMux
    port map (
            O => \N__23391\,
            I => \N__23376\
        );

    \I__4181\ : InMux
    port map (
            O => \N__23390\,
            I => \N__23373\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__23385\,
            I => \N__23370\
        );

    \I__4179\ : InMux
    port map (
            O => \N__23382\,
            I => \N__23367\
        );

    \I__4178\ : Span12Mux_h
    port map (
            O => \N__23379\,
            I => \N__23364\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__23376\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__23373\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__23370\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__23367\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__4173\ : Odrv12
    port map (
            O => \N__23364\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__23353\,
            I => \N__23350\
        );

    \I__4171\ : InMux
    port map (
            O => \N__23350\,
            I => \N__23347\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__23347\,
            I => \N__23340\
        );

    \I__4169\ : InMux
    port map (
            O => \N__23346\,
            I => \N__23337\
        );

    \I__4168\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23330\
        );

    \I__4167\ : InMux
    port map (
            O => \N__23344\,
            I => \N__23330\
        );

    \I__4166\ : InMux
    port map (
            O => \N__23343\,
            I => \N__23330\
        );

    \I__4165\ : Span4Mux_v
    port map (
            O => \N__23340\,
            I => \N__23327\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__23337\,
            I => \this_ppu.M_surface_x_qZ0Z_2\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__23330\,
            I => \this_ppu.M_surface_x_qZ0Z_2\
        );

    \I__4162\ : Odrv4
    port map (
            O => \N__23327\,
            I => \this_ppu.M_surface_x_qZ0Z_2\
        );

    \I__4161\ : CascadeMux
    port map (
            O => \N__23320\,
            I => \this_ppu.un1_M_surface_x_q_c1_cascade_\
        );

    \I__4160\ : CascadeMux
    port map (
            O => \N__23317\,
            I => \N__23313\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__23316\,
            I => \N__23307\
        );

    \I__4158\ : InMux
    port map (
            O => \N__23313\,
            I => \N__23304\
        );

    \I__4157\ : InMux
    port map (
            O => \N__23312\,
            I => \N__23301\
        );

    \I__4156\ : InMux
    port map (
            O => \N__23311\,
            I => \N__23296\
        );

    \I__4155\ : InMux
    port map (
            O => \N__23310\,
            I => \N__23296\
        );

    \I__4154\ : InMux
    port map (
            O => \N__23307\,
            I => \N__23293\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__23304\,
            I => \N__23290\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__23301\,
            I => \N__23285\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__23296\,
            I => \N__23285\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__23293\,
            I => \N__23282\
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__23290\,
            I => \this_ppu.M_surface_x_qZ0Z_1\
        );

    \I__4148\ : Odrv4
    port map (
            O => \N__23285\,
            I => \this_ppu.M_surface_x_qZ0Z_1\
        );

    \I__4147\ : Odrv4
    port map (
            O => \N__23282\,
            I => \this_ppu.M_surface_x_qZ0Z_1\
        );

    \I__4146\ : InMux
    port map (
            O => \N__23275\,
            I => \N__23272\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__23272\,
            I => \N__23268\
        );

    \I__4144\ : InMux
    port map (
            O => \N__23271\,
            I => \N__23265\
        );

    \I__4143\ : Span4Mux_v
    port map (
            O => \N__23268\,
            I => \N__23262\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__23265\,
            I => \N__23259\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__23262\,
            I => \this_ppu.un1_M_surface_x_q_c4\
        );

    \I__4140\ : Odrv12
    port map (
            O => \N__23259\,
            I => \this_ppu.un1_M_surface_x_q_c4\
        );

    \I__4139\ : InMux
    port map (
            O => \N__23254\,
            I => \N__23251\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23246\
        );

    \I__4137\ : InMux
    port map (
            O => \N__23250\,
            I => \N__23243\
        );

    \I__4136\ : CascadeMux
    port map (
            O => \N__23249\,
            I => \N__23239\
        );

    \I__4135\ : Span4Mux_v
    port map (
            O => \N__23246\,
            I => \N__23234\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__23243\,
            I => \N__23234\
        );

    \I__4133\ : InMux
    port map (
            O => \N__23242\,
            I => \N__23231\
        );

    \I__4132\ : InMux
    port map (
            O => \N__23239\,
            I => \N__23228\
        );

    \I__4131\ : Span4Mux_h
    port map (
            O => \N__23234\,
            I => \N__23223\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__23231\,
            I => \N__23223\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__23228\,
            I => \N__23219\
        );

    \I__4128\ : Span4Mux_h
    port map (
            O => \N__23223\,
            I => \N__23216\
        );

    \I__4127\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23213\
        );

    \I__4126\ : Span4Mux_h
    port map (
            O => \N__23219\,
            I => \N__23210\
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__23216\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__23213\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__4123\ : Odrv4
    port map (
            O => \N__23210\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__4122\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23197\
        );

    \I__4121\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23194\
        );

    \I__4120\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23191\
        );

    \I__4119\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23188\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__23197\,
            I => \this_ppu.M_state_qZ0Z_10\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__23194\,
            I => \this_ppu.M_state_qZ0Z_10\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__23191\,
            I => \this_ppu.M_state_qZ0Z_10\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__23188\,
            I => \this_ppu.M_state_qZ0Z_10\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__23179\,
            I => \N__23176\
        );

    \I__4113\ : InMux
    port map (
            O => \N__23176\,
            I => \N__23173\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__23173\,
            I => \N__23167\
        );

    \I__4111\ : InMux
    port map (
            O => \N__23172\,
            I => \N__23163\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__23171\,
            I => \N__23160\
        );

    \I__4109\ : CascadeMux
    port map (
            O => \N__23170\,
            I => \N__23157\
        );

    \I__4108\ : Span4Mux_h
    port map (
            O => \N__23167\,
            I => \N__23153\
        );

    \I__4107\ : InMux
    port map (
            O => \N__23166\,
            I => \N__23150\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__23163\,
            I => \N__23147\
        );

    \I__4105\ : InMux
    port map (
            O => \N__23160\,
            I => \N__23140\
        );

    \I__4104\ : InMux
    port map (
            O => \N__23157\,
            I => \N__23140\
        );

    \I__4103\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23140\
        );

    \I__4102\ : Span4Mux_h
    port map (
            O => \N__23153\,
            I => \N__23133\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__23150\,
            I => \N__23133\
        );

    \I__4100\ : Span4Mux_h
    port map (
            O => \N__23147\,
            I => \N__23133\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__23140\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__23133\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__23128\,
            I => \this_ppu.N_798_0_cascade_\
        );

    \I__4096\ : InMux
    port map (
            O => \N__23125\,
            I => \N__23122\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__23122\,
            I => \N__23119\
        );

    \I__4094\ : Span12Mux_h
    port map (
            O => \N__23119\,
            I => \N__23116\
        );

    \I__4093\ : Odrv12
    port map (
            O => \N__23116\,
            I => \M_this_ppu_vram_data_0\
        );

    \I__4092\ : InMux
    port map (
            O => \N__23113\,
            I => \N__23108\
        );

    \I__4091\ : InMux
    port map (
            O => \N__23112\,
            I => \N__23105\
        );

    \I__4090\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23102\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__23108\,
            I => \N__23099\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__23105\,
            I => \N__23096\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__23102\,
            I => \N__23093\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__23099\,
            I => \N__23088\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__23096\,
            I => \N__23088\
        );

    \I__4084\ : Odrv4
    port map (
            O => \N__23093\,
            I => \this_ppu.N_1182_1\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__23088\,
            I => \this_ppu.N_1182_1\
        );

    \I__4082\ : CascadeMux
    port map (
            O => \N__23083\,
            I => \N__23078\
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__23082\,
            I => \N__23075\
        );

    \I__4080\ : InMux
    port map (
            O => \N__23081\,
            I => \N__23068\
        );

    \I__4079\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23068\
        );

    \I__4078\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23065\
        );

    \I__4077\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23061\
        );

    \I__4076\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23058\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__23068\,
            I => \N__23055\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__23065\,
            I => \N__23052\
        );

    \I__4073\ : InMux
    port map (
            O => \N__23064\,
            I => \N__23049\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__23061\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__23058\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4070\ : Odrv4
    port map (
            O => \N__23055\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4069\ : Odrv4
    port map (
            O => \N__23052\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__23049\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4067\ : CascadeMux
    port map (
            O => \N__23038\,
            I => \this_vga_signals.M_lcounter_q_e_1_0_cascade_\
        );

    \I__4066\ : CEMux
    port map (
            O => \N__23035\,
            I => \N__23032\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__23032\,
            I => \N__23029\
        );

    \I__4064\ : Span4Mux_h
    port map (
            O => \N__23029\,
            I => \N__23026\
        );

    \I__4063\ : Span4Mux_h
    port map (
            O => \N__23026\,
            I => \N__23023\
        );

    \I__4062\ : Span4Mux_v
    port map (
            O => \N__23023\,
            I => \N__23020\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__23020\,
            I => \N_26\
        );

    \I__4060\ : InMux
    port map (
            O => \N__23017\,
            I => \N__23014\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__23014\,
            I => \this_ppu.N_1198\
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__23011\,
            I => \this_ppu.N_1198_cascade_\
        );

    \I__4057\ : CascadeMux
    port map (
            O => \N__23008\,
            I => \N__23005\
        );

    \I__4056\ : CascadeBuf
    port map (
            O => \N__23005\,
            I => \N__23001\
        );

    \I__4055\ : CascadeMux
    port map (
            O => \N__23004\,
            I => \N__22998\
        );

    \I__4054\ : CascadeMux
    port map (
            O => \N__23001\,
            I => \N__22994\
        );

    \I__4053\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22991\
        );

    \I__4052\ : CascadeMux
    port map (
            O => \N__22997\,
            I => \N__22988\
        );

    \I__4051\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22983\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__22991\,
            I => \N__22980\
        );

    \I__4049\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22977\
        );

    \I__4048\ : InMux
    port map (
            O => \N__22987\,
            I => \N__22974\
        );

    \I__4047\ : InMux
    port map (
            O => \N__22986\,
            I => \N__22971\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__22983\,
            I => \N__22968\
        );

    \I__4045\ : Span4Mux_h
    port map (
            O => \N__22980\,
            I => \N__22964\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__22977\,
            I => \N__22961\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__22974\,
            I => \N__22956\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__22971\,
            I => \N__22956\
        );

    \I__4041\ : Span12Mux_s2_v
    port map (
            O => \N__22968\,
            I => \N__22953\
        );

    \I__4040\ : InMux
    port map (
            O => \N__22967\,
            I => \N__22950\
        );

    \I__4039\ : Span4Mux_v
    port map (
            O => \N__22964\,
            I => \N__22947\
        );

    \I__4038\ : Span4Mux_h
    port map (
            O => \N__22961\,
            I => \N__22944\
        );

    \I__4037\ : Span12Mux_h
    port map (
            O => \N__22956\,
            I => \N__22939\
        );

    \I__4036\ : Span12Mux_h
    port map (
            O => \N__22953\,
            I => \N__22939\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__22950\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4034\ : Odrv4
    port map (
            O => \N__22947\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__22944\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4032\ : Odrv12
    port map (
            O => \N__22939\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4031\ : CascadeMux
    port map (
            O => \N__22930\,
            I => \this_ppu.un1_M_surface_x_q_c2_cascade_\
        );

    \I__4030\ : CascadeMux
    port map (
            O => \N__22927\,
            I => \this_ppu.un1_M_surface_x_q_c5_cascade_\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__22924\,
            I => \N__22921\
        );

    \I__4028\ : CascadeBuf
    port map (
            O => \N__22921\,
            I => \N__22918\
        );

    \I__4027\ : CascadeMux
    port map (
            O => \N__22918\,
            I => \N__22915\
        );

    \I__4026\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22911\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__22914\,
            I => \N__22908\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__22911\,
            I => \N__22905\
        );

    \I__4023\ : InMux
    port map (
            O => \N__22908\,
            I => \N__22901\
        );

    \I__4022\ : Span4Mux_s2_v
    port map (
            O => \N__22905\,
            I => \N__22898\
        );

    \I__4021\ : InMux
    port map (
            O => \N__22904\,
            I => \N__22895\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__22901\,
            I => \N__22892\
        );

    \I__4019\ : Sp12to4
    port map (
            O => \N__22898\,
            I => \N__22889\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__22895\,
            I => \N__22882\
        );

    \I__4017\ : Span4Mux_v
    port map (
            O => \N__22892\,
            I => \N__22882\
        );

    \I__4016\ : Span12Mux_h
    port map (
            O => \N__22889\,
            I => \N__22879\
        );

    \I__4015\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22876\
        );

    \I__4014\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22873\
        );

    \I__4013\ : Span4Mux_h
    port map (
            O => \N__22882\,
            I => \N__22870\
        );

    \I__4012\ : Span12Mux_v
    port map (
            O => \N__22879\,
            I => \N__22867\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__22876\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__22873\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__4009\ : Odrv4
    port map (
            O => \N__22870\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__4008\ : Odrv12
    port map (
            O => \N__22867\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__4007\ : InMux
    port map (
            O => \N__22858\,
            I => \N__22855\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__22855\,
            I => \this_ppu.un1_M_surface_x_q_c2\
        );

    \I__4005\ : InMux
    port map (
            O => \N__22852\,
            I => \N__22849\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__22849\,
            I => \N__22846\
        );

    \I__4003\ : Odrv4
    port map (
            O => \N__22846\,
            I => \M_this_data_count_q_s_13\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__22843\,
            I => \N__22839\
        );

    \I__4001\ : InMux
    port map (
            O => \N__22842\,
            I => \N__22835\
        );

    \I__4000\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22830\
        );

    \I__3999\ : InMux
    port map (
            O => \N__22838\,
            I => \N__22830\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__22835\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__22830\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__3996\ : InMux
    port map (
            O => \N__22825\,
            I => \N__22820\
        );

    \I__3995\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22815\
        );

    \I__3994\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22815\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__22820\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__22815\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__3991\ : CascadeMux
    port map (
            O => \N__22810\,
            I => \N__22806\
        );

    \I__3990\ : InMux
    port map (
            O => \N__22809\,
            I => \N__22803\
        );

    \I__3989\ : InMux
    port map (
            O => \N__22806\,
            I => \N__22800\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__22803\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__22800\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__3986\ : InMux
    port map (
            O => \N__22795\,
            I => \N__22791\
        );

    \I__3985\ : InMux
    port map (
            O => \N__22794\,
            I => \N__22788\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__22791\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__22788\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__3982\ : InMux
    port map (
            O => \N__22783\,
            I => \N__22780\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__22780\,
            I => \M_this_data_count_q_s_8\
        );

    \I__3980\ : InMux
    port map (
            O => \N__22777\,
            I => \N__22773\
        );

    \I__3979\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22770\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__22773\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__22770\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__3976\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22760\
        );

    \I__3975\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22757\
        );

    \I__3974\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22754\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__22760\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__22757\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__22754\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__22747\,
            I => \N__22743\
        );

    \I__3969\ : InMux
    port map (
            O => \N__22746\,
            I => \N__22739\
        );

    \I__3968\ : InMux
    port map (
            O => \N__22743\,
            I => \N__22736\
        );

    \I__3967\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22733\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__22739\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__22736\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__22733\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__3963\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22723\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__22723\,
            I => \un1_M_this_oam_address_q_c6\
        );

    \I__3961\ : InMux
    port map (
            O => \N__22720\,
            I => \N__22717\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__22717\,
            I => \N__22714\
        );

    \I__3959\ : Span12Mux_h
    port map (
            O => \N__22714\,
            I => \N__22711\
        );

    \I__3958\ : Odrv12
    port map (
            O => \N__22711\,
            I => \this_vga_signals.g0_1\
        );

    \I__3957\ : InMux
    port map (
            O => \N__22708\,
            I => \N__22704\
        );

    \I__3956\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22701\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__22704\,
            I => \N__22698\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__22701\,
            I => \this_vga_signals.N_3_0\
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__22698\,
            I => \this_vga_signals.N_3_0\
        );

    \I__3952\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22690\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__22690\,
            I => \N__22687\
        );

    \I__3950\ : Span4Mux_h
    port map (
            O => \N__22687\,
            I => \N__22683\
        );

    \I__3949\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22680\
        );

    \I__3948\ : Span4Mux_v
    port map (
            O => \N__22683\,
            I => \N__22677\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__22680\,
            I => \N__22674\
        );

    \I__3946\ : Odrv4
    port map (
            O => \N__22677\,
            I => \this_vga_signals.M_pcounter_q_i_2_1\
        );

    \I__3945\ : Odrv12
    port map (
            O => \N__22674\,
            I => \this_vga_signals.M_pcounter_q_i_2_1\
        );

    \I__3944\ : InMux
    port map (
            O => \N__22669\,
            I => \N__22666\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__22666\,
            I => \N__22663\
        );

    \I__3942\ : Span12Mux_v
    port map (
            O => \N__22663\,
            I => \N__22660\
        );

    \I__3941\ : Odrv12
    port map (
            O => \N__22660\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_CO\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__22657\,
            I => \N__22654\
        );

    \I__3939\ : CascadeBuf
    port map (
            O => \N__22654\,
            I => \N__22650\
        );

    \I__3938\ : CascadeMux
    port map (
            O => \N__22653\,
            I => \N__22647\
        );

    \I__3937\ : CascadeMux
    port map (
            O => \N__22650\,
            I => \N__22644\
        );

    \I__3936\ : InMux
    port map (
            O => \N__22647\,
            I => \N__22640\
        );

    \I__3935\ : InMux
    port map (
            O => \N__22644\,
            I => \N__22637\
        );

    \I__3934\ : CascadeMux
    port map (
            O => \N__22643\,
            I => \N__22633\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__22640\,
            I => \N__22630\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__22637\,
            I => \N__22627\
        );

    \I__3931\ : CascadeMux
    port map (
            O => \N__22636\,
            I => \N__22624\
        );

    \I__3930\ : InMux
    port map (
            O => \N__22633\,
            I => \N__22621\
        );

    \I__3929\ : Span4Mux_h
    port map (
            O => \N__22630\,
            I => \N__22618\
        );

    \I__3928\ : Span4Mux_h
    port map (
            O => \N__22627\,
            I => \N__22615\
        );

    \I__3927\ : InMux
    port map (
            O => \N__22624\,
            I => \N__22612\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__22621\,
            I => \N__22609\
        );

    \I__3925\ : Span4Mux_h
    port map (
            O => \N__22618\,
            I => \N__22606\
        );

    \I__3924\ : Span4Mux_h
    port map (
            O => \N__22615\,
            I => \N__22603\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__22612\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_2\
        );

    \I__3922\ : Odrv12
    port map (
            O => \N__22609\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_2\
        );

    \I__3921\ : Odrv4
    port map (
            O => \N__22606\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_2\
        );

    \I__3920\ : Odrv4
    port map (
            O => \N__22603\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_2\
        );

    \I__3919\ : InMux
    port map (
            O => \N__22594\,
            I => \N__22591\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__22591\,
            I => \M_this_data_count_q_cry_0_THRU_CO\
        );

    \I__3917\ : InMux
    port map (
            O => \N__22588\,
            I => \N__22583\
        );

    \I__3916\ : InMux
    port map (
            O => \N__22587\,
            I => \N__22578\
        );

    \I__3915\ : InMux
    port map (
            O => \N__22586\,
            I => \N__22578\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__22583\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__22578\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__3912\ : InMux
    port map (
            O => \N__22573\,
            I => \N__22570\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__22570\,
            I => \M_this_data_count_q_cry_1_THRU_CO\
        );

    \I__3910\ : CascadeMux
    port map (
            O => \N__22567\,
            I => \N__22564\
        );

    \I__3909\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22559\
        );

    \I__3908\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22554\
        );

    \I__3907\ : InMux
    port map (
            O => \N__22562\,
            I => \N__22554\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__22559\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__22554\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__3904\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22546\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__22546\,
            I => \M_this_data_count_q_cry_2_THRU_CO\
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__22543\,
            I => \N__22538\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__22542\,
            I => \N__22535\
        );

    \I__3900\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22532\
        );

    \I__3899\ : InMux
    port map (
            O => \N__22538\,
            I => \N__22527\
        );

    \I__3898\ : InMux
    port map (
            O => \N__22535\,
            I => \N__22527\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__22532\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__22527\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__3895\ : InMux
    port map (
            O => \N__22522\,
            I => \N__22519\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__22519\,
            I => \M_this_data_count_q_cry_3_THRU_CO\
        );

    \I__3893\ : InMux
    port map (
            O => \N__22516\,
            I => \N__22513\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__22513\,
            I => \M_this_data_count_q_cry_4_THRU_CO\
        );

    \I__3891\ : InMux
    port map (
            O => \N__22510\,
            I => \N__22507\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__22507\,
            I => \M_this_data_count_q_cry_5_THRU_CO\
        );

    \I__3889\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22501\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__22501\,
            I => \M_this_data_count_q_cry_10_THRU_CO\
        );

    \I__3887\ : InMux
    port map (
            O => \N__22498\,
            I => \N__22495\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__22495\,
            I => \N__22492\
        );

    \I__3885\ : Odrv4
    port map (
            O => \N__22492\,
            I => \M_this_data_count_q_s_10\
        );

    \I__3884\ : InMux
    port map (
            O => \N__22489\,
            I => \N__22486\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__22486\,
            I => \M_this_data_count_q_cry_11_THRU_CO\
        );

    \I__3882\ : CascadeMux
    port map (
            O => \N__22483\,
            I => \N__22480\
        );

    \I__3881\ : InMux
    port map (
            O => \N__22480\,
            I => \N__22477\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__22477\,
            I => \M_this_scroll_qZ0Z_2\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__22474\,
            I => \N__22471\
        );

    \I__3878\ : InMux
    port map (
            O => \N__22471\,
            I => \N__22467\
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__22470\,
            I => \N__22464\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__22467\,
            I => \N__22461\
        );

    \I__3875\ : InMux
    port map (
            O => \N__22464\,
            I => \N__22458\
        );

    \I__3874\ : Span4Mux_h
    port map (
            O => \N__22461\,
            I => \N__22455\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__22458\,
            I => \N__22452\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__22455\,
            I => \M_this_scroll_qZ0Z_4\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__22452\,
            I => \M_this_scroll_qZ0Z_4\
        );

    \I__3870\ : InMux
    port map (
            O => \N__22447\,
            I => \N__22444\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__22444\,
            I => \M_this_scroll_qZ0Z_7\
        );

    \I__3868\ : IoInMux
    port map (
            O => \N__22441\,
            I => \N__22438\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__22438\,
            I => \N__22435\
        );

    \I__3866\ : Span12Mux_s1_v
    port map (
            O => \N__22435\,
            I => \N__22432\
        );

    \I__3865\ : Span12Mux_h
    port map (
            O => \N__22432\,
            I => \N__22429\
        );

    \I__3864\ : Odrv12
    port map (
            O => \N__22429\,
            I => this_vga_signals_vsync_1_i
        );

    \I__3863\ : InMux
    port map (
            O => \N__22426\,
            I => \N__22421\
        );

    \I__3862\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22416\
        );

    \I__3861\ : InMux
    port map (
            O => \N__22424\,
            I => \N__22416\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__22421\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__22416\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__22411\,
            I => \N__22408\
        );

    \I__3857\ : InMux
    port map (
            O => \N__22408\,
            I => \N__22405\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__22405\,
            I => \N__22398\
        );

    \I__3855\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22395\
        );

    \I__3854\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22391\
        );

    \I__3853\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22388\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__22401\,
            I => \N__22385\
        );

    \I__3851\ : Span4Mux_v
    port map (
            O => \N__22398\,
            I => \N__22381\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__22395\,
            I => \N__22378\
        );

    \I__3849\ : InMux
    port map (
            O => \N__22394\,
            I => \N__22375\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__22391\,
            I => \N__22370\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__22388\,
            I => \N__22370\
        );

    \I__3846\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22367\
        );

    \I__3845\ : InMux
    port map (
            O => \N__22384\,
            I => \N__22364\
        );

    \I__3844\ : Span4Mux_h
    port map (
            O => \N__22381\,
            I => \N__22361\
        );

    \I__3843\ : Span4Mux_v
    port map (
            O => \N__22378\,
            I => \N__22354\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__22375\,
            I => \N__22354\
        );

    \I__3841\ : Span4Mux_v
    port map (
            O => \N__22370\,
            I => \N__22354\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__22367\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__22364\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__22361\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__22354\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__3836\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22342\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__22342\,
            I => \this_ppu.M_screen_y_q_RNIQ9FQ6Z0Z_0\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__22339\,
            I => \this_ppu.un1_M_screen_x_q_c4_cascade_\
        );

    \I__3833\ : InMux
    port map (
            O => \N__22336\,
            I => \N__22333\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__22333\,
            I => \this_ppu.un1_M_screen_x_q_c4\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__22330\,
            I => \N__22327\
        );

    \I__3830\ : InMux
    port map (
            O => \N__22327\,
            I => \N__22324\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__22324\,
            I => \N__22321\
        );

    \I__3828\ : Span4Mux_h
    port map (
            O => \N__22321\,
            I => \N__22317\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__22320\,
            I => \N__22314\
        );

    \I__3826\ : Span4Mux_h
    port map (
            O => \N__22317\,
            I => \N__22309\
        );

    \I__3825\ : InMux
    port map (
            O => \N__22314\,
            I => \N__22302\
        );

    \I__3824\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22302\
        );

    \I__3823\ : InMux
    port map (
            O => \N__22312\,
            I => \N__22302\
        );

    \I__3822\ : Odrv4
    port map (
            O => \N__22309\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__22302\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__22297\,
            I => \this_ppu.un1_M_screen_x_q_c5_cascade_\
        );

    \I__3819\ : CascadeMux
    port map (
            O => \N__22294\,
            I => \N__22291\
        );

    \I__3818\ : InMux
    port map (
            O => \N__22291\,
            I => \N__22288\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__22288\,
            I => \N__22285\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__22285\,
            I => \N__22282\
        );

    \I__3815\ : Span4Mux_h
    port map (
            O => \N__22282\,
            I => \N__22277\
        );

    \I__3814\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22272\
        );

    \I__3813\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22272\
        );

    \I__3812\ : Odrv4
    port map (
            O => \N__22277\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__22272\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__3810\ : CascadeMux
    port map (
            O => \N__22267\,
            I => \N__22264\
        );

    \I__3809\ : InMux
    port map (
            O => \N__22264\,
            I => \N__22261\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__22261\,
            I => \N__22258\
        );

    \I__3807\ : Span4Mux_v
    port map (
            O => \N__22258\,
            I => \N__22255\
        );

    \I__3806\ : Span4Mux_h
    port map (
            O => \N__22255\,
            I => \N__22251\
        );

    \I__3805\ : InMux
    port map (
            O => \N__22254\,
            I => \N__22248\
        );

    \I__3804\ : Odrv4
    port map (
            O => \N__22251\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__22248\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__3802\ : CascadeMux
    port map (
            O => \N__22243\,
            I => \N__22240\
        );

    \I__3801\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22237\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__22237\,
            I => \N__22234\
        );

    \I__3799\ : Span4Mux_v
    port map (
            O => \N__22234\,
            I => \N__22230\
        );

    \I__3798\ : CascadeMux
    port map (
            O => \N__22233\,
            I => \N__22226\
        );

    \I__3797\ : Span4Mux_h
    port map (
            O => \N__22230\,
            I => \N__22221\
        );

    \I__3796\ : InMux
    port map (
            O => \N__22229\,
            I => \N__22212\
        );

    \I__3795\ : InMux
    port map (
            O => \N__22226\,
            I => \N__22212\
        );

    \I__3794\ : InMux
    port map (
            O => \N__22225\,
            I => \N__22212\
        );

    \I__3793\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22212\
        );

    \I__3792\ : Odrv4
    port map (
            O => \N__22221\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__22212\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__3790\ : CascadeMux
    port map (
            O => \N__22207\,
            I => \N__22204\
        );

    \I__3789\ : InMux
    port map (
            O => \N__22204\,
            I => \N__22201\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__22201\,
            I => \M_this_scroll_qZ0Z_0\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__22198\,
            I => \N__22195\
        );

    \I__3786\ : InMux
    port map (
            O => \N__22195\,
            I => \N__22192\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__22192\,
            I => \N__22189\
        );

    \I__3784\ : Odrv4
    port map (
            O => \N__22189\,
            I => \M_this_scroll_qZ0Z_1\
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__22186\,
            I => \N__22182\
        );

    \I__3782\ : InMux
    port map (
            O => \N__22185\,
            I => \N__22175\
        );

    \I__3781\ : InMux
    port map (
            O => \N__22182\,
            I => \N__22175\
        );

    \I__3780\ : InMux
    port map (
            O => \N__22181\,
            I => \N__22172\
        );

    \I__3779\ : InMux
    port map (
            O => \N__22180\,
            I => \N__22169\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__22175\,
            I => \N__22166\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__22172\,
            I => \N__22161\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__22169\,
            I => \N__22157\
        );

    \I__3775\ : Span4Mux_v
    port map (
            O => \N__22166\,
            I => \N__22154\
        );

    \I__3774\ : InMux
    port map (
            O => \N__22165\,
            I => \N__22149\
        );

    \I__3773\ : InMux
    port map (
            O => \N__22164\,
            I => \N__22149\
        );

    \I__3772\ : Span4Mux_h
    port map (
            O => \N__22161\,
            I => \N__22146\
        );

    \I__3771\ : InMux
    port map (
            O => \N__22160\,
            I => \N__22143\
        );

    \I__3770\ : Span4Mux_h
    port map (
            O => \N__22157\,
            I => \N__22136\
        );

    \I__3769\ : Span4Mux_h
    port map (
            O => \N__22154\,
            I => \N__22136\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__22149\,
            I => \N__22136\
        );

    \I__3767\ : Odrv4
    port map (
            O => \N__22146\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__22143\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__22136\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__3764\ : InMux
    port map (
            O => \N__22129\,
            I => \N__22126\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__22126\,
            I => \N__22123\
        );

    \I__3762\ : Span4Mux_h
    port map (
            O => \N__22123\,
            I => \N__22120\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__22120\,
            I => \this_ppu.M_state_q_srsts_1_8\
        );

    \I__3760\ : InMux
    port map (
            O => \N__22117\,
            I => \N__22113\
        );

    \I__3759\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22110\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__22113\,
            I => \N__22107\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__22110\,
            I => \this_ppu.N_1145\
        );

    \I__3756\ : Odrv12
    port map (
            O => \N__22107\,
            I => \this_ppu.N_1145\
        );

    \I__3755\ : CascadeMux
    port map (
            O => \N__22102\,
            I => \N__22099\
        );

    \I__3754\ : InMux
    port map (
            O => \N__22099\,
            I => \N__22095\
        );

    \I__3753\ : CascadeMux
    port map (
            O => \N__22098\,
            I => \N__22092\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__22095\,
            I => \N__22089\
        );

    \I__3751\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22086\
        );

    \I__3750\ : Odrv4
    port map (
            O => \N__22089\,
            I => \this_ppu.M_screen_y_qZ0Z_7\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__22086\,
            I => \this_ppu.M_screen_y_qZ0Z_7\
        );

    \I__3748\ : InMux
    port map (
            O => \N__22081\,
            I => \N__22073\
        );

    \I__3747\ : InMux
    port map (
            O => \N__22080\,
            I => \N__22073\
        );

    \I__3746\ : InMux
    port map (
            O => \N__22079\,
            I => \N__22070\
        );

    \I__3745\ : InMux
    port map (
            O => \N__22078\,
            I => \N__22067\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__22073\,
            I => \N__22060\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__22070\,
            I => \N__22060\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__22067\,
            I => \N__22060\
        );

    \I__3741\ : Span4Mux_v
    port map (
            O => \N__22060\,
            I => \N__22057\
        );

    \I__3740\ : Odrv4
    port map (
            O => \N__22057\,
            I => \this_ppu.M_screen_y_qZ0Z_1\
        );

    \I__3739\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22051\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__22051\,
            I => \N__22048\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__22048\,
            I => \this_ppu.un3_M_screen_y_d_0_c2\
        );

    \I__3736\ : CascadeMux
    port map (
            O => \N__22045\,
            I => \this_ppu.un3_M_screen_y_d_0_c2_cascade_\
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__22042\,
            I => \this_ppu.un3_M_screen_y_d_0_c4_cascade_\
        );

    \I__3734\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22036\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__22036\,
            I => \this_ppu.un3_M_screen_y_d_0_c6\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__22033\,
            I => \N_861_0_cascade_\
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__22030\,
            I => \N__22026\
        );

    \I__3730\ : InMux
    port map (
            O => \N__22029\,
            I => \N__22022\
        );

    \I__3729\ : InMux
    port map (
            O => \N__22026\,
            I => \N__22017\
        );

    \I__3728\ : InMux
    port map (
            O => \N__22025\,
            I => \N__22017\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__22022\,
            I => \N__22014\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__22017\,
            I => \this_ppu.M_screen_y_qZ0Z_2\
        );

    \I__3725\ : Odrv4
    port map (
            O => \N__22014\,
            I => \this_ppu.M_screen_y_qZ0Z_2\
        );

    \I__3724\ : CascadeMux
    port map (
            O => \N__22009\,
            I => \N__22006\
        );

    \I__3723\ : InMux
    port map (
            O => \N__22006\,
            I => \N__22003\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__22003\,
            I => \N__21999\
        );

    \I__3721\ : InMux
    port map (
            O => \N__22002\,
            I => \N__21996\
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__21999\,
            I => \this_ppu.un3_M_screen_y_d_a_2\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__21996\,
            I => \this_ppu.un3_M_screen_y_d_a_2\
        );

    \I__3718\ : CascadeMux
    port map (
            O => \N__21991\,
            I => \N__21988\
        );

    \I__3717\ : InMux
    port map (
            O => \N__21988\,
            I => \N__21984\
        );

    \I__3716\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21981\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__21984\,
            I => \N__21978\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__21981\,
            I => \N__21975\
        );

    \I__3713\ : Span4Mux_v
    port map (
            O => \N__21978\,
            I => \N__21970\
        );

    \I__3712\ : Span4Mux_h
    port map (
            O => \N__21975\,
            I => \N__21970\
        );

    \I__3711\ : Odrv4
    port map (
            O => \N__21970\,
            I => \this_ppu.N_762_0\
        );

    \I__3710\ : InMux
    port map (
            O => \N__21967\,
            I => \N__21964\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__21964\,
            I => \N__21960\
        );

    \I__3708\ : InMux
    port map (
            O => \N__21963\,
            I => \N__21957\
        );

    \I__3707\ : Odrv12
    port map (
            O => \N__21960\,
            I => \this_ppu.N_91_0\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__21957\,
            I => \this_ppu.N_91_0\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__21952\,
            I => \this_ppu.N_91_0_cascade_\
        );

    \I__3704\ : InMux
    port map (
            O => \N__21949\,
            I => \N__21946\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__21946\,
            I => \this_ppu.un1_M_surface_x_q_c3\
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__21943\,
            I => \this_ppu.un1_M_surface_x_q_c3_cascade_\
        );

    \I__3701\ : InMux
    port map (
            O => \N__21940\,
            I => \N__21937\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__21937\,
            I => \this_ppu.un1_M_surface_x_q_c6\
        );

    \I__3699\ : CascadeMux
    port map (
            O => \N__21934\,
            I => \N__21931\
        );

    \I__3698\ : InMux
    port map (
            O => \N__21931\,
            I => \N__21928\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__21928\,
            I => \N__21925\
        );

    \I__3696\ : Odrv4
    port map (
            O => \N__21925\,
            I => \this_ppu.N_1202\
        );

    \I__3695\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21919\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__21919\,
            I => \N__21913\
        );

    \I__3693\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21910\
        );

    \I__3692\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21905\
        );

    \I__3691\ : InMux
    port map (
            O => \N__21916\,
            I => \N__21905\
        );

    \I__3690\ : Span4Mux_v
    port map (
            O => \N__21913\,
            I => \N__21900\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__21910\,
            I => \N__21900\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__21905\,
            I => \N__21897\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__21900\,
            I => \N__21894\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__21897\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__3685\ : Odrv4
    port map (
            O => \N__21894\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__3684\ : CascadeMux
    port map (
            O => \N__21889\,
            I => \N__21886\
        );

    \I__3683\ : InMux
    port map (
            O => \N__21886\,
            I => \N__21882\
        );

    \I__3682\ : CascadeMux
    port map (
            O => \N__21885\,
            I => \N__21879\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__21882\,
            I => \N__21875\
        );

    \I__3680\ : InMux
    port map (
            O => \N__21879\,
            I => \N__21872\
        );

    \I__3679\ : InMux
    port map (
            O => \N__21878\,
            I => \N__21869\
        );

    \I__3678\ : Span4Mux_v
    port map (
            O => \N__21875\,
            I => \N__21866\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__21872\,
            I => \N__21863\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__21869\,
            I => \N__21860\
        );

    \I__3675\ : Span4Mux_v
    port map (
            O => \N__21866\,
            I => \N__21857\
        );

    \I__3674\ : Span4Mux_h
    port map (
            O => \N__21863\,
            I => \N__21853\
        );

    \I__3673\ : Span12Mux_s7_v
    port map (
            O => \N__21860\,
            I => \N__21850\
        );

    \I__3672\ : Span4Mux_h
    port map (
            O => \N__21857\,
            I => \N__21847\
        );

    \I__3671\ : InMux
    port map (
            O => \N__21856\,
            I => \N__21844\
        );

    \I__3670\ : Span4Mux_v
    port map (
            O => \N__21853\,
            I => \N__21841\
        );

    \I__3669\ : Odrv12
    port map (
            O => \N__21850\,
            I => \M_this_status_flags_qZ0Z_0\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__21847\,
            I => \M_this_status_flags_qZ0Z_0\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__21844\,
            I => \M_this_status_flags_qZ0Z_0\
        );

    \I__3666\ : Odrv4
    port map (
            O => \N__21841\,
            I => \M_this_status_flags_qZ0Z_0\
        );

    \I__3665\ : InMux
    port map (
            O => \N__21832\,
            I => \N__21829\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__21829\,
            I => \this_ppu.N_1201\
        );

    \I__3663\ : InMux
    port map (
            O => \N__21826\,
            I => \M_this_data_count_q_cry_9\
        );

    \I__3662\ : InMux
    port map (
            O => \N__21823\,
            I => \M_this_data_count_q_cry_10\
        );

    \I__3661\ : InMux
    port map (
            O => \N__21820\,
            I => \M_this_data_count_q_cry_11\
        );

    \I__3660\ : InMux
    port map (
            O => \N__21817\,
            I => \M_this_data_count_q_cry_12\
        );

    \I__3659\ : CascadeMux
    port map (
            O => \N__21814\,
            I => \N__21811\
        );

    \I__3658\ : CascadeBuf
    port map (
            O => \N__21811\,
            I => \N__21808\
        );

    \I__3657\ : CascadeMux
    port map (
            O => \N__21808\,
            I => \N__21804\
        );

    \I__3656\ : CascadeMux
    port map (
            O => \N__21807\,
            I => \N__21801\
        );

    \I__3655\ : InMux
    port map (
            O => \N__21804\,
            I => \N__21798\
        );

    \I__3654\ : InMux
    port map (
            O => \N__21801\,
            I => \N__21795\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__21798\,
            I => \N__21792\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__21795\,
            I => \M_this_oam_address_qZ0Z_7\
        );

    \I__3651\ : Odrv12
    port map (
            O => \N__21792\,
            I => \M_this_oam_address_qZ0Z_7\
        );

    \I__3650\ : IoInMux
    port map (
            O => \N__21787\,
            I => \N__21784\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__21784\,
            I => \N__21781\
        );

    \I__3648\ : Odrv12
    port map (
            O => \N__21781\,
            I => \IO_port_data_write_i_m2_i_m2_0\
        );

    \I__3647\ : IoInMux
    port map (
            O => \N__21778\,
            I => \N__21775\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__21775\,
            I => \N__21772\
        );

    \I__3645\ : IoSpan4Mux
    port map (
            O => \N__21772\,
            I => \N__21769\
        );

    \I__3644\ : Sp12to4
    port map (
            O => \N__21769\,
            I => \N__21766\
        );

    \I__3643\ : Span12Mux_v
    port map (
            O => \N__21766\,
            I => \N__21763\
        );

    \I__3642\ : Odrv12
    port map (
            O => \N__21763\,
            I => \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\
        );

    \I__3641\ : InMux
    port map (
            O => \N__21760\,
            I => \N__21757\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__21757\,
            I => \this_ppu.M_state_qZ0Z_8\
        );

    \I__3639\ : InMux
    port map (
            O => \N__21754\,
            I => \M_this_data_count_q_cry_0\
        );

    \I__3638\ : InMux
    port map (
            O => \N__21751\,
            I => \M_this_data_count_q_cry_1\
        );

    \I__3637\ : InMux
    port map (
            O => \N__21748\,
            I => \M_this_data_count_q_cry_2\
        );

    \I__3636\ : InMux
    port map (
            O => \N__21745\,
            I => \M_this_data_count_q_cry_3\
        );

    \I__3635\ : InMux
    port map (
            O => \N__21742\,
            I => \M_this_data_count_q_cry_4\
        );

    \I__3634\ : InMux
    port map (
            O => \N__21739\,
            I => \M_this_data_count_q_cry_5\
        );

    \I__3633\ : InMux
    port map (
            O => \N__21736\,
            I => \M_this_data_count_q_cry_6\
        );

    \I__3632\ : InMux
    port map (
            O => \N__21733\,
            I => \bfn_14_25_0_\
        );

    \I__3631\ : InMux
    port map (
            O => \N__21730\,
            I => \M_this_data_count_q_cry_8\
        );

    \I__3630\ : InMux
    port map (
            O => \N__21727\,
            I => \bfn_14_22_0_\
        );

    \I__3629\ : CascadeMux
    port map (
            O => \N__21724\,
            I => \N__21721\
        );

    \I__3628\ : CascadeBuf
    port map (
            O => \N__21721\,
            I => \N__21718\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__21718\,
            I => \N__21715\
        );

    \I__3626\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21712\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__21712\,
            I => \N__21709\
        );

    \I__3624\ : Span4Mux_s2_v
    port map (
            O => \N__21709\,
            I => \N__21706\
        );

    \I__3623\ : Sp12to4
    port map (
            O => \N__21706\,
            I => \N__21702\
        );

    \I__3622\ : InMux
    port map (
            O => \N__21705\,
            I => \N__21699\
        );

    \I__3621\ : Span12Mux_s6_h
    port map (
            O => \N__21702\,
            I => \N__21696\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__21699\,
            I => \N__21693\
        );

    \I__3619\ : Span12Mux_h
    port map (
            O => \N__21696\,
            I => \N__21690\
        );

    \I__3618\ : Odrv12
    port map (
            O => \N__21693\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__3617\ : Odrv12
    port map (
            O => \N__21690\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__3616\ : InMux
    port map (
            O => \N__21685\,
            I => \N__21682\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__21682\,
            I => \N__21679\
        );

    \I__3614\ : Odrv4
    port map (
            O => \N__21679\,
            I => \this_ppu.M_screen_y_q_esr_RNI563Q6Z0Z_2\
        );

    \I__3613\ : InMux
    port map (
            O => \N__21676\,
            I => \N__21673\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__21673\,
            I => \N__21669\
        );

    \I__3611\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21666\
        );

    \I__3610\ : Span4Mux_h
    port map (
            O => \N__21669\,
            I => \N__21661\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__21666\,
            I => \N__21661\
        );

    \I__3608\ : Span4Mux_h
    port map (
            O => \N__21661\,
            I => \N__21658\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__21658\,
            I => \M_this_oam_ram_read_data_23\
        );

    \I__3606\ : InMux
    port map (
            O => \N__21655\,
            I => \N__21652\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__21652\,
            I => \N__21649\
        );

    \I__3604\ : Span4Mux_h
    port map (
            O => \N__21649\,
            I => \N__21646\
        );

    \I__3603\ : Span4Mux_h
    port map (
            O => \N__21646\,
            I => \N__21643\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__21643\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_23\
        );

    \I__3601\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21637\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__21637\,
            I => \N__21633\
        );

    \I__3599\ : InMux
    port map (
            O => \N__21636\,
            I => \N__21630\
        );

    \I__3598\ : Span4Mux_h
    port map (
            O => \N__21633\,
            I => \N__21627\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__21630\,
            I => \N__21624\
        );

    \I__3596\ : Span4Mux_h
    port map (
            O => \N__21627\,
            I => \N__21621\
        );

    \I__3595\ : Span4Mux_h
    port map (
            O => \N__21624\,
            I => \N__21618\
        );

    \I__3594\ : Odrv4
    port map (
            O => \N__21621\,
            I => \M_this_oam_ram_read_data_1\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__21618\,
            I => \M_this_oam_ram_read_data_1\
        );

    \I__3592\ : InMux
    port map (
            O => \N__21613\,
            I => \N__21610\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__21610\,
            I => \N__21607\
        );

    \I__3590\ : Span4Mux_h
    port map (
            O => \N__21607\,
            I => \N__21604\
        );

    \I__3589\ : Span4Mux_v
    port map (
            O => \N__21604\,
            I => \N__21601\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__21601\,
            I => \this_ppu.oam_cache.N_581_0\
        );

    \I__3587\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21595\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__21595\,
            I => \M_this_data_tmp_qZ0Z_13\
        );

    \I__3585\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21589\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__21589\,
            I => \this_ppu.m13_0_i_1\
        );

    \I__3583\ : InMux
    port map (
            O => \N__21586\,
            I => \N__21582\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__21585\,
            I => \N__21579\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__21582\,
            I => \N__21576\
        );

    \I__3580\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21573\
        );

    \I__3579\ : Span4Mux_h
    port map (
            O => \N__21576\,
            I => \N__21569\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__21573\,
            I => \N__21566\
        );

    \I__3577\ : InMux
    port map (
            O => \N__21572\,
            I => \N__21563\
        );

    \I__3576\ : Span4Mux_h
    port map (
            O => \N__21569\,
            I => \N__21560\
        );

    \I__3575\ : Span4Mux_h
    port map (
            O => \N__21566\,
            I => \N__21557\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__21563\,
            I => \this_ppu.offset_y\
        );

    \I__3573\ : Odrv4
    port map (
            O => \N__21560\,
            I => \this_ppu.offset_y\
        );

    \I__3572\ : Odrv4
    port map (
            O => \N__21557\,
            I => \this_ppu.offset_y\
        );

    \I__3571\ : InMux
    port map (
            O => \N__21550\,
            I => \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO\
        );

    \I__3570\ : InMux
    port map (
            O => \N__21547\,
            I => \N__21544\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__21544\,
            I => \this_ppu.M_screen_y_q_esr_RNI453Q6Z0Z_1\
        );

    \I__3568\ : CascadeMux
    port map (
            O => \N__21541\,
            I => \N__21537\
        );

    \I__3567\ : CascadeMux
    port map (
            O => \N__21540\,
            I => \N__21534\
        );

    \I__3566\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21531\
        );

    \I__3565\ : InMux
    port map (
            O => \N__21534\,
            I => \N__21528\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__21531\,
            I => \N__21525\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__21528\,
            I => \N__21522\
        );

    \I__3562\ : Span12Mux_h
    port map (
            O => \N__21525\,
            I => \N__21519\
        );

    \I__3561\ : Span4Mux_h
    port map (
            O => \N__21522\,
            I => \N__21516\
        );

    \I__3560\ : Odrv12
    port map (
            O => \N__21519\,
            I => \this_ppu.M_surface_y_qZ0Z_1\
        );

    \I__3559\ : Odrv4
    port map (
            O => \N__21516\,
            I => \this_ppu.M_surface_y_qZ0Z_1\
        );

    \I__3558\ : InMux
    port map (
            O => \N__21511\,
            I => \this_ppu.un1_M_surface_y_d_cry_0\
        );

    \I__3557\ : CascadeMux
    port map (
            O => \N__21508\,
            I => \N__21505\
        );

    \I__3556\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21501\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__21504\,
            I => \N__21498\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__21501\,
            I => \N__21495\
        );

    \I__3553\ : InMux
    port map (
            O => \N__21498\,
            I => \N__21492\
        );

    \I__3552\ : Span4Mux_v
    port map (
            O => \N__21495\,
            I => \N__21489\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__21492\,
            I => \N__21486\
        );

    \I__3550\ : Span4Mux_h
    port map (
            O => \N__21489\,
            I => \N__21481\
        );

    \I__3549\ : Span4Mux_v
    port map (
            O => \N__21486\,
            I => \N__21481\
        );

    \I__3548\ : Odrv4
    port map (
            O => \N__21481\,
            I => \this_ppu.M_surface_y_qZ0Z_2\
        );

    \I__3547\ : InMux
    port map (
            O => \N__21478\,
            I => \this_ppu.un1_M_surface_y_d_cry_1\
        );

    \I__3546\ : CascadeMux
    port map (
            O => \N__21475\,
            I => \N__21472\
        );

    \I__3545\ : CascadeBuf
    port map (
            O => \N__21472\,
            I => \N__21469\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__21469\,
            I => \N__21465\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__21468\,
            I => \N__21462\
        );

    \I__3542\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21459\
        );

    \I__3541\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21456\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__21459\,
            I => \N__21453\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__21456\,
            I => \N__21450\
        );

    \I__3538\ : Sp12to4
    port map (
            O => \N__21453\,
            I => \N__21447\
        );

    \I__3537\ : Span4Mux_v
    port map (
            O => \N__21450\,
            I => \N__21444\
        );

    \I__3536\ : Span12Mux_s11_v
    port map (
            O => \N__21447\,
            I => \N__21441\
        );

    \I__3535\ : Odrv4
    port map (
            O => \N__21444\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__3534\ : Odrv12
    port map (
            O => \N__21441\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__3533\ : InMux
    port map (
            O => \N__21436\,
            I => \this_ppu.un1_M_surface_y_d_cry_2\
        );

    \I__3532\ : InMux
    port map (
            O => \N__21433\,
            I => \N__21430\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__21430\,
            I => \this_ppu.M_screen_y_q_RNI8FJF7Z0Z_4\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__21427\,
            I => \N__21424\
        );

    \I__3529\ : CascadeBuf
    port map (
            O => \N__21424\,
            I => \N__21420\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__21423\,
            I => \N__21417\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__21420\,
            I => \N__21414\
        );

    \I__3526\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21411\
        );

    \I__3525\ : InMux
    port map (
            O => \N__21414\,
            I => \N__21408\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__21411\,
            I => \N__21405\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__21408\,
            I => \N__21402\
        );

    \I__3522\ : Span4Mux_v
    port map (
            O => \N__21405\,
            I => \N__21399\
        );

    \I__3521\ : Span12Mux_s11_v
    port map (
            O => \N__21402\,
            I => \N__21396\
        );

    \I__3520\ : Odrv4
    port map (
            O => \N__21399\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__3519\ : Odrv12
    port map (
            O => \N__21396\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__3518\ : InMux
    port map (
            O => \N__21391\,
            I => \this_ppu.un1_M_surface_y_d_cry_3\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__21388\,
            I => \N__21385\
        );

    \I__3516\ : CascadeBuf
    port map (
            O => \N__21385\,
            I => \N__21382\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__21382\,
            I => \N__21379\
        );

    \I__3514\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21375\
        );

    \I__3513\ : InMux
    port map (
            O => \N__21378\,
            I => \N__21372\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__21375\,
            I => \N__21369\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__21372\,
            I => \N__21366\
        );

    \I__3510\ : Span4Mux_h
    port map (
            O => \N__21369\,
            I => \N__21363\
        );

    \I__3509\ : Span4Mux_h
    port map (
            O => \N__21366\,
            I => \N__21360\
        );

    \I__3508\ : Sp12to4
    port map (
            O => \N__21363\,
            I => \N__21357\
        );

    \I__3507\ : Span4Mux_h
    port map (
            O => \N__21360\,
            I => \N__21354\
        );

    \I__3506\ : Span12Mux_s11_v
    port map (
            O => \N__21357\,
            I => \N__21351\
        );

    \I__3505\ : Odrv4
    port map (
            O => \N__21354\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__3504\ : Odrv12
    port map (
            O => \N__21351\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__3503\ : InMux
    port map (
            O => \N__21346\,
            I => \this_ppu.un1_M_surface_y_d_cry_4\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__21343\,
            I => \N__21340\
        );

    \I__3501\ : CascadeBuf
    port map (
            O => \N__21340\,
            I => \N__21337\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__21337\,
            I => \N__21334\
        );

    \I__3499\ : InMux
    port map (
            O => \N__21334\,
            I => \N__21331\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__21331\,
            I => \N__21327\
        );

    \I__3497\ : InMux
    port map (
            O => \N__21330\,
            I => \N__21324\
        );

    \I__3496\ : Sp12to4
    port map (
            O => \N__21327\,
            I => \N__21321\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__21324\,
            I => \N__21318\
        );

    \I__3494\ : Span12Mux_s4_v
    port map (
            O => \N__21321\,
            I => \N__21315\
        );

    \I__3493\ : Span4Mux_h
    port map (
            O => \N__21318\,
            I => \N__21312\
        );

    \I__3492\ : Span12Mux_h
    port map (
            O => \N__21315\,
            I => \N__21309\
        );

    \I__3491\ : Odrv4
    port map (
            O => \N__21312\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__3490\ : Odrv12
    port map (
            O => \N__21309\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__3489\ : InMux
    port map (
            O => \N__21304\,
            I => \this_ppu.un1_M_surface_y_d_cry_5\
        );

    \I__3488\ : InMux
    port map (
            O => \N__21301\,
            I => \N__21298\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__21298\,
            I => \N__21295\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__21295\,
            I => \this_ppu.M_oam_cache_read_data_i_12\
        );

    \I__3485\ : InMux
    port map (
            O => \N__21292\,
            I => \N__21289\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__21289\,
            I => \this_ppu.offset_x_4\
        );

    \I__3483\ : InMux
    port map (
            O => \N__21286\,
            I => \this_ppu.offset_x_cry_3\
        );

    \I__3482\ : InMux
    port map (
            O => \N__21283\,
            I => \N__21280\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__21280\,
            I => \this_ppu.M_oam_cache_read_data_i_13\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__21277\,
            I => \N__21274\
        );

    \I__3479\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21271\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__21271\,
            I => \this_ppu.offset_x_5\
        );

    \I__3477\ : InMux
    port map (
            O => \N__21268\,
            I => \this_ppu.offset_x_cry_4\
        );

    \I__3476\ : InMux
    port map (
            O => \N__21265\,
            I => \N__21262\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__21262\,
            I => \this_ppu.M_oam_cache_read_data_i_14\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__21259\,
            I => \N__21256\
        );

    \I__3473\ : CascadeBuf
    port map (
            O => \N__21256\,
            I => \N__21253\
        );

    \I__3472\ : CascadeMux
    port map (
            O => \N__21253\,
            I => \N__21250\
        );

    \I__3471\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21247\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__21247\,
            I => \N__21244\
        );

    \I__3469\ : Span4Mux_s2_v
    port map (
            O => \N__21244\,
            I => \N__21239\
        );

    \I__3468\ : InMux
    port map (
            O => \N__21243\,
            I => \N__21235\
        );

    \I__3467\ : CascadeMux
    port map (
            O => \N__21242\,
            I => \N__21232\
        );

    \I__3466\ : Sp12to4
    port map (
            O => \N__21239\,
            I => \N__21229\
        );

    \I__3465\ : InMux
    port map (
            O => \N__21238\,
            I => \N__21226\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__21235\,
            I => \N__21223\
        );

    \I__3463\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21220\
        );

    \I__3462\ : Span12Mux_v
    port map (
            O => \N__21229\,
            I => \N__21217\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__21226\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__3460\ : Odrv12
    port map (
            O => \N__21223\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__21220\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__3458\ : Odrv12
    port map (
            O => \N__21217\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__3457\ : InMux
    port map (
            O => \N__21208\,
            I => \N__21205\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__21205\,
            I => \this_ppu.offset_x_6\
        );

    \I__3455\ : InMux
    port map (
            O => \N__21202\,
            I => \this_ppu.offset_x_cry_5\
        );

    \I__3454\ : InMux
    port map (
            O => \N__21199\,
            I => \N__21196\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__21196\,
            I => \N__21193\
        );

    \I__3452\ : Span4Mux_v
    port map (
            O => \N__21193\,
            I => \N__21190\
        );

    \I__3451\ : Odrv4
    port map (
            O => \N__21190\,
            I => \this_ppu.M_oam_cache_read_data_15\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__21187\,
            I => \N__21184\
        );

    \I__3449\ : CascadeBuf
    port map (
            O => \N__21184\,
            I => \N__21181\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__21181\,
            I => \N__21178\
        );

    \I__3447\ : InMux
    port map (
            O => \N__21178\,
            I => \N__21175\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__21175\,
            I => \N__21172\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__21172\,
            I => \N__21168\
        );

    \I__3444\ : InMux
    port map (
            O => \N__21171\,
            I => \N__21164\
        );

    \I__3443\ : Sp12to4
    port map (
            O => \N__21168\,
            I => \N__21161\
        );

    \I__3442\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21158\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__21164\,
            I => \N__21153\
        );

    \I__3440\ : Span12Mux_h
    port map (
            O => \N__21161\,
            I => \N__21153\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__21158\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__3438\ : Odrv12
    port map (
            O => \N__21153\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__3437\ : InMux
    port map (
            O => \N__21148\,
            I => \bfn_14_20_0_\
        );

    \I__3436\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21142\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__21142\,
            I => \this_ppu.offset_x_7\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__21139\,
            I => \N__21136\
        );

    \I__3433\ : InMux
    port map (
            O => \N__21136\,
            I => \N__21129\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__21135\,
            I => \N__21123\
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__21134\,
            I => \N__21120\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__21133\,
            I => \N__21117\
        );

    \I__3429\ : CascadeMux
    port map (
            O => \N__21132\,
            I => \N__21113\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__21129\,
            I => \N__21108\
        );

    \I__3427\ : CascadeMux
    port map (
            O => \N__21128\,
            I => \N__21105\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__21127\,
            I => \N__21100\
        );

    \I__3425\ : CascadeMux
    port map (
            O => \N__21126\,
            I => \N__21097\
        );

    \I__3424\ : InMux
    port map (
            O => \N__21123\,
            I => \N__21094\
        );

    \I__3423\ : InMux
    port map (
            O => \N__21120\,
            I => \N__21091\
        );

    \I__3422\ : InMux
    port map (
            O => \N__21117\,
            I => \N__21088\
        );

    \I__3421\ : CascadeMux
    port map (
            O => \N__21116\,
            I => \N__21085\
        );

    \I__3420\ : InMux
    port map (
            O => \N__21113\,
            I => \N__21079\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__21112\,
            I => \N__21076\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__21111\,
            I => \N__21073\
        );

    \I__3417\ : Span4Mux_h
    port map (
            O => \N__21108\,
            I => \N__21070\
        );

    \I__3416\ : InMux
    port map (
            O => \N__21105\,
            I => \N__21067\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__21104\,
            I => \N__21064\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__21103\,
            I => \N__21061\
        );

    \I__3413\ : InMux
    port map (
            O => \N__21100\,
            I => \N__21058\
        );

    \I__3412\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21055\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__21094\,
            I => \N__21052\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__21091\,
            I => \N__21047\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__21088\,
            I => \N__21047\
        );

    \I__3408\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21044\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__21084\,
            I => \N__21041\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__21083\,
            I => \N__21038\
        );

    \I__3405\ : CascadeMux
    port map (
            O => \N__21082\,
            I => \N__21035\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__21079\,
            I => \N__21032\
        );

    \I__3403\ : InMux
    port map (
            O => \N__21076\,
            I => \N__21029\
        );

    \I__3402\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21026\
        );

    \I__3401\ : IoSpan4Mux
    port map (
            O => \N__21070\,
            I => \N__21023\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__21067\,
            I => \N__21020\
        );

    \I__3399\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21017\
        );

    \I__3398\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21014\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__21058\,
            I => \N__21011\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__21055\,
            I => \N__21002\
        );

    \I__3395\ : Span4Mux_v
    port map (
            O => \N__21052\,
            I => \N__21002\
        );

    \I__3394\ : Span4Mux_v
    port map (
            O => \N__21047\,
            I => \N__21002\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__21044\,
            I => \N__21002\
        );

    \I__3392\ : InMux
    port map (
            O => \N__21041\,
            I => \N__20999\
        );

    \I__3391\ : InMux
    port map (
            O => \N__21038\,
            I => \N__20996\
        );

    \I__3390\ : InMux
    port map (
            O => \N__21035\,
            I => \N__20993\
        );

    \I__3389\ : Span4Mux_v
    port map (
            O => \N__21032\,
            I => \N__20990\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__21029\,
            I => \N__20985\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__21026\,
            I => \N__20985\
        );

    \I__3386\ : IoSpan4Mux
    port map (
            O => \N__21023\,
            I => \N__20982\
        );

    \I__3385\ : Span4Mux_h
    port map (
            O => \N__21020\,
            I => \N__20979\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__21017\,
            I => \N__20974\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__21014\,
            I => \N__20974\
        );

    \I__3382\ : Span4Mux_v
    port map (
            O => \N__21011\,
            I => \N__20971\
        );

    \I__3381\ : Span4Mux_v
    port map (
            O => \N__21002\,
            I => \N__20966\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20966\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__20996\,
            I => \N__20961\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__20993\,
            I => \N__20961\
        );

    \I__3377\ : Span4Mux_h
    port map (
            O => \N__20990\,
            I => \N__20956\
        );

    \I__3376\ : Span4Mux_v
    port map (
            O => \N__20985\,
            I => \N__20956\
        );

    \I__3375\ : Span4Mux_s3_v
    port map (
            O => \N__20982\,
            I => \N__20951\
        );

    \I__3374\ : Span4Mux_h
    port map (
            O => \N__20979\,
            I => \N__20951\
        );

    \I__3373\ : Span4Mux_v
    port map (
            O => \N__20974\,
            I => \N__20948\
        );

    \I__3372\ : Span4Mux_h
    port map (
            O => \N__20971\,
            I => \N__20945\
        );

    \I__3371\ : Span4Mux_v
    port map (
            O => \N__20966\,
            I => \N__20940\
        );

    \I__3370\ : Span4Mux_v
    port map (
            O => \N__20961\,
            I => \N__20940\
        );

    \I__3369\ : Sp12to4
    port map (
            O => \N__20956\,
            I => \N__20937\
        );

    \I__3368\ : Span4Mux_v
    port map (
            O => \N__20951\,
            I => \N__20934\
        );

    \I__3367\ : Sp12to4
    port map (
            O => \N__20948\,
            I => \N__20931\
        );

    \I__3366\ : Sp12to4
    port map (
            O => \N__20945\,
            I => \N__20926\
        );

    \I__3365\ : Sp12to4
    port map (
            O => \N__20940\,
            I => \N__20926\
        );

    \I__3364\ : Span12Mux_h
    port map (
            O => \N__20937\,
            I => \N__20923\
        );

    \I__3363\ : Span4Mux_v
    port map (
            O => \N__20934\,
            I => \N__20920\
        );

    \I__3362\ : Span12Mux_h
    port map (
            O => \N__20931\,
            I => \N__20915\
        );

    \I__3361\ : Span12Mux_h
    port map (
            O => \N__20926\,
            I => \N__20915\
        );

    \I__3360\ : Span12Mux_v
    port map (
            O => \N__20923\,
            I => \N__20912\
        );

    \I__3359\ : Odrv4
    port map (
            O => \N__20920\,
            I => \M_this_ppu_spr_addr_0\
        );

    \I__3358\ : Odrv12
    port map (
            O => \N__20915\,
            I => \M_this_ppu_spr_addr_0\
        );

    \I__3357\ : Odrv12
    port map (
            O => \N__20912\,
            I => \M_this_ppu_spr_addr_0\
        );

    \I__3356\ : CascadeMux
    port map (
            O => \N__20905\,
            I => \N__20902\
        );

    \I__3355\ : InMux
    port map (
            O => \N__20902\,
            I => \N__20898\
        );

    \I__3354\ : InMux
    port map (
            O => \N__20901\,
            I => \N__20895\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__20898\,
            I => \this_ppu.M_oam_cache_read_data_8\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__20895\,
            I => \this_ppu.M_oam_cache_read_data_8\
        );

    \I__3351\ : InMux
    port map (
            O => \N__20890\,
            I => \N__20887\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__20887\,
            I => \this_ppu.M_oam_cache_read_data_i_8\
        );

    \I__3349\ : InMux
    port map (
            O => \N__20884\,
            I => \N__20881\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__20881\,
            I => \this_ppu.M_oam_cache_read_data_i_9\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__20878\,
            I => \N__20875\
        );

    \I__3346\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20871\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__20874\,
            I => \N__20868\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__20871\,
            I => \N__20864\
        );

    \I__3343\ : InMux
    port map (
            O => \N__20868\,
            I => \N__20861\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__20867\,
            I => \N__20858\
        );

    \I__3341\ : Span4Mux_s2_v
    port map (
            O => \N__20864\,
            I => \N__20852\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__20861\,
            I => \N__20852\
        );

    \I__3339\ : InMux
    port map (
            O => \N__20858\,
            I => \N__20849\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__20857\,
            I => \N__20846\
        );

    \I__3337\ : Span4Mux_v
    port map (
            O => \N__20852\,
            I => \N__20840\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__20849\,
            I => \N__20840\
        );

    \I__3335\ : InMux
    port map (
            O => \N__20846\,
            I => \N__20837\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__20845\,
            I => \N__20834\
        );

    \I__3333\ : Span4Mux_h
    port map (
            O => \N__20840\,
            I => \N__20824\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__20837\,
            I => \N__20824\
        );

    \I__3331\ : InMux
    port map (
            O => \N__20834\,
            I => \N__20821\
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__20833\,
            I => \N__20818\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__20832\,
            I => \N__20814\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__20831\,
            I => \N__20811\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__20830\,
            I => \N__20807\
        );

    \I__3326\ : CascadeMux
    port map (
            O => \N__20829\,
            I => \N__20804\
        );

    \I__3325\ : Span4Mux_v
    port map (
            O => \N__20824\,
            I => \N__20797\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__20821\,
            I => \N__20797\
        );

    \I__3323\ : InMux
    port map (
            O => \N__20818\,
            I => \N__20794\
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__20817\,
            I => \N__20791\
        );

    \I__3321\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20787\
        );

    \I__3320\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20784\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__20810\,
            I => \N__20781\
        );

    \I__3318\ : InMux
    port map (
            O => \N__20807\,
            I => \N__20778\
        );

    \I__3317\ : InMux
    port map (
            O => \N__20804\,
            I => \N__20775\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__20803\,
            I => \N__20772\
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__20802\,
            I => \N__20769\
        );

    \I__3314\ : Span4Mux_h
    port map (
            O => \N__20797\,
            I => \N__20764\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__20794\,
            I => \N__20764\
        );

    \I__3312\ : InMux
    port map (
            O => \N__20791\,
            I => \N__20761\
        );

    \I__3311\ : CascadeMux
    port map (
            O => \N__20790\,
            I => \N__20758\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__20787\,
            I => \N__20752\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__20784\,
            I => \N__20752\
        );

    \I__3308\ : InMux
    port map (
            O => \N__20781\,
            I => \N__20749\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__20778\,
            I => \N__20744\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__20775\,
            I => \N__20744\
        );

    \I__3305\ : InMux
    port map (
            O => \N__20772\,
            I => \N__20741\
        );

    \I__3304\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20738\
        );

    \I__3303\ : Span4Mux_v
    port map (
            O => \N__20764\,
            I => \N__20733\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__20761\,
            I => \N__20733\
        );

    \I__3301\ : InMux
    port map (
            O => \N__20758\,
            I => \N__20730\
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__20757\,
            I => \N__20727\
        );

    \I__3299\ : Span4Mux_v
    port map (
            O => \N__20752\,
            I => \N__20722\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__20749\,
            I => \N__20722\
        );

    \I__3297\ : Span4Mux_v
    port map (
            O => \N__20744\,
            I => \N__20715\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__20741\,
            I => \N__20715\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__20738\,
            I => \N__20715\
        );

    \I__3294\ : Span4Mux_h
    port map (
            O => \N__20733\,
            I => \N__20710\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__20730\,
            I => \N__20710\
        );

    \I__3292\ : InMux
    port map (
            O => \N__20727\,
            I => \N__20707\
        );

    \I__3291\ : Span4Mux_v
    port map (
            O => \N__20722\,
            I => \N__20704\
        );

    \I__3290\ : Span4Mux_v
    port map (
            O => \N__20715\,
            I => \N__20697\
        );

    \I__3289\ : Span4Mux_v
    port map (
            O => \N__20710\,
            I => \N__20697\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__20707\,
            I => \N__20697\
        );

    \I__3287\ : Span4Mux_h
    port map (
            O => \N__20704\,
            I => \N__20694\
        );

    \I__3286\ : Span4Mux_h
    port map (
            O => \N__20697\,
            I => \N__20691\
        );

    \I__3285\ : Span4Mux_v
    port map (
            O => \N__20694\,
            I => \N__20688\
        );

    \I__3284\ : Span4Mux_h
    port map (
            O => \N__20691\,
            I => \N__20685\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__20688\,
            I => \M_this_ppu_spr_addr_1\
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__20685\,
            I => \M_this_ppu_spr_addr_1\
        );

    \I__3281\ : InMux
    port map (
            O => \N__20680\,
            I => \this_ppu.offset_x_cry_0\
        );

    \I__3280\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20674\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__20674\,
            I => \N__20671\
        );

    \I__3278\ : Span4Mux_h
    port map (
            O => \N__20671\,
            I => \N__20668\
        );

    \I__3277\ : Odrv4
    port map (
            O => \N__20668\,
            I => \this_ppu.M_oam_cache_read_data_i_10\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__20665\,
            I => \N__20662\
        );

    \I__3275\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20658\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__20661\,
            I => \N__20655\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__20658\,
            I => \N__20649\
        );

    \I__3272\ : InMux
    port map (
            O => \N__20655\,
            I => \N__20646\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__20654\,
            I => \N__20643\
        );

    \I__3270\ : CascadeMux
    port map (
            O => \N__20653\,
            I => \N__20636\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__20652\,
            I => \N__20633\
        );

    \I__3268\ : Span4Mux_h
    port map (
            O => \N__20649\,
            I => \N__20627\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__20646\,
            I => \N__20627\
        );

    \I__3266\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20624\
        );

    \I__3265\ : CascadeMux
    port map (
            O => \N__20642\,
            I => \N__20621\
        );

    \I__3264\ : CascadeMux
    port map (
            O => \N__20641\,
            I => \N__20617\
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__20640\,
            I => \N__20614\
        );

    \I__3262\ : CascadeMux
    port map (
            O => \N__20639\,
            I => \N__20611\
        );

    \I__3261\ : InMux
    port map (
            O => \N__20636\,
            I => \N__20606\
        );

    \I__3260\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20602\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__20632\,
            I => \N__20599\
        );

    \I__3258\ : Span4Mux_v
    port map (
            O => \N__20627\,
            I => \N__20594\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__20624\,
            I => \N__20594\
        );

    \I__3256\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20591\
        );

    \I__3255\ : CascadeMux
    port map (
            O => \N__20620\,
            I => \N__20588\
        );

    \I__3254\ : InMux
    port map (
            O => \N__20617\,
            I => \N__20585\
        );

    \I__3253\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20582\
        );

    \I__3252\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20579\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__20610\,
            I => \N__20576\
        );

    \I__3250\ : CascadeMux
    port map (
            O => \N__20609\,
            I => \N__20573\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__20606\,
            I => \N__20569\
        );

    \I__3248\ : CascadeMux
    port map (
            O => \N__20605\,
            I => \N__20566\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__20602\,
            I => \N__20562\
        );

    \I__3246\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20559\
        );

    \I__3245\ : Span4Mux_h
    port map (
            O => \N__20594\,
            I => \N__20554\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__20591\,
            I => \N__20554\
        );

    \I__3243\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20551\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__20585\,
            I => \N__20548\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__20582\,
            I => \N__20545\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__20579\,
            I => \N__20542\
        );

    \I__3239\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20539\
        );

    \I__3238\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20536\
        );

    \I__3237\ : CascadeMux
    port map (
            O => \N__20572\,
            I => \N__20533\
        );

    \I__3236\ : Span4Mux_v
    port map (
            O => \N__20569\,
            I => \N__20530\
        );

    \I__3235\ : InMux
    port map (
            O => \N__20566\,
            I => \N__20527\
        );

    \I__3234\ : CascadeMux
    port map (
            O => \N__20565\,
            I => \N__20524\
        );

    \I__3233\ : Span4Mux_h
    port map (
            O => \N__20562\,
            I => \N__20521\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__20559\,
            I => \N__20518\
        );

    \I__3231\ : Span4Mux_v
    port map (
            O => \N__20554\,
            I => \N__20513\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20513\
        );

    \I__3229\ : Span4Mux_v
    port map (
            O => \N__20548\,
            I => \N__20504\
        );

    \I__3228\ : Span4Mux_v
    port map (
            O => \N__20545\,
            I => \N__20504\
        );

    \I__3227\ : Span4Mux_h
    port map (
            O => \N__20542\,
            I => \N__20504\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__20539\,
            I => \N__20504\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__20536\,
            I => \N__20501\
        );

    \I__3224\ : InMux
    port map (
            O => \N__20533\,
            I => \N__20498\
        );

    \I__3223\ : Sp12to4
    port map (
            O => \N__20530\,
            I => \N__20493\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__20527\,
            I => \N__20493\
        );

    \I__3221\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20490\
        );

    \I__3220\ : Span4Mux_v
    port map (
            O => \N__20521\,
            I => \N__20485\
        );

    \I__3219\ : Span4Mux_h
    port map (
            O => \N__20518\,
            I => \N__20485\
        );

    \I__3218\ : Span4Mux_h
    port map (
            O => \N__20513\,
            I => \N__20482\
        );

    \I__3217\ : Span4Mux_v
    port map (
            O => \N__20504\,
            I => \N__20475\
        );

    \I__3216\ : Span4Mux_v
    port map (
            O => \N__20501\,
            I => \N__20475\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__20498\,
            I => \N__20475\
        );

    \I__3214\ : Span12Mux_h
    port map (
            O => \N__20493\,
            I => \N__20472\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__20490\,
            I => \N__20469\
        );

    \I__3212\ : Span4Mux_h
    port map (
            O => \N__20485\,
            I => \N__20466\
        );

    \I__3211\ : Span4Mux_v
    port map (
            O => \N__20482\,
            I => \N__20461\
        );

    \I__3210\ : Span4Mux_h
    port map (
            O => \N__20475\,
            I => \N__20461\
        );

    \I__3209\ : Span12Mux_v
    port map (
            O => \N__20472\,
            I => \N__20454\
        );

    \I__3208\ : Span12Mux_h
    port map (
            O => \N__20469\,
            I => \N__20454\
        );

    \I__3207\ : Sp12to4
    port map (
            O => \N__20466\,
            I => \N__20454\
        );

    \I__3206\ : Span4Mux_h
    port map (
            O => \N__20461\,
            I => \N__20451\
        );

    \I__3205\ : Odrv12
    port map (
            O => \N__20454\,
            I => \M_this_ppu_spr_addr_2\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__20451\,
            I => \M_this_ppu_spr_addr_2\
        );

    \I__3203\ : InMux
    port map (
            O => \N__20446\,
            I => \this_ppu.offset_x_cry_1\
        );

    \I__3202\ : InMux
    port map (
            O => \N__20443\,
            I => \N__20440\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__20440\,
            I => \this_ppu.M_oam_cache_read_data_i_11\
        );

    \I__3200\ : InMux
    port map (
            O => \N__20437\,
            I => \N__20434\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__20434\,
            I => \this_ppu.m68_0_o2_0\
        );

    \I__3198\ : InMux
    port map (
            O => \N__20431\,
            I => \this_ppu.offset_x_cry_2\
        );

    \I__3197\ : InMux
    port map (
            O => \N__20428\,
            I => \N__20425\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__20425\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__3195\ : InMux
    port map (
            O => \N__20422\,
            I => \N__20413\
        );

    \I__3194\ : InMux
    port map (
            O => \N__20421\,
            I => \N__20413\
        );

    \I__3193\ : InMux
    port map (
            O => \N__20420\,
            I => \N__20413\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__20413\,
            I => \N__20409\
        );

    \I__3191\ : InMux
    port map (
            O => \N__20412\,
            I => \N__20406\
        );

    \I__3190\ : Span4Mux_h
    port map (
            O => \N__20409\,
            I => \N__20403\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__20406\,
            I => \N__20400\
        );

    \I__3188\ : Span4Mux_v
    port map (
            O => \N__20403\,
            I => \N__20397\
        );

    \I__3187\ : Span12Mux_h
    port map (
            O => \N__20400\,
            I => \N__20394\
        );

    \I__3186\ : Span4Mux_v
    port map (
            O => \N__20397\,
            I => \N__20391\
        );

    \I__3185\ : Span12Mux_v
    port map (
            O => \N__20394\,
            I => \N__20388\
        );

    \I__3184\ : Span4Mux_v
    port map (
            O => \N__20391\,
            I => \N__20385\
        );

    \I__3183\ : Odrv12
    port map (
            O => \N__20388\,
            I => rst_n_c
        );

    \I__3182\ : Odrv4
    port map (
            O => \N__20385\,
            I => rst_n_c
        );

    \I__3181\ : InMux
    port map (
            O => \N__20380\,
            I => \N__20377\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__20377\,
            I => \N__20374\
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__20374\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__20371\,
            I => \N__20367\
        );

    \I__3177\ : CascadeMux
    port map (
            O => \N__20370\,
            I => \N__20363\
        );

    \I__3176\ : InMux
    port map (
            O => \N__20367\,
            I => \N__20360\
        );

    \I__3175\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20355\
        );

    \I__3174\ : InMux
    port map (
            O => \N__20363\,
            I => \N__20355\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__20360\,
            I => \this_vga_signals.N_1417\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__20355\,
            I => \this_vga_signals.N_1417\
        );

    \I__3171\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20347\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__20347\,
            I => \N__20343\
        );

    \I__3169\ : InMux
    port map (
            O => \N__20346\,
            I => \N__20338\
        );

    \I__3168\ : Span4Mux_v
    port map (
            O => \N__20343\,
            I => \N__20335\
        );

    \I__3167\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20332\
        );

    \I__3166\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20329\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__20338\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__20335\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__20332\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__20329\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__3161\ : InMux
    port map (
            O => \N__20320\,
            I => \N__20317\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__20317\,
            I => \N__20314\
        );

    \I__3159\ : Span12Mux_h
    port map (
            O => \N__20314\,
            I => \N__20311\
        );

    \I__3158\ : Odrv12
    port map (
            O => \N__20311\,
            I => \this_vga_ramdac.i2_mux_0\
        );

    \I__3157\ : InMux
    port map (
            O => \N__20308\,
            I => \N__20300\
        );

    \I__3156\ : InMux
    port map (
            O => \N__20307\,
            I => \N__20297\
        );

    \I__3155\ : InMux
    port map (
            O => \N__20306\,
            I => \N__20294\
        );

    \I__3154\ : InMux
    port map (
            O => \N__20305\,
            I => \N__20291\
        );

    \I__3153\ : InMux
    port map (
            O => \N__20304\,
            I => \N__20286\
        );

    \I__3152\ : InMux
    port map (
            O => \N__20303\,
            I => \N__20286\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__20300\,
            I => \N__20281\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__20297\,
            I => \N__20281\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__20294\,
            I => \M_pcounter_q_ret_1_RNIOILK7\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__20291\,
            I => \M_pcounter_q_ret_1_RNIOILK7\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__20286\,
            I => \M_pcounter_q_ret_1_RNIOILK7\
        );

    \I__3146\ : Odrv4
    port map (
            O => \N__20281\,
            I => \M_pcounter_q_ret_1_RNIOILK7\
        );

    \I__3145\ : InMux
    port map (
            O => \N__20272\,
            I => \N__20269\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__20269\,
            I => \N__20266\
        );

    \I__3143\ : Span4Mux_h
    port map (
            O => \N__20266\,
            I => \N__20262\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__20265\,
            I => \N__20259\
        );

    \I__3141\ : Span4Mux_h
    port map (
            O => \N__20262\,
            I => \N__20256\
        );

    \I__3140\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20253\
        );

    \I__3139\ : Odrv4
    port map (
            O => \N__20256\,
            I => \this_vga_ramdac.N_3861_reto\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__20253\,
            I => \this_vga_ramdac.N_3861_reto\
        );

    \I__3137\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20245\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__20245\,
            I => \N__20242\
        );

    \I__3135\ : Odrv12
    port map (
            O => \N__20242\,
            I => \this_ppu.un1_M_surface_x_q_ac0_11\
        );

    \I__3134\ : InMux
    port map (
            O => \N__20239\,
            I => \N__20236\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__20236\,
            I => \M_this_data_tmp_qZ0Z_12\
        );

    \I__3132\ : InMux
    port map (
            O => \N__20233\,
            I => \N__20230\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__20230\,
            I => \M_this_data_tmp_qZ0Z_14\
        );

    \I__3130\ : InMux
    port map (
            O => \N__20227\,
            I => \N__20224\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__20224\,
            I => \M_this_data_tmp_qZ0Z_1\
        );

    \I__3128\ : InMux
    port map (
            O => \N__20221\,
            I => \N__20218\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__20218\,
            I => \N__20215\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__20215\,
            I => \N__20212\
        );

    \I__3125\ : Span4Mux_h
    port map (
            O => \N__20212\,
            I => \N__20209\
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__20209\,
            I => \M_this_oam_ram_write_data_22\
        );

    \I__3123\ : InMux
    port map (
            O => \N__20206\,
            I => \N__20203\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__20203\,
            I => \M_this_data_tmp_qZ0Z_22\
        );

    \I__3121\ : InMux
    port map (
            O => \N__20200\,
            I => \N__20196\
        );

    \I__3120\ : InMux
    port map (
            O => \N__20199\,
            I => \N__20193\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__20196\,
            I => \N__20190\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__20193\,
            I => \N__20187\
        );

    \I__3117\ : Span12Mux_v
    port map (
            O => \N__20190\,
            I => \N__20184\
        );

    \I__3116\ : Span12Mux_h
    port map (
            O => \N__20187\,
            I => \N__20181\
        );

    \I__3115\ : Span12Mux_h
    port map (
            O => \N__20184\,
            I => \N__20178\
        );

    \I__3114\ : Odrv12
    port map (
            O => \N__20181\,
            I => \M_this_map_ram_read_data_1\
        );

    \I__3113\ : Odrv12
    port map (
            O => \N__20178\,
            I => \M_this_map_ram_read_data_1\
        );

    \I__3112\ : IoInMux
    port map (
            O => \N__20173\,
            I => \N__20170\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__20170\,
            I => \N__20167\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__20167\,
            I => \N_724_0\
        );

    \I__3109\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20161\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__20161\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__3107\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20155\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__20155\,
            I => \N__20152\
        );

    \I__3105\ : Span12Mux_h
    port map (
            O => \N__20152\,
            I => \N__20148\
        );

    \I__3104\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20145\
        );

    \I__3103\ : Odrv12
    port map (
            O => \N__20148\,
            I => \this_ppu.M_oam_cache_read_data_16\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__20145\,
            I => \this_ppu.M_oam_cache_read_data_16\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__20140\,
            I => \N__20136\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__20139\,
            I => \N__20133\
        );

    \I__3099\ : InMux
    port map (
            O => \N__20136\,
            I => \N__20125\
        );

    \I__3098\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20122\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__20132\,
            I => \N__20119\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__20131\,
            I => \N__20108\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__20130\,
            I => \N__20105\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__20129\,
            I => \N__20101\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__20128\,
            I => \N__20098\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__20125\,
            I => \N__20093\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__20122\,
            I => \N__20093\
        );

    \I__3090\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20090\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__20118\,
            I => \N__20087\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__20117\,
            I => \N__20084\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__20116\,
            I => \N__20081\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__20115\,
            I => \N__20078\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__20114\,
            I => \N__20075\
        );

    \I__3084\ : CascadeMux
    port map (
            O => \N__20113\,
            I => \N__20072\
        );

    \I__3083\ : CascadeMux
    port map (
            O => \N__20112\,
            I => \N__20069\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__20111\,
            I => \N__20066\
        );

    \I__3081\ : InMux
    port map (
            O => \N__20108\,
            I => \N__20063\
        );

    \I__3080\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20060\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__20104\,
            I => \N__20057\
        );

    \I__3078\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20054\
        );

    \I__3077\ : InMux
    port map (
            O => \N__20098\,
            I => \N__20051\
        );

    \I__3076\ : Span4Mux_v
    port map (
            O => \N__20093\,
            I => \N__20046\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__20090\,
            I => \N__20046\
        );

    \I__3074\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20043\
        );

    \I__3073\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20040\
        );

    \I__3072\ : InMux
    port map (
            O => \N__20081\,
            I => \N__20037\
        );

    \I__3071\ : InMux
    port map (
            O => \N__20078\,
            I => \N__20034\
        );

    \I__3070\ : InMux
    port map (
            O => \N__20075\,
            I => \N__20031\
        );

    \I__3069\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20028\
        );

    \I__3068\ : InMux
    port map (
            O => \N__20069\,
            I => \N__20025\
        );

    \I__3067\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20022\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__20063\,
            I => \N__20019\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__20060\,
            I => \N__20016\
        );

    \I__3064\ : InMux
    port map (
            O => \N__20057\,
            I => \N__20013\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__20054\,
            I => \N__20008\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__20051\,
            I => \N__20008\
        );

    \I__3061\ : Sp12to4
    port map (
            O => \N__20046\,
            I => \N__19997\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__20043\,
            I => \N__19997\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__20040\,
            I => \N__19997\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__20037\,
            I => \N__19997\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__20034\,
            I => \N__19997\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__20031\,
            I => \N__19988\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__20028\,
            I => \N__19988\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__20025\,
            I => \N__19988\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__20022\,
            I => \N__19988\
        );

    \I__3052\ : Span4Mux_s3_v
    port map (
            O => \N__20019\,
            I => \N__19981\
        );

    \I__3051\ : Span4Mux_h
    port map (
            O => \N__20016\,
            I => \N__19981\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__20013\,
            I => \N__19981\
        );

    \I__3049\ : Span12Mux_s11_v
    port map (
            O => \N__20008\,
            I => \N__19978\
        );

    \I__3048\ : Span12Mux_v
    port map (
            O => \N__19997\,
            I => \N__19975\
        );

    \I__3047\ : Span12Mux_v
    port map (
            O => \N__19988\,
            I => \N__19972\
        );

    \I__3046\ : Span4Mux_v
    port map (
            O => \N__19981\,
            I => \N__19969\
        );

    \I__3045\ : Span12Mux_h
    port map (
            O => \N__19978\,
            I => \N__19964\
        );

    \I__3044\ : Span12Mux_h
    port map (
            O => \N__19975\,
            I => \N__19964\
        );

    \I__3043\ : Span12Mux_h
    port map (
            O => \N__19972\,
            I => \N__19961\
        );

    \I__3042\ : Span4Mux_h
    port map (
            O => \N__19969\,
            I => \N__19958\
        );

    \I__3041\ : Odrv12
    port map (
            O => \N__19964\,
            I => \M_this_ppu_spr_addr_3\
        );

    \I__3040\ : Odrv12
    port map (
            O => \N__19961\,
            I => \M_this_ppu_spr_addr_3\
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__19958\,
            I => \M_this_ppu_spr_addr_3\
        );

    \I__3038\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19948\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__19948\,
            I => \N__19945\
        );

    \I__3036\ : Span4Mux_v
    port map (
            O => \N__19945\,
            I => \N__19942\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__19942\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_2\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__19939\,
            I => \N__19933\
        );

    \I__3033\ : CascadeMux
    port map (
            O => \N__19938\,
            I => \N__19930\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__19937\,
            I => \N__19925\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__19936\,
            I => \N__19919\
        );

    \I__3030\ : InMux
    port map (
            O => \N__19933\,
            I => \N__19915\
        );

    \I__3029\ : InMux
    port map (
            O => \N__19930\,
            I => \N__19912\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__19929\,
            I => \N__19909\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__19928\,
            I => \N__19906\
        );

    \I__3026\ : InMux
    port map (
            O => \N__19925\,
            I => \N__19902\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__19924\,
            I => \N__19899\
        );

    \I__3024\ : CascadeMux
    port map (
            O => \N__19923\,
            I => \N__19896\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__19922\,
            I => \N__19893\
        );

    \I__3022\ : InMux
    port map (
            O => \N__19919\,
            I => \N__19890\
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__19918\,
            I => \N__19887\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__19915\,
            I => \N__19882\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__19912\,
            I => \N__19879\
        );

    \I__3018\ : InMux
    port map (
            O => \N__19909\,
            I => \N__19876\
        );

    \I__3017\ : InMux
    port map (
            O => \N__19906\,
            I => \N__19873\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__19905\,
            I => \N__19870\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__19902\,
            I => \N__19866\
        );

    \I__3014\ : InMux
    port map (
            O => \N__19899\,
            I => \N__19863\
        );

    \I__3013\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19860\
        );

    \I__3012\ : InMux
    port map (
            O => \N__19893\,
            I => \N__19857\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__19890\,
            I => \N__19854\
        );

    \I__3010\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19851\
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__19886\,
            I => \N__19848\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__19885\,
            I => \N__19845\
        );

    \I__3007\ : Span4Mux_v
    port map (
            O => \N__19882\,
            I => \N__19836\
        );

    \I__3006\ : Span4Mux_v
    port map (
            O => \N__19879\,
            I => \N__19836\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__19876\,
            I => \N__19836\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__19873\,
            I => \N__19833\
        );

    \I__3003\ : InMux
    port map (
            O => \N__19870\,
            I => \N__19830\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__19869\,
            I => \N__19827\
        );

    \I__3001\ : Span4Mux_v
    port map (
            O => \N__19866\,
            I => \N__19822\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__19863\,
            I => \N__19822\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__19860\,
            I => \N__19819\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__19857\,
            I => \N__19816\
        );

    \I__2997\ : Span4Mux_v
    port map (
            O => \N__19854\,
            I => \N__19811\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__19851\,
            I => \N__19811\
        );

    \I__2995\ : InMux
    port map (
            O => \N__19848\,
            I => \N__19808\
        );

    \I__2994\ : InMux
    port map (
            O => \N__19845\,
            I => \N__19805\
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__19844\,
            I => \N__19802\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__19843\,
            I => \N__19799\
        );

    \I__2991\ : Span4Mux_v
    port map (
            O => \N__19836\,
            I => \N__19792\
        );

    \I__2990\ : Span4Mux_h
    port map (
            O => \N__19833\,
            I => \N__19792\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__19830\,
            I => \N__19792\
        );

    \I__2988\ : InMux
    port map (
            O => \N__19827\,
            I => \N__19789\
        );

    \I__2987\ : Span4Mux_h
    port map (
            O => \N__19822\,
            I => \N__19786\
        );

    \I__2986\ : Span4Mux_v
    port map (
            O => \N__19819\,
            I => \N__19777\
        );

    \I__2985\ : Span4Mux_v
    port map (
            O => \N__19816\,
            I => \N__19777\
        );

    \I__2984\ : Span4Mux_v
    port map (
            O => \N__19811\,
            I => \N__19777\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__19808\,
            I => \N__19777\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__19805\,
            I => \N__19774\
        );

    \I__2981\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19771\
        );

    \I__2980\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19768\
        );

    \I__2979\ : Span4Mux_v
    port map (
            O => \N__19792\,
            I => \N__19765\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__19789\,
            I => \N__19762\
        );

    \I__2977\ : Span4Mux_v
    port map (
            O => \N__19786\,
            I => \N__19757\
        );

    \I__2976\ : Span4Mux_h
    port map (
            O => \N__19777\,
            I => \N__19757\
        );

    \I__2975\ : Span4Mux_s3_v
    port map (
            O => \N__19774\,
            I => \N__19750\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__19771\,
            I => \N__19750\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__19768\,
            I => \N__19750\
        );

    \I__2972\ : Sp12to4
    port map (
            O => \N__19765\,
            I => \N__19745\
        );

    \I__2971\ : Span12Mux_s7_h
    port map (
            O => \N__19762\,
            I => \N__19745\
        );

    \I__2970\ : Span4Mux_h
    port map (
            O => \N__19757\,
            I => \N__19742\
        );

    \I__2969\ : Span4Mux_v
    port map (
            O => \N__19750\,
            I => \N__19739\
        );

    \I__2968\ : Span12Mux_h
    port map (
            O => \N__19745\,
            I => \N__19736\
        );

    \I__2967\ : Span4Mux_h
    port map (
            O => \N__19742\,
            I => \N__19733\
        );

    \I__2966\ : Span4Mux_h
    port map (
            O => \N__19739\,
            I => \N__19730\
        );

    \I__2965\ : Odrv12
    port map (
            O => \N__19736\,
            I => \read_data_RNI6RFJ1_2\
        );

    \I__2964\ : Odrv4
    port map (
            O => \N__19733\,
            I => \read_data_RNI6RFJ1_2\
        );

    \I__2963\ : Odrv4
    port map (
            O => \N__19730\,
            I => \read_data_RNI6RFJ1_2\
        );

    \I__2962\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19720\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__19720\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_3\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__19717\,
            I => \N__19710\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__19716\,
            I => \N__19706\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__19715\,
            I => \N__19701\
        );

    \I__2957\ : CascadeMux
    port map (
            O => \N__19714\,
            I => \N__19698\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__19713\,
            I => \N__19695\
        );

    \I__2955\ : InMux
    port map (
            O => \N__19710\,
            I => \N__19689\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__19709\,
            I => \N__19686\
        );

    \I__2953\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19678\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__19705\,
            I => \N__19675\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__19704\,
            I => \N__19672\
        );

    \I__2950\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19669\
        );

    \I__2949\ : InMux
    port map (
            O => \N__19698\,
            I => \N__19666\
        );

    \I__2948\ : InMux
    port map (
            O => \N__19695\,
            I => \N__19663\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__19694\,
            I => \N__19660\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__19693\,
            I => \N__19657\
        );

    \I__2945\ : CascadeMux
    port map (
            O => \N__19692\,
            I => \N__19654\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__19689\,
            I => \N__19651\
        );

    \I__2943\ : InMux
    port map (
            O => \N__19686\,
            I => \N__19648\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__19685\,
            I => \N__19645\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__19684\,
            I => \N__19642\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__19683\,
            I => \N__19639\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__19682\,
            I => \N__19636\
        );

    \I__2938\ : CascadeMux
    port map (
            O => \N__19681\,
            I => \N__19633\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__19678\,
            I => \N__19630\
        );

    \I__2936\ : InMux
    port map (
            O => \N__19675\,
            I => \N__19627\
        );

    \I__2935\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19624\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__19669\,
            I => \N__19617\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__19666\,
            I => \N__19617\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__19663\,
            I => \N__19617\
        );

    \I__2931\ : InMux
    port map (
            O => \N__19660\,
            I => \N__19614\
        );

    \I__2930\ : InMux
    port map (
            O => \N__19657\,
            I => \N__19611\
        );

    \I__2929\ : InMux
    port map (
            O => \N__19654\,
            I => \N__19608\
        );

    \I__2928\ : Span4Mux_v
    port map (
            O => \N__19651\,
            I => \N__19603\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__19648\,
            I => \N__19603\
        );

    \I__2926\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19600\
        );

    \I__2925\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19597\
        );

    \I__2924\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19594\
        );

    \I__2923\ : InMux
    port map (
            O => \N__19636\,
            I => \N__19591\
        );

    \I__2922\ : InMux
    port map (
            O => \N__19633\,
            I => \N__19588\
        );

    \I__2921\ : Span4Mux_s3_v
    port map (
            O => \N__19630\,
            I => \N__19581\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__19627\,
            I => \N__19581\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__19624\,
            I => \N__19581\
        );

    \I__2918\ : Span12Mux_v
    port map (
            O => \N__19617\,
            I => \N__19578\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__19614\,
            I => \N__19571\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__19611\,
            I => \N__19571\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__19608\,
            I => \N__19571\
        );

    \I__2914\ : Sp12to4
    port map (
            O => \N__19603\,
            I => \N__19558\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__19600\,
            I => \N__19558\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__19597\,
            I => \N__19558\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__19594\,
            I => \N__19558\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__19591\,
            I => \N__19558\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__19588\,
            I => \N__19558\
        );

    \I__2908\ : Span4Mux_v
    port map (
            O => \N__19581\,
            I => \N__19555\
        );

    \I__2907\ : Span12Mux_h
    port map (
            O => \N__19578\,
            I => \N__19552\
        );

    \I__2906\ : Span12Mux_s10_v
    port map (
            O => \N__19571\,
            I => \N__19547\
        );

    \I__2905\ : Span12Mux_v
    port map (
            O => \N__19558\,
            I => \N__19547\
        );

    \I__2904\ : Span4Mux_h
    port map (
            O => \N__19555\,
            I => \N__19544\
        );

    \I__2903\ : Odrv12
    port map (
            O => \N__19552\,
            I => \read_data_RNI7SFJ1_3\
        );

    \I__2902\ : Odrv12
    port map (
            O => \N__19547\,
            I => \read_data_RNI7SFJ1_3\
        );

    \I__2901\ : Odrv4
    port map (
            O => \N__19544\,
            I => \read_data_RNI7SFJ1_3\
        );

    \I__2900\ : InMux
    port map (
            O => \N__19537\,
            I => \N__19534\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__19534\,
            I => \N__19531\
        );

    \I__2898\ : Span4Mux_h
    port map (
            O => \N__19531\,
            I => \N__19528\
        );

    \I__2897\ : Span4Mux_v
    port map (
            O => \N__19528\,
            I => \N__19525\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__19525\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_4\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__19522\,
            I => \N__19519\
        );

    \I__2894\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19513\
        );

    \I__2893\ : CascadeMux
    port map (
            O => \N__19518\,
            I => \N__19510\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__19517\,
            I => \N__19505\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__19516\,
            I => \N__19502\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__19513\,
            I => \N__19493\
        );

    \I__2889\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19490\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__19509\,
            I => \N__19487\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__19508\,
            I => \N__19482\
        );

    \I__2886\ : InMux
    port map (
            O => \N__19505\,
            I => \N__19477\
        );

    \I__2885\ : InMux
    port map (
            O => \N__19502\,
            I => \N__19474\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__19501\,
            I => \N__19471\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__19500\,
            I => \N__19468\
        );

    \I__2882\ : CascadeMux
    port map (
            O => \N__19499\,
            I => \N__19465\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__19498\,
            I => \N__19462\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__19497\,
            I => \N__19459\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__19496\,
            I => \N__19456\
        );

    \I__2878\ : Span4Mux_v
    port map (
            O => \N__19493\,
            I => \N__19451\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__19490\,
            I => \N__19451\
        );

    \I__2876\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19448\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__19486\,
            I => \N__19445\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__19485\,
            I => \N__19442\
        );

    \I__2873\ : InMux
    port map (
            O => \N__19482\,
            I => \N__19439\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__19481\,
            I => \N__19436\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__19480\,
            I => \N__19433\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__19477\,
            I => \N__19430\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__19474\,
            I => \N__19427\
        );

    \I__2868\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19424\
        );

    \I__2867\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19421\
        );

    \I__2866\ : InMux
    port map (
            O => \N__19465\,
            I => \N__19418\
        );

    \I__2865\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19415\
        );

    \I__2864\ : InMux
    port map (
            O => \N__19459\,
            I => \N__19412\
        );

    \I__2863\ : InMux
    port map (
            O => \N__19456\,
            I => \N__19409\
        );

    \I__2862\ : Span4Mux_v
    port map (
            O => \N__19451\,
            I => \N__19404\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__19448\,
            I => \N__19404\
        );

    \I__2860\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19401\
        );

    \I__2859\ : InMux
    port map (
            O => \N__19442\,
            I => \N__19398\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__19439\,
            I => \N__19395\
        );

    \I__2857\ : InMux
    port map (
            O => \N__19436\,
            I => \N__19392\
        );

    \I__2856\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19389\
        );

    \I__2855\ : Span12Mux_s4_v
    port map (
            O => \N__19430\,
            I => \N__19384\
        );

    \I__2854\ : Span12Mux_s7_h
    port map (
            O => \N__19427\,
            I => \N__19384\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__19424\,
            I => \N__19377\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__19421\,
            I => \N__19377\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__19418\,
            I => \N__19377\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__19415\,
            I => \N__19374\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__19412\,
            I => \N__19363\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__19409\,
            I => \N__19363\
        );

    \I__2847\ : Sp12to4
    port map (
            O => \N__19404\,
            I => \N__19363\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__19401\,
            I => \N__19363\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__19398\,
            I => \N__19363\
        );

    \I__2844\ : Span4Mux_s3_v
    port map (
            O => \N__19395\,
            I => \N__19358\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__19392\,
            I => \N__19358\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__19389\,
            I => \N__19355\
        );

    \I__2841\ : Span12Mux_h
    port map (
            O => \N__19384\,
            I => \N__19352\
        );

    \I__2840\ : Span12Mux_v
    port map (
            O => \N__19377\,
            I => \N__19345\
        );

    \I__2839\ : Sp12to4
    port map (
            O => \N__19374\,
            I => \N__19345\
        );

    \I__2838\ : Span12Mux_v
    port map (
            O => \N__19363\,
            I => \N__19345\
        );

    \I__2837\ : Span4Mux_v
    port map (
            O => \N__19358\,
            I => \N__19340\
        );

    \I__2836\ : Span4Mux_v
    port map (
            O => \N__19355\,
            I => \N__19340\
        );

    \I__2835\ : Span12Mux_v
    port map (
            O => \N__19352\,
            I => \N__19335\
        );

    \I__2834\ : Span12Mux_h
    port map (
            O => \N__19345\,
            I => \N__19335\
        );

    \I__2833\ : Span4Mux_h
    port map (
            O => \N__19340\,
            I => \N__19332\
        );

    \I__2832\ : Odrv12
    port map (
            O => \N__19335\,
            I => \read_data_RNI9TFJ1_4\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__19332\,
            I => \read_data_RNI9TFJ1_4\
        );

    \I__2830\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19324\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__19324\,
            I => \N__19321\
        );

    \I__2828\ : Span4Mux_v
    port map (
            O => \N__19321\,
            I => \N__19318\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__19318\,
            I => \this_vga_signals.M_pcounter_q_0Z0Z_1\
        );

    \I__2826\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19312\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__19312\,
            I => \N__19309\
        );

    \I__2824\ : Span4Mux_v
    port map (
            O => \N__19309\,
            I => \N__19306\
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__19306\,
            I => \M_this_data_tmp_qZ0Z_11\
        );

    \I__2822\ : InMux
    port map (
            O => \N__19303\,
            I => \N__19300\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__19300\,
            I => \N__19297\
        );

    \I__2820\ : Odrv12
    port map (
            O => \N__19297\,
            I => \M_this_oam_ram_write_data_11\
        );

    \I__2819\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19291\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__19291\,
            I => \N__19288\
        );

    \I__2817\ : Odrv12
    port map (
            O => \N__19288\,
            I => \M_this_oam_ram_write_data_12\
        );

    \I__2816\ : InMux
    port map (
            O => \N__19285\,
            I => \N__19282\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__19282\,
            I => \N__19279\
        );

    \I__2814\ : Odrv12
    port map (
            O => \N__19279\,
            I => \M_this_oam_ram_write_data_13\
        );

    \I__2813\ : InMux
    port map (
            O => \N__19276\,
            I => \N__19273\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__19273\,
            I => \N__19270\
        );

    \I__2811\ : Odrv12
    port map (
            O => \N__19270\,
            I => \M_this_oam_ram_write_data_14\
        );

    \I__2810\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19264\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__19264\,
            I => \N__19260\
        );

    \I__2808\ : InMux
    port map (
            O => \N__19263\,
            I => \N__19257\
        );

    \I__2807\ : Span4Mux_v
    port map (
            O => \N__19260\,
            I => \N__19251\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__19257\,
            I => \N__19251\
        );

    \I__2805\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19248\
        );

    \I__2804\ : Span4Mux_v
    port map (
            O => \N__19251\,
            I => \N__19245\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__19248\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__2802\ : Odrv4
    port map (
            O => \N__19245\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__2801\ : InMux
    port map (
            O => \N__19240\,
            I => \N__19236\
        );

    \I__2800\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19233\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__19236\,
            I => \N__19230\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__19233\,
            I => \this_pixel_clk_M_counter_q_i_1\
        );

    \I__2797\ : Odrv12
    port map (
            O => \N__19230\,
            I => \this_pixel_clk_M_counter_q_i_1\
        );

    \I__2796\ : InMux
    port map (
            O => \N__19225\,
            I => \N__19217\
        );

    \I__2795\ : CascadeMux
    port map (
            O => \N__19224\,
            I => \N__19212\
        );

    \I__2794\ : InMux
    port map (
            O => \N__19223\,
            I => \N__19206\
        );

    \I__2793\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19201\
        );

    \I__2792\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19201\
        );

    \I__2791\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19198\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__19217\,
            I => \N__19195\
        );

    \I__2789\ : InMux
    port map (
            O => \N__19216\,
            I => \N__19192\
        );

    \I__2788\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19189\
        );

    \I__2787\ : InMux
    port map (
            O => \N__19212\,
            I => \N__19186\
        );

    \I__2786\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19183\
        );

    \I__2785\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19178\
        );

    \I__2784\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19178\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__19206\,
            I => \N__19171\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__19201\,
            I => \N__19171\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__19198\,
            I => \N__19171\
        );

    \I__2780\ : Span4Mux_h
    port map (
            O => \N__19195\,
            I => \N__19164\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__19192\,
            I => \N__19164\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__19189\,
            I => \N__19164\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__19186\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__19183\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__19178\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2774\ : Odrv4
    port map (
            O => \N__19171\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2773\ : Odrv4
    port map (
            O => \N__19164\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2772\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19146\
        );

    \I__2771\ : InMux
    port map (
            O => \N__19152\,
            I => \N__19143\
        );

    \I__2770\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19138\
        );

    \I__2769\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19138\
        );

    \I__2768\ : InMux
    port map (
            O => \N__19149\,
            I => \N__19135\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__19146\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__19143\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__19138\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__19135\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\
        );

    \I__2763\ : InMux
    port map (
            O => \N__19126\,
            I => \N__19115\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__19125\,
            I => \N__19112\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__19124\,
            I => \N__19109\
        );

    \I__2760\ : InMux
    port map (
            O => \N__19123\,
            I => \N__19101\
        );

    \I__2759\ : InMux
    port map (
            O => \N__19122\,
            I => \N__19101\
        );

    \I__2758\ : InMux
    port map (
            O => \N__19121\,
            I => \N__19101\
        );

    \I__2757\ : InMux
    port map (
            O => \N__19120\,
            I => \N__19098\
        );

    \I__2756\ : InMux
    port map (
            O => \N__19119\,
            I => \N__19095\
        );

    \I__2755\ : InMux
    port map (
            O => \N__19118\,
            I => \N__19092\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__19115\,
            I => \N__19089\
        );

    \I__2753\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19086\
        );

    \I__2752\ : InMux
    port map (
            O => \N__19109\,
            I => \N__19083\
        );

    \I__2751\ : InMux
    port map (
            O => \N__19108\,
            I => \N__19080\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__19101\,
            I => \N__19073\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__19098\,
            I => \N__19073\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__19095\,
            I => \N__19073\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__19092\,
            I => \N__19067\
        );

    \I__2746\ : Span4Mux_v
    port map (
            O => \N__19089\,
            I => \N__19067\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__19086\,
            I => \N__19064\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__19083\,
            I => \N__19059\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__19080\,
            I => \N__19059\
        );

    \I__2742\ : Span4Mux_h
    port map (
            O => \N__19073\,
            I => \N__19056\
        );

    \I__2741\ : InMux
    port map (
            O => \N__19072\,
            I => \N__19053\
        );

    \I__2740\ : Odrv4
    port map (
            O => \N__19067\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2739\ : Odrv12
    port map (
            O => \N__19064\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2738\ : Odrv4
    port map (
            O => \N__19059\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2737\ : Odrv4
    port map (
            O => \N__19056\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__19053\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2735\ : InMux
    port map (
            O => \N__19042\,
            I => \N__19038\
        );

    \I__2734\ : InMux
    port map (
            O => \N__19041\,
            I => \N__19035\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__19038\,
            I => \N__19031\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__19035\,
            I => \N__19024\
        );

    \I__2731\ : InMux
    port map (
            O => \N__19034\,
            I => \N__19021\
        );

    \I__2730\ : Span4Mux_h
    port map (
            O => \N__19031\,
            I => \N__19018\
        );

    \I__2729\ : InMux
    port map (
            O => \N__19030\,
            I => \N__19015\
        );

    \I__2728\ : InMux
    port map (
            O => \N__19029\,
            I => \N__19008\
        );

    \I__2727\ : InMux
    port map (
            O => \N__19028\,
            I => \N__19008\
        );

    \I__2726\ : InMux
    port map (
            O => \N__19027\,
            I => \N__19008\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__19024\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_3\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__19021\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_3\
        );

    \I__2723\ : Odrv4
    port map (
            O => \N__19018\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_3\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__19015\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_3\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__19008\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_3\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__18997\,
            I => \N__18993\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__18996\,
            I => \N__18990\
        );

    \I__2718\ : InMux
    port map (
            O => \N__18993\,
            I => \N__18985\
        );

    \I__2717\ : InMux
    port map (
            O => \N__18990\,
            I => \N__18985\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__18985\,
            I => \N__18982\
        );

    \I__2715\ : Odrv4
    port map (
            O => \N__18982\,
            I => \this_vga_signals.M_hcounter_q_RNII1437Z0Z_3\
        );

    \I__2714\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18976\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__18976\,
            I => \N__18973\
        );

    \I__2712\ : Span4Mux_h
    port map (
            O => \N__18973\,
            I => \N__18970\
        );

    \I__2711\ : Span4Mux_h
    port map (
            O => \N__18970\,
            I => \N__18967\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__18967\,
            I => \M_this_oam_ram_read_data_30\
        );

    \I__2709\ : InMux
    port map (
            O => \N__18964\,
            I => \N__18961\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__18961\,
            I => \N__18958\
        );

    \I__2707\ : Span4Mux_h
    port map (
            O => \N__18958\,
            I => \N__18955\
        );

    \I__2706\ : Span4Mux_h
    port map (
            O => \N__18955\,
            I => \N__18952\
        );

    \I__2705\ : Odrv4
    port map (
            O => \N__18952\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_30\
        );

    \I__2704\ : InMux
    port map (
            O => \N__18949\,
            I => \N__18946\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__18946\,
            I => \N__18943\
        );

    \I__2702\ : Span4Mux_h
    port map (
            O => \N__18943\,
            I => \N__18940\
        );

    \I__2701\ : Span4Mux_h
    port map (
            O => \N__18940\,
            I => \N__18937\
        );

    \I__2700\ : Odrv4
    port map (
            O => \N__18937\,
            I => \this_ppu.oam_cache.mem_3\
        );

    \I__2699\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18931\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__18931\,
            I => \N__18928\
        );

    \I__2697\ : Span4Mux_v
    port map (
            O => \N__18928\,
            I => \N__18925\
        );

    \I__2696\ : Odrv4
    port map (
            O => \N__18925\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_1\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__18922\,
            I => \N__18918\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__18921\,
            I => \N__18913\
        );

    \I__2693\ : InMux
    port map (
            O => \N__18918\,
            I => \N__18910\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__18917\,
            I => \N__18907\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__18916\,
            I => \N__18900\
        );

    \I__2690\ : InMux
    port map (
            O => \N__18913\,
            I => \N__18891\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__18910\,
            I => \N__18888\
        );

    \I__2688\ : InMux
    port map (
            O => \N__18907\,
            I => \N__18885\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__18906\,
            I => \N__18882\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__18905\,
            I => \N__18879\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__18904\,
            I => \N__18876\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__18903\,
            I => \N__18873\
        );

    \I__2683\ : InMux
    port map (
            O => \N__18900\,
            I => \N__18870\
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__18899\,
            I => \N__18867\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__18898\,
            I => \N__18864\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__18897\,
            I => \N__18861\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__18896\,
            I => \N__18858\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__18895\,
            I => \N__18855\
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__18894\,
            I => \N__18851\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__18891\,
            I => \N__18847\
        );

    \I__2675\ : Span4Mux_v
    port map (
            O => \N__18888\,
            I => \N__18844\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__18885\,
            I => \N__18841\
        );

    \I__2673\ : InMux
    port map (
            O => \N__18882\,
            I => \N__18838\
        );

    \I__2672\ : InMux
    port map (
            O => \N__18879\,
            I => \N__18835\
        );

    \I__2671\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18832\
        );

    \I__2670\ : InMux
    port map (
            O => \N__18873\,
            I => \N__18829\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__18870\,
            I => \N__18826\
        );

    \I__2668\ : InMux
    port map (
            O => \N__18867\,
            I => \N__18823\
        );

    \I__2667\ : InMux
    port map (
            O => \N__18864\,
            I => \N__18820\
        );

    \I__2666\ : InMux
    port map (
            O => \N__18861\,
            I => \N__18817\
        );

    \I__2665\ : InMux
    port map (
            O => \N__18858\,
            I => \N__18814\
        );

    \I__2664\ : InMux
    port map (
            O => \N__18855\,
            I => \N__18811\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__18854\,
            I => \N__18808\
        );

    \I__2662\ : InMux
    port map (
            O => \N__18851\,
            I => \N__18805\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__18850\,
            I => \N__18802\
        );

    \I__2660\ : Span12Mux_s6_v
    port map (
            O => \N__18847\,
            I => \N__18795\
        );

    \I__2659\ : Sp12to4
    port map (
            O => \N__18844\,
            I => \N__18795\
        );

    \I__2658\ : Span12Mux_s7_h
    port map (
            O => \N__18841\,
            I => \N__18795\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__18838\,
            I => \N__18786\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__18835\,
            I => \N__18786\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__18832\,
            I => \N__18786\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__18829\,
            I => \N__18786\
        );

    \I__2653\ : Span4Mux_v
    port map (
            O => \N__18826\,
            I => \N__18783\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__18823\,
            I => \N__18780\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__18820\,
            I => \N__18771\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__18817\,
            I => \N__18771\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__18814\,
            I => \N__18771\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__18811\,
            I => \N__18771\
        );

    \I__2647\ : InMux
    port map (
            O => \N__18808\,
            I => \N__18768\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__18805\,
            I => \N__18765\
        );

    \I__2645\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18762\
        );

    \I__2644\ : Span12Mux_h
    port map (
            O => \N__18795\,
            I => \N__18759\
        );

    \I__2643\ : Span12Mux_v
    port map (
            O => \N__18786\,
            I => \N__18750\
        );

    \I__2642\ : Sp12to4
    port map (
            O => \N__18783\,
            I => \N__18750\
        );

    \I__2641\ : Sp12to4
    port map (
            O => \N__18780\,
            I => \N__18750\
        );

    \I__2640\ : Span12Mux_v
    port map (
            O => \N__18771\,
            I => \N__18750\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__18768\,
            I => \N__18743\
        );

    \I__2638\ : Sp12to4
    port map (
            O => \N__18765\,
            I => \N__18743\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__18762\,
            I => \N__18743\
        );

    \I__2636\ : Span12Mux_v
    port map (
            O => \N__18759\,
            I => \N__18738\
        );

    \I__2635\ : Span12Mux_h
    port map (
            O => \N__18750\,
            I => \N__18738\
        );

    \I__2634\ : Span12Mux_s10_v
    port map (
            O => \N__18743\,
            I => \N__18735\
        );

    \I__2633\ : Odrv12
    port map (
            O => \N__18738\,
            I => \read_data_RNI5QFJ1_1\
        );

    \I__2632\ : Odrv12
    port map (
            O => \N__18735\,
            I => \read_data_RNI5QFJ1_1\
        );

    \I__2631\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18726\
        );

    \I__2630\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18723\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__18726\,
            I => \N__18718\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__18723\,
            I => \N__18718\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__18718\,
            I => \this_ppu.N_1196_1\
        );

    \I__2626\ : InMux
    port map (
            O => \N__18715\,
            I => \N__18708\
        );

    \I__2625\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18708\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__18713\,
            I => \N__18705\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__18708\,
            I => \N__18702\
        );

    \I__2622\ : InMux
    port map (
            O => \N__18705\,
            I => \N__18699\
        );

    \I__2621\ : Span4Mux_h
    port map (
            O => \N__18702\,
            I => \N__18696\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__18699\,
            I => \this_ppu.M_oam_curr_qZ0Z_6\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__18696\,
            I => \this_ppu.M_oam_curr_qZ0Z_6\
        );

    \I__2618\ : InMux
    port map (
            O => \N__18691\,
            I => \N__18688\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__18688\,
            I => \N__18685\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__18685\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_13\
        );

    \I__2615\ : SRMux
    port map (
            O => \N__18682\,
            I => \N__18678\
        );

    \I__2614\ : SRMux
    port map (
            O => \N__18681\,
            I => \N__18675\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__18678\,
            I => \N__18671\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__18675\,
            I => \N__18668\
        );

    \I__2611\ : SRMux
    port map (
            O => \N__18674\,
            I => \N__18665\
        );

    \I__2610\ : Span4Mux_v
    port map (
            O => \N__18671\,
            I => \N__18658\
        );

    \I__2609\ : Span4Mux_h
    port map (
            O => \N__18668\,
            I => \N__18658\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__18665\,
            I => \N__18658\
        );

    \I__2607\ : Sp12to4
    port map (
            O => \N__18658\,
            I => \N__18655\
        );

    \I__2606\ : Odrv12
    port map (
            O => \N__18655\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIRSG13Z0Z_9\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__18652\,
            I => \this_vga_signals.M_hcounter_q_esr_RNIRSG13Z0Z_9_cascade_\
        );

    \I__2604\ : CEMux
    port map (
            O => \N__18649\,
            I => \N__18646\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__18646\,
            I => \this_vga_signals.N_1307_1\
        );

    \I__2602\ : InMux
    port map (
            O => \N__18643\,
            I => \N__18640\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__18640\,
            I => \N__18637\
        );

    \I__2600\ : Span4Mux_h
    port map (
            O => \N__18637\,
            I => \N__18634\
        );

    \I__2599\ : Span4Mux_h
    port map (
            O => \N__18634\,
            I => \N__18631\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__18631\,
            I => \this_ppu.oam_cache.mem_8\
        );

    \I__2597\ : InMux
    port map (
            O => \N__18628\,
            I => \N__18625\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__18625\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_11\
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__18622\,
            I => \N__18615\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__18621\,
            I => \N__18611\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__18620\,
            I => \N__18607\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__18619\,
            I => \N__18604\
        );

    \I__2591\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18600\
        );

    \I__2590\ : InMux
    port map (
            O => \N__18615\,
            I => \N__18595\
        );

    \I__2589\ : InMux
    port map (
            O => \N__18614\,
            I => \N__18595\
        );

    \I__2588\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18589\
        );

    \I__2587\ : InMux
    port map (
            O => \N__18610\,
            I => \N__18589\
        );

    \I__2586\ : InMux
    port map (
            O => \N__18607\,
            I => \N__18586\
        );

    \I__2585\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18583\
        );

    \I__2584\ : InMux
    port map (
            O => \N__18603\,
            I => \N__18580\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__18600\,
            I => \N__18577\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__18595\,
            I => \N__18574\
        );

    \I__2581\ : InMux
    port map (
            O => \N__18594\,
            I => \N__18571\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__18589\,
            I => \N__18568\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__18586\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__18583\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__18580\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__18577\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2575\ : Odrv12
    port map (
            O => \N__18574\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__18571\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2573\ : Odrv4
    port map (
            O => \N__18568\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2572\ : InMux
    port map (
            O => \N__18553\,
            I => \N__18550\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__18550\,
            I => \N__18546\
        );

    \I__2570\ : InMux
    port map (
            O => \N__18549\,
            I => \N__18543\
        );

    \I__2569\ : Odrv4
    port map (
            O => \N__18546\,
            I => \this_vga_signals.mult1_un61_sum_axbxc1_0\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__18543\,
            I => \this_vga_signals.mult1_un61_sum_axbxc1_0\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__18538\,
            I => \this_vga_signals.N_2_0_cascade_\
        );

    \I__2566\ : InMux
    port map (
            O => \N__18535\,
            I => \N__18532\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__18532\,
            I => \N__18529\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__18529\,
            I => \this_vga_ramdac.m19\
        );

    \I__2563\ : InMux
    port map (
            O => \N__18526\,
            I => \N__18522\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__18525\,
            I => \N__18519\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__18522\,
            I => \N__18516\
        );

    \I__2560\ : InMux
    port map (
            O => \N__18519\,
            I => \N__18513\
        );

    \I__2559\ : Odrv12
    port map (
            O => \N__18516\,
            I => \this_vga_ramdac.N_3860_reto\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__18513\,
            I => \this_vga_ramdac.N_3860_reto\
        );

    \I__2557\ : InMux
    port map (
            O => \N__18508\,
            I => \N__18505\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__18505\,
            I => \N__18502\
        );

    \I__2555\ : Span12Mux_h
    port map (
            O => \N__18502\,
            I => \N__18499\
        );

    \I__2554\ : Odrv12
    port map (
            O => \N__18499\,
            I => \this_ppu.oam_cache.mem_14\
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__18496\,
            I => \this_ppu.m35_i_0_a3_0_cascade_\
        );

    \I__2552\ : InMux
    port map (
            O => \N__18493\,
            I => \N__18490\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__18490\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_9\
        );

    \I__2550\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18484\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__18484\,
            I => \N__18481\
        );

    \I__2548\ : Span4Mux_v
    port map (
            O => \N__18481\,
            I => \N__18478\
        );

    \I__2547\ : Span4Mux_h
    port map (
            O => \N__18478\,
            I => \N__18475\
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__18475\,
            I => \this_ppu.oam_cache.mem_11\
        );

    \I__2545\ : InMux
    port map (
            O => \N__18472\,
            I => \N__18469\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__18469\,
            I => \N__18466\
        );

    \I__2543\ : Span4Mux_h
    port map (
            O => \N__18466\,
            I => \N__18463\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__18463\,
            I => \this_ppu.oam_cache.mem_1\
        );

    \I__2541\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18457\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__18457\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_14\
        );

    \I__2539\ : InMux
    port map (
            O => \N__18454\,
            I => \N__18451\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__18451\,
            I => \this_vga_ramdac.N_24_mux\
        );

    \I__2537\ : InMux
    port map (
            O => \N__18448\,
            I => \N__18439\
        );

    \I__2536\ : InMux
    port map (
            O => \N__18447\,
            I => \N__18439\
        );

    \I__2535\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18439\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__18439\,
            I => \N__18434\
        );

    \I__2533\ : InMux
    port map (
            O => \N__18438\,
            I => \N__18429\
        );

    \I__2532\ : InMux
    port map (
            O => \N__18437\,
            I => \N__18429\
        );

    \I__2531\ : Span4Mux_v
    port map (
            O => \N__18434\,
            I => \N__18423\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__18429\,
            I => \N__18423\
        );

    \I__2529\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18420\
        );

    \I__2528\ : Span4Mux_h
    port map (
            O => \N__18423\,
            I => \N__18415\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__18420\,
            I => \N__18415\
        );

    \I__2526\ : Span4Mux_v
    port map (
            O => \N__18415\,
            I => \N__18412\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__18412\,
            I => \M_this_vram_read_data_0\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__18409\,
            I => \N__18405\
        );

    \I__2523\ : InMux
    port map (
            O => \N__18408\,
            I => \N__18399\
        );

    \I__2522\ : InMux
    port map (
            O => \N__18405\,
            I => \N__18399\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__18404\,
            I => \N__18395\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__18399\,
            I => \N__18391\
        );

    \I__2519\ : InMux
    port map (
            O => \N__18398\,
            I => \N__18386\
        );

    \I__2518\ : InMux
    port map (
            O => \N__18395\,
            I => \N__18386\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__18394\,
            I => \N__18383\
        );

    \I__2516\ : Span4Mux_h
    port map (
            O => \N__18391\,
            I => \N__18380\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__18386\,
            I => \N__18377\
        );

    \I__2514\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18374\
        );

    \I__2513\ : Span4Mux_h
    port map (
            O => \N__18380\,
            I => \N__18371\
        );

    \I__2512\ : Span4Mux_v
    port map (
            O => \N__18377\,
            I => \N__18366\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__18374\,
            I => \N__18366\
        );

    \I__2510\ : Span4Mux_v
    port map (
            O => \N__18371\,
            I => \N__18363\
        );

    \I__2509\ : Span4Mux_h
    port map (
            O => \N__18366\,
            I => \N__18360\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__18363\,
            I => \M_this_vram_read_data_2\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__18360\,
            I => \M_this_vram_read_data_2\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__18355\,
            I => \N__18350\
        );

    \I__2505\ : InMux
    port map (
            O => \N__18354\,
            I => \N__18343\
        );

    \I__2504\ : InMux
    port map (
            O => \N__18353\,
            I => \N__18343\
        );

    \I__2503\ : InMux
    port map (
            O => \N__18350\,
            I => \N__18335\
        );

    \I__2502\ : InMux
    port map (
            O => \N__18349\,
            I => \N__18335\
        );

    \I__2501\ : InMux
    port map (
            O => \N__18348\,
            I => \N__18335\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__18343\,
            I => \N__18332\
        );

    \I__2499\ : InMux
    port map (
            O => \N__18342\,
            I => \N__18329\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__18335\,
            I => \N__18326\
        );

    \I__2497\ : Span4Mux_h
    port map (
            O => \N__18332\,
            I => \N__18323\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__18329\,
            I => \N__18318\
        );

    \I__2495\ : Span4Mux_v
    port map (
            O => \N__18326\,
            I => \N__18318\
        );

    \I__2494\ : Span4Mux_v
    port map (
            O => \N__18323\,
            I => \N__18315\
        );

    \I__2493\ : Span4Mux_h
    port map (
            O => \N__18318\,
            I => \N__18312\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__18315\,
            I => \M_this_vram_read_data_3\
        );

    \I__2491\ : Odrv4
    port map (
            O => \N__18312\,
            I => \M_this_vram_read_data_3\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__18307\,
            I => \N__18304\
        );

    \I__2489\ : InMux
    port map (
            O => \N__18304\,
            I => \N__18295\
        );

    \I__2488\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18295\
        );

    \I__2487\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18287\
        );

    \I__2486\ : InMux
    port map (
            O => \N__18301\,
            I => \N__18287\
        );

    \I__2485\ : InMux
    port map (
            O => \N__18300\,
            I => \N__18287\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__18295\,
            I => \N__18284\
        );

    \I__2483\ : InMux
    port map (
            O => \N__18294\,
            I => \N__18281\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__18287\,
            I => \N__18278\
        );

    \I__2481\ : Span4Mux_h
    port map (
            O => \N__18284\,
            I => \N__18275\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__18281\,
            I => \N__18272\
        );

    \I__2479\ : Span12Mux_h
    port map (
            O => \N__18278\,
            I => \N__18269\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__18275\,
            I => \N__18266\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__18272\,
            I => \N__18263\
        );

    \I__2476\ : Odrv12
    port map (
            O => \N__18269\,
            I => \M_this_vram_read_data_1\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__18266\,
            I => \M_this_vram_read_data_1\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__18263\,
            I => \M_this_vram_read_data_1\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__18256\,
            I => \this_vga_ramdac.m6_cascade_\
        );

    \I__2472\ : InMux
    port map (
            O => \N__18253\,
            I => \N__18250\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__18250\,
            I => \N__18246\
        );

    \I__2470\ : InMux
    port map (
            O => \N__18249\,
            I => \N__18243\
        );

    \I__2469\ : Odrv4
    port map (
            O => \N__18246\,
            I => \this_vga_ramdac.N_3857_reto\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__18243\,
            I => \this_vga_ramdac.N_3857_reto\
        );

    \I__2467\ : InMux
    port map (
            O => \N__18238\,
            I => \N__18235\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__18235\,
            I => \N__18232\
        );

    \I__2465\ : Odrv12
    port map (
            O => \N__18232\,
            I => \this_ppu.oam_cache.mem_9\
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__18229\,
            I => \this_vga_signals.M_pcounter_q_ret_RNIB85CZ0Z3_cascade_\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__18226\,
            I => \this_vga_signals.N_3_0_cascade_\
        );

    \I__2462\ : InMux
    port map (
            O => \N__18223\,
            I => \N__18220\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__18220\,
            I => \N__18217\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__18217\,
            I => \this_vga_ramdac.m16\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__18214\,
            I => \M_pcounter_q_ret_1_RNIOILK7_cascade_\
        );

    \I__2458\ : InMux
    port map (
            O => \N__18211\,
            I => \N__18208\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__18208\,
            I => \N__18204\
        );

    \I__2456\ : InMux
    port map (
            O => \N__18207\,
            I => \N__18201\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__18204\,
            I => \this_vga_ramdac.N_3859_reto\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__18201\,
            I => \this_vga_ramdac.N_3859_reto\
        );

    \I__2453\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18193\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__18193\,
            I => \this_vga_signals.N_2_0\
        );

    \I__2451\ : InMux
    port map (
            O => \N__18190\,
            I => \N__18187\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__18187\,
            I => \N__18184\
        );

    \I__2449\ : Span4Mux_h
    port map (
            O => \N__18184\,
            I => \N__18181\
        );

    \I__2448\ : Odrv4
    port map (
            O => \N__18181\,
            I => \M_this_oam_ram_write_data_1\
        );

    \I__2447\ : InMux
    port map (
            O => \N__18178\,
            I => \N__18175\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__18175\,
            I => \N__18172\
        );

    \I__2445\ : Odrv12
    port map (
            O => \N__18172\,
            I => \M_this_oam_ram_write_data_25\
        );

    \I__2444\ : InMux
    port map (
            O => \N__18169\,
            I => \N__18166\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__18166\,
            I => \M_this_data_tmp_qZ0Z_21\
        );

    \I__2442\ : InMux
    port map (
            O => \N__18163\,
            I => \N__18160\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__18160\,
            I => \N__18157\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__18157\,
            I => \M_this_data_tmp_qZ0Z_23\
        );

    \I__2439\ : InMux
    port map (
            O => \N__18154\,
            I => \N__18151\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__18151\,
            I => \M_this_data_tmp_qZ0Z_0\
        );

    \I__2437\ : InMux
    port map (
            O => \N__18148\,
            I => \N__18144\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__18147\,
            I => \N__18141\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__18144\,
            I => \N__18138\
        );

    \I__2434\ : InMux
    port map (
            O => \N__18141\,
            I => \N__18135\
        );

    \I__2433\ : Odrv12
    port map (
            O => \N__18138\,
            I => \this_vga_ramdac.N_3856_reto\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__18135\,
            I => \this_vga_ramdac.N_3856_reto\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__18130\,
            I => \this_vga_ramdac.i2_mux_cascade_\
        );

    \I__2430\ : InMux
    port map (
            O => \N__18127\,
            I => \N__18124\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__18124\,
            I => \N__18121\
        );

    \I__2428\ : Span4Mux_h
    port map (
            O => \N__18121\,
            I => \N__18117\
        );

    \I__2427\ : InMux
    port map (
            O => \N__18120\,
            I => \N__18114\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__18117\,
            I => \this_vga_ramdac.N_3858_reto\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__18114\,
            I => \this_vga_ramdac.N_3858_reto\
        );

    \I__2424\ : InMux
    port map (
            O => \N__18109\,
            I => \N__18106\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__18106\,
            I => \N__18101\
        );

    \I__2422\ : InMux
    port map (
            O => \N__18105\,
            I => \N__18098\
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__18104\,
            I => \N__18093\
        );

    \I__2420\ : Span4Mux_v
    port map (
            O => \N__18101\,
            I => \N__18088\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__18098\,
            I => \N__18085\
        );

    \I__2418\ : InMux
    port map (
            O => \N__18097\,
            I => \N__18080\
        );

    \I__2417\ : InMux
    port map (
            O => \N__18096\,
            I => \N__18080\
        );

    \I__2416\ : InMux
    port map (
            O => \N__18093\,
            I => \N__18075\
        );

    \I__2415\ : InMux
    port map (
            O => \N__18092\,
            I => \N__18075\
        );

    \I__2414\ : InMux
    port map (
            O => \N__18091\,
            I => \N__18072\
        );

    \I__2413\ : Odrv4
    port map (
            O => \N__18088\,
            I => \N_852_0\
        );

    \I__2412\ : Odrv4
    port map (
            O => \N__18085\,
            I => \N_852_0\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__18080\,
            I => \N_852_0\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__18075\,
            I => \N_852_0\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__18072\,
            I => \N_852_0\
        );

    \I__2408\ : CascadeMux
    port map (
            O => \N__18061\,
            I => \N__18058\
        );

    \I__2407\ : InMux
    port map (
            O => \N__18058\,
            I => \N__18054\
        );

    \I__2406\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18051\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__18054\,
            I => \N__18048\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__18051\,
            I => \this_vga_signals.mult1_un54_sum_c3\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__18048\,
            I => \this_vga_signals.mult1_un54_sum_c3\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__18043\,
            I => \N__18040\
        );

    \I__2401\ : InMux
    port map (
            O => \N__18040\,
            I => \N__18037\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__18037\,
            I => \N__18034\
        );

    \I__2399\ : Span4Mux_h
    port map (
            O => \N__18034\,
            I => \N__18031\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__18031\,
            I => \M_this_vga_signals_address_5\
        );

    \I__2397\ : InMux
    port map (
            O => \N__18028\,
            I => \N__18025\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__18025\,
            I => \N__18022\
        );

    \I__2395\ : Span4Mux_h
    port map (
            O => \N__18022\,
            I => \N__18019\
        );

    \I__2394\ : Odrv4
    port map (
            O => \N__18019\,
            I => \M_this_oam_ram_write_data_3\
        );

    \I__2393\ : InMux
    port map (
            O => \N__18016\,
            I => \N__18013\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__18013\,
            I => \M_this_data_tmp_qZ0Z_3\
        );

    \I__2391\ : InMux
    port map (
            O => \N__18010\,
            I => \N__18007\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__18007\,
            I => \N__18004\
        );

    \I__2389\ : Span4Mux_v
    port map (
            O => \N__18004\,
            I => \N__18001\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__18001\,
            I => \M_this_oam_ram_write_data_4\
        );

    \I__2387\ : InMux
    port map (
            O => \N__17998\,
            I => \N__17995\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__17995\,
            I => \M_this_data_tmp_qZ0Z_4\
        );

    \I__2385\ : InMux
    port map (
            O => \N__17992\,
            I => \N__17989\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__17989\,
            I => \N__17986\
        );

    \I__2383\ : Span4Mux_h
    port map (
            O => \N__17986\,
            I => \N__17983\
        );

    \I__2382\ : Odrv4
    port map (
            O => \N__17983\,
            I => \M_this_data_tmp_qZ0Z_5\
        );

    \I__2381\ : InMux
    port map (
            O => \N__17980\,
            I => \N__17977\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__17977\,
            I => \N__17974\
        );

    \I__2379\ : Odrv12
    port map (
            O => \N__17974\,
            I => \M_this_oam_ram_write_data_29\
        );

    \I__2378\ : InMux
    port map (
            O => \N__17971\,
            I => \N__17968\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__17968\,
            I => \N__17965\
        );

    \I__2376\ : Span4Mux_h
    port map (
            O => \N__17965\,
            I => \N__17962\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__17962\,
            I => \M_this_oam_ram_write_data_21\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__17959\,
            I => \this_vga_signals.mult1_un54_sum_c3_cascade_\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__17956\,
            I => \N__17953\
        );

    \I__2372\ : InMux
    port map (
            O => \N__17953\,
            I => \N__17949\
        );

    \I__2371\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17946\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__17949\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0_0\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__17946\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0_0\
        );

    \I__2368\ : InMux
    port map (
            O => \N__17941\,
            I => \N__17938\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__17938\,
            I => \N__17934\
        );

    \I__2366\ : InMux
    port map (
            O => \N__17937\,
            I => \N__17931\
        );

    \I__2365\ : Span4Mux_v
    port map (
            O => \N__17934\,
            I => \N__17924\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__17931\,
            I => \N__17924\
        );

    \I__2363\ : InMux
    port map (
            O => \N__17930\,
            I => \N__17921\
        );

    \I__2362\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17917\
        );

    \I__2361\ : Span4Mux_h
    port map (
            O => \N__17924\,
            I => \N__17909\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__17921\,
            I => \N__17909\
        );

    \I__2359\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17906\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__17917\,
            I => \N__17902\
        );

    \I__2357\ : InMux
    port map (
            O => \N__17916\,
            I => \N__17899\
        );

    \I__2356\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17894\
        );

    \I__2355\ : InMux
    port map (
            O => \N__17914\,
            I => \N__17894\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__17909\,
            I => \N__17889\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__17906\,
            I => \N__17889\
        );

    \I__2352\ : InMux
    port map (
            O => \N__17905\,
            I => \N__17886\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__17902\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__17899\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__17894\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__17889\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__17886\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2346\ : InMux
    port map (
            O => \N__17875\,
            I => \N__17871\
        );

    \I__2345\ : InMux
    port map (
            O => \N__17874\,
            I => \N__17867\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__17871\,
            I => \N__17864\
        );

    \I__2343\ : InMux
    port map (
            O => \N__17870\,
            I => \N__17861\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__17867\,
            I => \N__17857\
        );

    \I__2341\ : Span4Mux_h
    port map (
            O => \N__17864\,
            I => \N__17848\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__17861\,
            I => \N__17848\
        );

    \I__2339\ : InMux
    port map (
            O => \N__17860\,
            I => \N__17845\
        );

    \I__2338\ : Span12Mux_s11_h
    port map (
            O => \N__17857\,
            I => \N__17841\
        );

    \I__2337\ : InMux
    port map (
            O => \N__17856\,
            I => \N__17838\
        );

    \I__2336\ : InMux
    port map (
            O => \N__17855\,
            I => \N__17835\
        );

    \I__2335\ : InMux
    port map (
            O => \N__17854\,
            I => \N__17832\
        );

    \I__2334\ : InMux
    port map (
            O => \N__17853\,
            I => \N__17829\
        );

    \I__2333\ : Span4Mux_v
    port map (
            O => \N__17848\,
            I => \N__17824\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__17845\,
            I => \N__17824\
        );

    \I__2331\ : InMux
    port map (
            O => \N__17844\,
            I => \N__17821\
        );

    \I__2330\ : Odrv12
    port map (
            O => \N__17841\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__17838\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__17835\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__17832\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__17829\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__17824\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__17821\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2323\ : InMux
    port map (
            O => \N__17806\,
            I => \N__17802\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__17805\,
            I => \N__17799\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__17802\,
            I => \N__17796\
        );

    \I__2320\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17793\
        );

    \I__2319\ : Span4Mux_h
    port map (
            O => \N__17796\,
            I => \N__17788\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__17793\,
            I => \N__17788\
        );

    \I__2317\ : Span4Mux_h
    port map (
            O => \N__17788\,
            I => \N__17781\
        );

    \I__2316\ : InMux
    port map (
            O => \N__17787\,
            I => \N__17778\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__17786\,
            I => \N__17775\
        );

    \I__2314\ : InMux
    port map (
            O => \N__17785\,
            I => \N__17770\
        );

    \I__2313\ : CascadeMux
    port map (
            O => \N__17784\,
            I => \N__17766\
        );

    \I__2312\ : Span4Mux_v
    port map (
            O => \N__17781\,
            I => \N__17761\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__17778\,
            I => \N__17761\
        );

    \I__2310\ : InMux
    port map (
            O => \N__17775\,
            I => \N__17758\
        );

    \I__2309\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17755\
        );

    \I__2308\ : InMux
    port map (
            O => \N__17773\,
            I => \N__17752\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__17770\,
            I => \N__17749\
        );

    \I__2306\ : InMux
    port map (
            O => \N__17769\,
            I => \N__17744\
        );

    \I__2305\ : InMux
    port map (
            O => \N__17766\,
            I => \N__17744\
        );

    \I__2304\ : Span4Mux_v
    port map (
            O => \N__17761\,
            I => \N__17739\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__17758\,
            I => \N__17739\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__17755\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__17752\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__17749\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__17744\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__17739\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2297\ : InMux
    port map (
            O => \N__17728\,
            I => \N__17724\
        );

    \I__2296\ : InMux
    port map (
            O => \N__17727\,
            I => \N__17721\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__17724\,
            I => \this_vga_signals.N_968\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__17721\,
            I => \this_vga_signals.N_968\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__17716\,
            I => \N__17713\
        );

    \I__2292\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17703\
        );

    \I__2291\ : InMux
    port map (
            O => \N__17712\,
            I => \N__17694\
        );

    \I__2290\ : InMux
    port map (
            O => \N__17711\,
            I => \N__17694\
        );

    \I__2289\ : InMux
    port map (
            O => \N__17710\,
            I => \N__17694\
        );

    \I__2288\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17689\
        );

    \I__2287\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17689\
        );

    \I__2286\ : InMux
    port map (
            O => \N__17707\,
            I => \N__17686\
        );

    \I__2285\ : InMux
    port map (
            O => \N__17706\,
            I => \N__17683\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__17703\,
            I => \N__17680\
        );

    \I__2283\ : InMux
    port map (
            O => \N__17702\,
            I => \N__17675\
        );

    \I__2282\ : InMux
    port map (
            O => \N__17701\,
            I => \N__17675\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__17694\,
            I => \N__17670\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__17689\,
            I => \N__17670\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__17686\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__17683\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__17680\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__17675\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__17670\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__17659\,
            I => \this_vga_signals.N_968_cascade_\
        );

    \I__2273\ : InMux
    port map (
            O => \N__17656\,
            I => \N__17650\
        );

    \I__2272\ : InMux
    port map (
            O => \N__17655\,
            I => \N__17650\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__17650\,
            I => \N__17646\
        );

    \I__2270\ : InMux
    port map (
            O => \N__17649\,
            I => \N__17643\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__17646\,
            I => \this_vga_signals.N_291_0\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__17643\,
            I => \this_vga_signals.N_291_0\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__17638\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_\
        );

    \I__2266\ : InMux
    port map (
            O => \N__17635\,
            I => \N__17629\
        );

    \I__2265\ : InMux
    port map (
            O => \N__17634\,
            I => \N__17629\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__17629\,
            I => \this_vga_signals.mult1_un68_sum_axb1\
        );

    \I__2263\ : InMux
    port map (
            O => \N__17626\,
            I => \N__17623\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__17623\,
            I => \this_vga_signals.mult1_un68_sum_ac0_2\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__17620\,
            I => \this_vga_signals.mult1_un68_sum_axb1_cascade_\
        );

    \I__2260\ : InMux
    port map (
            O => \N__17617\,
            I => \N__17613\
        );

    \I__2259\ : InMux
    port map (
            O => \N__17616\,
            I => \N__17610\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__17613\,
            I => \this_vga_signals.mult1_un68_sum_axb2\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__17610\,
            I => \this_vga_signals.mult1_un68_sum_axb2\
        );

    \I__2256\ : InMux
    port map (
            O => \N__17605\,
            I => \N__17601\
        );

    \I__2255\ : InMux
    port map (
            O => \N__17604\,
            I => \N__17598\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__17601\,
            I => \N__17595\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__17598\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__17595\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0\
        );

    \I__2251\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17587\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__17587\,
            I => \N__17584\
        );

    \I__2249\ : Span4Mux_h
    port map (
            O => \N__17584\,
            I => \N__17580\
        );

    \I__2248\ : InMux
    port map (
            O => \N__17583\,
            I => \N__17577\
        );

    \I__2247\ : Span4Mux_v
    port map (
            O => \N__17580\,
            I => \N__17572\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__17577\,
            I => \N__17572\
        );

    \I__2245\ : Span4Mux_h
    port map (
            O => \N__17572\,
            I => \N__17569\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__17569\,
            I => \M_this_oam_ram_read_data_20\
        );

    \I__2243\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17563\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__17563\,
            I => \N__17560\
        );

    \I__2241\ : Span4Mux_v
    port map (
            O => \N__17560\,
            I => \N__17557\
        );

    \I__2240\ : Span4Mux_h
    port map (
            O => \N__17557\,
            I => \N__17554\
        );

    \I__2239\ : Odrv4
    port map (
            O => \N__17554\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_20\
        );

    \I__2238\ : InMux
    port map (
            O => \N__17551\,
            I => \N__17548\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__17548\,
            I => \N__17545\
        );

    \I__2236\ : Span4Mux_v
    port map (
            O => \N__17545\,
            I => \N__17542\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__17542\,
            I => \this_ppu.oam_cache.mem_13\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__17539\,
            I => \N__17536\
        );

    \I__2233\ : InMux
    port map (
            O => \N__17536\,
            I => \N__17533\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__17533\,
            I => \N__17530\
        );

    \I__2231\ : Odrv12
    port map (
            O => \N__17530\,
            I => \M_this_vga_signals_address_4\
        );

    \I__2230\ : InMux
    port map (
            O => \N__17527\,
            I => \bfn_12_18_0_\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__17524\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_3_1_0_cascade_\
        );

    \I__2228\ : InMux
    port map (
            O => \N__17521\,
            I => \N__17518\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__17518\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0_0_tz\
        );

    \I__2226\ : InMux
    port map (
            O => \N__17515\,
            I => \N__17512\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__17512\,
            I => \N__17509\
        );

    \I__2224\ : Span4Mux_h
    port map (
            O => \N__17509\,
            I => \N__17505\
        );

    \I__2223\ : InMux
    port map (
            O => \N__17508\,
            I => \N__17502\
        );

    \I__2222\ : Odrv4
    port map (
            O => \N__17505\,
            I => \this_ppu.N_1184_7\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__17502\,
            I => \this_ppu.N_1184_7\
        );

    \I__2220\ : InMux
    port map (
            O => \N__17497\,
            I => \N__17494\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__17494\,
            I => \N__17491\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__17491\,
            I => \this_ppu.un1_M_state_q_7_i_0\
        );

    \I__2217\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17485\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__17485\,
            I => \N__17482\
        );

    \I__2215\ : Span12Mux_v
    port map (
            O => \N__17482\,
            I => \N__17479\
        );

    \I__2214\ : Odrv12
    port map (
            O => \N__17479\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__2213\ : InMux
    port map (
            O => \N__17476\,
            I => \N__17473\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__17473\,
            I => \N__17470\
        );

    \I__2211\ : Span4Mux_h
    port map (
            O => \N__17470\,
            I => \N__17467\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__17467\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_11\
        );

    \I__2209\ : InMux
    port map (
            O => \N__17464\,
            I => \N__17461\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__17461\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_12\
        );

    \I__2207\ : InMux
    port map (
            O => \N__17458\,
            I => \N__17455\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__17455\,
            I => \N__17452\
        );

    \I__2205\ : Span4Mux_h
    port map (
            O => \N__17452\,
            I => \N__17449\
        );

    \I__2204\ : Span4Mux_h
    port map (
            O => \N__17449\,
            I => \N__17446\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__17446\,
            I => \this_ppu.oam_cache.mem_15\
        );

    \I__2202\ : InMux
    port map (
            O => \N__17443\,
            I => \N__17439\
        );

    \I__2201\ : InMux
    port map (
            O => \N__17442\,
            I => \N__17436\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__17439\,
            I => \this_vga_signals.N_298_0\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__17436\,
            I => \this_vga_signals.N_298_0\
        );

    \I__2198\ : InMux
    port map (
            O => \N__17431\,
            I => \N__17428\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__17428\,
            I => \this_vga_signals.hsync_1_i_0_0_a3_0\
        );

    \I__2196\ : InMux
    port map (
            O => \N__17425\,
            I => \N__17422\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__17422\,
            I => \N__17419\
        );

    \I__2194\ : Span4Mux_h
    port map (
            O => \N__17419\,
            I => \N__17413\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__17418\,
            I => \N__17410\
        );

    \I__2192\ : InMux
    port map (
            O => \N__17417\,
            I => \N__17405\
        );

    \I__2191\ : InMux
    port map (
            O => \N__17416\,
            I => \N__17402\
        );

    \I__2190\ : Span4Mux_v
    port map (
            O => \N__17413\,
            I => \N__17399\
        );

    \I__2189\ : InMux
    port map (
            O => \N__17410\,
            I => \N__17392\
        );

    \I__2188\ : InMux
    port map (
            O => \N__17409\,
            I => \N__17392\
        );

    \I__2187\ : InMux
    port map (
            O => \N__17408\,
            I => \N__17392\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__17405\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__17402\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__17399\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__17392\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2182\ : InMux
    port map (
            O => \N__17383\,
            I => \N__17380\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__17380\,
            I => \N__17375\
        );

    \I__2180\ : InMux
    port map (
            O => \N__17379\,
            I => \N__17372\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__17378\,
            I => \N__17369\
        );

    \I__2178\ : Span4Mux_h
    port map (
            O => \N__17375\,
            I => \N__17365\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__17372\,
            I => \N__17362\
        );

    \I__2176\ : InMux
    port map (
            O => \N__17369\,
            I => \N__17359\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__17368\,
            I => \N__17355\
        );

    \I__2174\ : Span4Mux_h
    port map (
            O => \N__17365\,
            I => \N__17348\
        );

    \I__2173\ : Span4Mux_h
    port map (
            O => \N__17362\,
            I => \N__17348\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__17359\,
            I => \N__17348\
        );

    \I__2171\ : InMux
    port map (
            O => \N__17358\,
            I => \N__17342\
        );

    \I__2170\ : InMux
    port map (
            O => \N__17355\,
            I => \N__17339\
        );

    \I__2169\ : Span4Mux_v
    port map (
            O => \N__17348\,
            I => \N__17336\
        );

    \I__2168\ : InMux
    port map (
            O => \N__17347\,
            I => \N__17329\
        );

    \I__2167\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17329\
        );

    \I__2166\ : InMux
    port map (
            O => \N__17345\,
            I => \N__17329\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__17342\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__17339\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__17336\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__17329\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2161\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17314\
        );

    \I__2160\ : InMux
    port map (
            O => \N__17319\,
            I => \N__17307\
        );

    \I__2159\ : InMux
    port map (
            O => \N__17318\,
            I => \N__17307\
        );

    \I__2158\ : InMux
    port map (
            O => \N__17317\,
            I => \N__17307\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__17314\,
            I => \N__17299\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__17307\,
            I => \N__17299\
        );

    \I__2155\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17294\
        );

    \I__2154\ : InMux
    port map (
            O => \N__17305\,
            I => \N__17294\
        );

    \I__2153\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17291\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__17299\,
            I => \N__17288\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__17294\,
            I => \N__17285\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__17291\,
            I => \N__17277\
        );

    \I__2149\ : Span4Mux_h
    port map (
            O => \N__17288\,
            I => \N__17277\
        );

    \I__2148\ : Span4Mux_v
    port map (
            O => \N__17285\,
            I => \N__17277\
        );

    \I__2147\ : InMux
    port map (
            O => \N__17284\,
            I => \N__17274\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__17277\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__17274\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2144\ : InMux
    port map (
            O => \N__17269\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__2143\ : InMux
    port map (
            O => \N__17266\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__2142\ : InMux
    port map (
            O => \N__17263\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__2141\ : InMux
    port map (
            O => \N__17260\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__2140\ : InMux
    port map (
            O => \N__17257\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__2139\ : InMux
    port map (
            O => \N__17254\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__2138\ : InMux
    port map (
            O => \N__17251\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__2137\ : InMux
    port map (
            O => \N__17248\,
            I => \N__17245\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__17245\,
            I => \N__17242\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__17242\,
            I => \M_this_data_tmp_qZ0Z_20\
        );

    \I__2134\ : InMux
    port map (
            O => \N__17239\,
            I => \N__17236\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__17236\,
            I => \N__17233\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__17233\,
            I => \M_this_data_tmp_qZ0Z_18\
        );

    \I__2131\ : InMux
    port map (
            O => \N__17230\,
            I => \N__17227\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__17227\,
            I => \N__17224\
        );

    \I__2129\ : Span4Mux_h
    port map (
            O => \N__17224\,
            I => \N__17221\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__17221\,
            I => \M_this_oam_ram_write_data_0\
        );

    \I__2127\ : InMux
    port map (
            O => \N__17218\,
            I => \N__17213\
        );

    \I__2126\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17208\
        );

    \I__2125\ : InMux
    port map (
            O => \N__17216\,
            I => \N__17208\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__17213\,
            I => \N__17201\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__17208\,
            I => \N__17201\
        );

    \I__2122\ : InMux
    port map (
            O => \N__17207\,
            I => \N__17198\
        );

    \I__2121\ : InMux
    port map (
            O => \N__17206\,
            I => \N__17195\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__17201\,
            I => \N__17190\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__17198\,
            I => \N__17187\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__17195\,
            I => \N__17184\
        );

    \I__2117\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17181\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__17193\,
            I => \N__17178\
        );

    \I__2115\ : Span4Mux_h
    port map (
            O => \N__17190\,
            I => \N__17171\
        );

    \I__2114\ : Span4Mux_v
    port map (
            O => \N__17187\,
            I => \N__17171\
        );

    \I__2113\ : Span4Mux_v
    port map (
            O => \N__17184\,
            I => \N__17171\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__17181\,
            I => \N__17168\
        );

    \I__2111\ : InMux
    port map (
            O => \N__17178\,
            I => \N__17165\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__17171\,
            I => \this_vga_ramdac.N_852_i_reto\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__17168\,
            I => \this_vga_ramdac.N_852_i_reto\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__17165\,
            I => \this_vga_ramdac.N_852_i_reto\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__17158\,
            I => \this_vga_signals.N_298_0_cascade_\
        );

    \I__2106\ : InMux
    port map (
            O => \N__17155\,
            I => \N__17152\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__17152\,
            I => \N__17149\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__17149\,
            I => \this_vga_signals.M_hcounter_d7_0_i_0_o3_0_o3_4_a2_0\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__17146\,
            I => \this_vga_signals.N_1044_0_cascade_\
        );

    \I__2102\ : InMux
    port map (
            O => \N__17143\,
            I => \N__17140\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__17140\,
            I => \M_this_data_tmp_qZ0Z_8\
        );

    \I__2100\ : InMux
    port map (
            O => \N__17137\,
            I => \N__17134\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__17134\,
            I => \M_this_data_tmp_qZ0Z_9\
        );

    \I__2098\ : InMux
    port map (
            O => \N__17131\,
            I => \N__17128\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__17128\,
            I => \N__17125\
        );

    \I__2096\ : Odrv12
    port map (
            O => \N__17125\,
            I => \M_this_oam_ram_write_data_26\
        );

    \I__2095\ : InMux
    port map (
            O => \N__17122\,
            I => \N__17119\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__17119\,
            I => \N__17116\
        );

    \I__2093\ : Odrv4
    port map (
            O => \N__17116\,
            I => \M_this_oam_ram_write_data_27\
        );

    \I__2092\ : InMux
    port map (
            O => \N__17113\,
            I => \N__17110\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__17110\,
            I => \N__17107\
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__17107\,
            I => \M_this_oam_ram_write_data_30\
        );

    \I__2089\ : InMux
    port map (
            O => \N__17104\,
            I => \N__17101\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__17101\,
            I => \M_this_data_tmp_qZ0Z_15\
        );

    \I__2087\ : InMux
    port map (
            O => \N__17098\,
            I => \N__17095\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__17095\,
            I => \N__17092\
        );

    \I__2085\ : Span4Mux_h
    port map (
            O => \N__17092\,
            I => \N__17089\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__17089\,
            I => \M_this_oam_ram_write_data_15\
        );

    \I__2083\ : InMux
    port map (
            O => \N__17086\,
            I => \N__17083\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__17083\,
            I => \M_this_data_tmp_qZ0Z_16\
        );

    \I__2081\ : InMux
    port map (
            O => \N__17080\,
            I => \N__17077\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__17077\,
            I => \N__17074\
        );

    \I__2079\ : Span4Mux_h
    port map (
            O => \N__17074\,
            I => \N__17071\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__17071\,
            I => \M_this_data_tmp_qZ0Z_17\
        );

    \I__2077\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17065\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__17065\,
            I => \N__17062\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__17062\,
            I => \M_this_data_tmp_qZ0Z_19\
        );

    \I__2074\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17056\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__17056\,
            I => \N__17053\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__17053\,
            I => \this_ppu.un1_oam_data_1_axb_7\
        );

    \I__2071\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17047\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__17047\,
            I => \N__17044\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__17044\,
            I => \N__17041\
        );

    \I__2068\ : Span4Mux_h
    port map (
            O => \N__17041\,
            I => \N__17038\
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__17038\,
            I => \M_this_oam_ram_write_data_6\
        );

    \I__2066\ : InMux
    port map (
            O => \N__17035\,
            I => \N__17032\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__17032\,
            I => \M_this_data_tmp_qZ0Z_6\
        );

    \I__2064\ : InMux
    port map (
            O => \N__17029\,
            I => \N__17026\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__17026\,
            I => \N__17023\
        );

    \I__2062\ : Span4Mux_h
    port map (
            O => \N__17023\,
            I => \N__17020\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__17020\,
            I => \M_this_oam_ram_write_data_7\
        );

    \I__2060\ : InMux
    port map (
            O => \N__17017\,
            I => \N__17014\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__17014\,
            I => \M_this_data_tmp_qZ0Z_7\
        );

    \I__2058\ : InMux
    port map (
            O => \N__17011\,
            I => \N__17007\
        );

    \I__2057\ : InMux
    port map (
            O => \N__17010\,
            I => \N__17004\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__17007\,
            I => \N__17001\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__17004\,
            I => \N__16998\
        );

    \I__2054\ : Span4Mux_h
    port map (
            O => \N__17001\,
            I => \N__16995\
        );

    \I__2053\ : Span12Mux_v
    port map (
            O => \N__16998\,
            I => \N__16992\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__16995\,
            I => \M_this_oam_ram_read_data_17\
        );

    \I__2051\ : Odrv12
    port map (
            O => \N__16992\,
            I => \M_this_oam_ram_read_data_17\
        );

    \I__2050\ : InMux
    port map (
            O => \N__16987\,
            I => \N__16984\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__16984\,
            I => \N__16981\
        );

    \I__2048\ : Span12Mux_v
    port map (
            O => \N__16981\,
            I => \N__16978\
        );

    \I__2047\ : Odrv12
    port map (
            O => \N__16978\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_17\
        );

    \I__2046\ : InMux
    port map (
            O => \N__16975\,
            I => \N__16972\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__16972\,
            I => \M_this_data_tmp_qZ0Z_10\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__16969\,
            I => \this_vga_signals.mult1_un68_sum_ac0_2_cascade_\
        );

    \I__2043\ : InMux
    port map (
            O => \N__16966\,
            I => \N__16963\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__16963\,
            I => \this_vga_signals.mult1_un68_sum_c3_1\
        );

    \I__2041\ : InMux
    port map (
            O => \N__16960\,
            I => \N__16952\
        );

    \I__2040\ : InMux
    port map (
            O => \N__16959\,
            I => \N__16947\
        );

    \I__2039\ : InMux
    port map (
            O => \N__16958\,
            I => \N__16947\
        );

    \I__2038\ : InMux
    port map (
            O => \N__16957\,
            I => \N__16942\
        );

    \I__2037\ : InMux
    port map (
            O => \N__16956\,
            I => \N__16942\
        );

    \I__2036\ : InMux
    port map (
            O => \N__16955\,
            I => \N__16939\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__16952\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__16947\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__16942\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__16939\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__2031\ : InMux
    port map (
            O => \N__16930\,
            I => \N__16927\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__16927\,
            I => \this_vga_signals.mult1_un75_sum_c2_0\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__16924\,
            I => \this_vga_signals.mult1_un75_sum_c2_0_cascade_\
        );

    \I__2028\ : InMux
    port map (
            O => \N__16921\,
            I => \N__16918\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__16918\,
            I => \this_vga_signals.if_N_8_i\
        );

    \I__2026\ : InMux
    port map (
            O => \N__16915\,
            I => \N__16912\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__16912\,
            I => \N__16909\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__16909\,
            I => \N__16906\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__16906\,
            I => \this_delay_clk.M_pipe_qZ0Z_2\
        );

    \I__2022\ : InMux
    port map (
            O => \N__16903\,
            I => \N__16900\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__16900\,
            I => \N__16897\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__16897\,
            I => \N__16894\
        );

    \I__2019\ : Span4Mux_h
    port map (
            O => \N__16894\,
            I => \N__16891\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__16891\,
            I => \M_this_oam_ram_read_data_27\
        );

    \I__2017\ : InMux
    port map (
            O => \N__16888\,
            I => \N__16885\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__16885\,
            I => \N__16882\
        );

    \I__2015\ : Span4Mux_h
    port map (
            O => \N__16882\,
            I => \N__16879\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__16879\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_27\
        );

    \I__2013\ : InMux
    port map (
            O => \N__16876\,
            I => \N__16873\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__16873\,
            I => \N__16870\
        );

    \I__2011\ : Span4Mux_v
    port map (
            O => \N__16870\,
            I => \N__16867\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__16867\,
            I => \this_ppu.oam_cache.mem_0\
        );

    \I__2009\ : InMux
    port map (
            O => \N__16864\,
            I => \N__16861\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__16861\,
            I => \N__16857\
        );

    \I__2007\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16854\
        );

    \I__2006\ : Span4Mux_h
    port map (
            O => \N__16857\,
            I => \N__16851\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__16854\,
            I => \N__16848\
        );

    \I__2004\ : Span4Mux_v
    port map (
            O => \N__16851\,
            I => \N__16845\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__16848\,
            I => \M_this_oam_ram_read_data_2\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__16845\,
            I => \M_this_oam_ram_read_data_2\
        );

    \I__2001\ : InMux
    port map (
            O => \N__16840\,
            I => \N__16837\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__16837\,
            I => \N__16834\
        );

    \I__1999\ : Span4Mux_h
    port map (
            O => \N__16834\,
            I => \N__16831\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__16831\,
            I => \this_ppu.m28_e_i_a3_4\
        );

    \I__1997\ : InMux
    port map (
            O => \N__16828\,
            I => \N__16825\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__16825\,
            I => \this_ppu.m28_e_i_a3_3\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__16822\,
            I => \this_ppu.N_1184_7_cascade_\
        );

    \I__1994\ : InMux
    port map (
            O => \N__16819\,
            I => \N__16816\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__16816\,
            I => \this_ppu.m18_i_1\
        );

    \I__1992\ : InMux
    port map (
            O => \N__16813\,
            I => \N__16810\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__16810\,
            I => \N__16806\
        );

    \I__1990\ : InMux
    port map (
            O => \N__16809\,
            I => \N__16803\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__16806\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0_2\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__16803\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0_2\
        );

    \I__1987\ : InMux
    port map (
            O => \N__16798\,
            I => \N__16795\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__16795\,
            I => \N__16792\
        );

    \I__1985\ : Span4Mux_v
    port map (
            O => \N__16792\,
            I => \N__16789\
        );

    \I__1984\ : Odrv4
    port map (
            O => \N__16789\,
            I => \this_ppu.oam_cache.mem_12\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__16786\,
            I => \N__16782\
        );

    \I__1982\ : InMux
    port map (
            O => \N__16785\,
            I => \N__16777\
        );

    \I__1981\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16777\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__16777\,
            I => \N__16774\
        );

    \I__1979\ : Span4Mux_h
    port map (
            O => \N__16774\,
            I => \N__16771\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__16771\,
            I => \N__16768\
        );

    \I__1977\ : Odrv4
    port map (
            O => \N__16768\,
            I => \M_this_oam_ram_read_data_5\
        );

    \I__1976\ : InMux
    port map (
            O => \N__16765\,
            I => \N__16762\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__16762\,
            I => \N__16759\
        );

    \I__1974\ : Span4Mux_h
    port map (
            O => \N__16759\,
            I => \N__16756\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__16756\,
            I => \this_ppu.oam_cache.N_569_0\
        );

    \I__1972\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16749\
        );

    \I__1971\ : InMux
    port map (
            O => \N__16752\,
            I => \N__16746\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__16749\,
            I => \N__16741\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__16746\,
            I => \N__16741\
        );

    \I__1968\ : Span4Mux_h
    port map (
            O => \N__16741\,
            I => \N__16738\
        );

    \I__1967\ : Span4Mux_v
    port map (
            O => \N__16738\,
            I => \N__16735\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__16735\,
            I => \M_this_oam_ram_read_data_4\
        );

    \I__1965\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16729\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__16729\,
            I => \N__16726\
        );

    \I__1963\ : Span4Mux_h
    port map (
            O => \N__16726\,
            I => \N__16723\
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__16723\,
            I => \this_ppu.oam_cache.N_575_0\
        );

    \I__1961\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16717\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__16717\,
            I => \this_ppu.N_1182\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__16714\,
            I => \this_vga_signals.if_N_9_0_0_cascade_\
        );

    \I__1958\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16708\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__16708\,
            I => \this_vga_signals.mult1_un82_sum_c3\
        );

    \I__1956\ : InMux
    port map (
            O => \N__16705\,
            I => \N__16702\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__16702\,
            I => \this_vga_signals.N_811_0\
        );

    \I__1954\ : IoInMux
    port map (
            O => \N__16699\,
            I => \N__16696\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__16696\,
            I => \N__16693\
        );

    \I__1952\ : Span4Mux_s3_h
    port map (
            O => \N__16693\,
            I => \N__16690\
        );

    \I__1951\ : Span4Mux_v
    port map (
            O => \N__16690\,
            I => \N__16687\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__16687\,
            I => \N__16684\
        );

    \I__1949\ : Span4Mux_h
    port map (
            O => \N__16684\,
            I => \N__16681\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__16681\,
            I => rgb_c_3
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__16678\,
            I => \N__16675\
        );

    \I__1946\ : CascadeBuf
    port map (
            O => \N__16675\,
            I => \N__16672\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__16672\,
            I => \N__16669\
        );

    \I__1944\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16666\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__16666\,
            I => \N__16663\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__16663\,
            I => \N__16657\
        );

    \I__1941\ : InMux
    port map (
            O => \N__16662\,
            I => \N__16652\
        );

    \I__1940\ : InMux
    port map (
            O => \N__16661\,
            I => \N__16652\
        );

    \I__1939\ : InMux
    port map (
            O => \N__16660\,
            I => \N__16649\
        );

    \I__1938\ : Span4Mux_v
    port map (
            O => \N__16657\,
            I => \N__16646\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__16652\,
            I => \M_this_ppu_oam_addr_5\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__16649\,
            I => \M_this_ppu_oam_addr_5\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__16646\,
            I => \M_this_ppu_oam_addr_5\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__16639\,
            I => \N__16636\
        );

    \I__1933\ : CascadeBuf
    port map (
            O => \N__16636\,
            I => \N__16633\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__16633\,
            I => \N__16628\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__16632\,
            I => \N__16625\
        );

    \I__1930\ : InMux
    port map (
            O => \N__16631\,
            I => \N__16620\
        );

    \I__1929\ : InMux
    port map (
            O => \N__16628\,
            I => \N__16617\
        );

    \I__1928\ : InMux
    port map (
            O => \N__16625\,
            I => \N__16610\
        );

    \I__1927\ : InMux
    port map (
            O => \N__16624\,
            I => \N__16610\
        );

    \I__1926\ : InMux
    port map (
            O => \N__16623\,
            I => \N__16610\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__16620\,
            I => \N__16604\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__16617\,
            I => \N__16601\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__16610\,
            I => \N__16598\
        );

    \I__1922\ : InMux
    port map (
            O => \N__16609\,
            I => \N__16593\
        );

    \I__1921\ : InMux
    port map (
            O => \N__16608\,
            I => \N__16593\
        );

    \I__1920\ : InMux
    port map (
            O => \N__16607\,
            I => \N__16590\
        );

    \I__1919\ : Span4Mux_h
    port map (
            O => \N__16604\,
            I => \N__16585\
        );

    \I__1918\ : Span4Mux_v
    port map (
            O => \N__16601\,
            I => \N__16585\
        );

    \I__1917\ : Odrv4
    port map (
            O => \N__16598\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__16593\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__16590\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__16585\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__1913\ : InMux
    port map (
            O => \N__16576\,
            I => \N__16573\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__16573\,
            I => \N__16570\
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__16570\,
            I => \this_ppu.m35_i_0_a3_1_3\
        );

    \I__1910\ : InMux
    port map (
            O => \N__16567\,
            I => \N__16563\
        );

    \I__1909\ : InMux
    port map (
            O => \N__16566\,
            I => \N__16560\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__16563\,
            I => \N__16557\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__16560\,
            I => \N__16554\
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__16557\,
            I => \this_ppu.N_1394\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__16554\,
            I => \this_ppu.N_1394\
        );

    \I__1904\ : InMux
    port map (
            O => \N__16549\,
            I => \N__16546\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__16546\,
            I => \N__16543\
        );

    \I__1902\ : Span4Mux_h
    port map (
            O => \N__16543\,
            I => \N__16540\
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__16540\,
            I => \M_this_oam_ram_write_data_9\
        );

    \I__1900\ : InMux
    port map (
            O => \N__16537\,
            I => \N__16534\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__16534\,
            I => \N__16531\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__16531\,
            I => \M_this_oam_ram_read_data_i_20\
        );

    \I__1897\ : InMux
    port map (
            O => \N__16528\,
            I => \N__16525\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__16525\,
            I => \N__16522\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__16522\,
            I => \M_this_oam_ram_write_data_28\
        );

    \I__1894\ : InMux
    port map (
            O => \N__16519\,
            I => \N__16516\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__16516\,
            I => \N__16513\
        );

    \I__1892\ : Span4Mux_h
    port map (
            O => \N__16513\,
            I => \N__16510\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__16510\,
            I => \M_this_oam_ram_write_data_8\
        );

    \I__1890\ : InMux
    port map (
            O => \N__16507\,
            I => \N__16504\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__16504\,
            I => \N__16501\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__16501\,
            I => \M_this_oam_ram_write_data_31\
        );

    \I__1887\ : InMux
    port map (
            O => \N__16498\,
            I => \N__16495\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__16495\,
            I => \N__16492\
        );

    \I__1885\ : Odrv4
    port map (
            O => \N__16492\,
            I => \M_this_oam_ram_write_data_16\
        );

    \I__1884\ : InMux
    port map (
            O => \N__16489\,
            I => \N__16486\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__16486\,
            I => \N__16483\
        );

    \I__1882\ : Span4Mux_h
    port map (
            O => \N__16483\,
            I => \N__16480\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__16480\,
            I => \M_this_oam_ram_write_data_24\
        );

    \I__1880\ : InMux
    port map (
            O => \N__16477\,
            I => \N__16474\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__16474\,
            I => \N__16471\
        );

    \I__1878\ : Sp12to4
    port map (
            O => \N__16471\,
            I => \N__16468\
        );

    \I__1877\ : Odrv12
    port map (
            O => \N__16468\,
            I => \this_vga_signals.hsync_1_i_0_0_1\
        );

    \I__1876\ : InMux
    port map (
            O => \N__16465\,
            I => \N__16462\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__16462\,
            I => \N__16459\
        );

    \I__1874\ : Span4Mux_h
    port map (
            O => \N__16459\,
            I => \N__16456\
        );

    \I__1873\ : Span4Mux_v
    port map (
            O => \N__16456\,
            I => \N__16453\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__16453\,
            I => \M_this_oam_ram_read_data_14\
        );

    \I__1871\ : InMux
    port map (
            O => \N__16450\,
            I => \N__16447\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__16447\,
            I => \N__16444\
        );

    \I__1869\ : Span4Mux_h
    port map (
            O => \N__16444\,
            I => \N__16441\
        );

    \I__1868\ : Odrv4
    port map (
            O => \N__16441\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_14\
        );

    \I__1867\ : InMux
    port map (
            O => \N__16438\,
            I => \N__16435\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__16435\,
            I => \this_vga_signals.hsync_1_i_0_0_a3_0_0\
        );

    \I__1865\ : InMux
    port map (
            O => \N__16432\,
            I => \N__16429\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__16429\,
            I => \N__16426\
        );

    \I__1863\ : Span12Mux_h
    port map (
            O => \N__16426\,
            I => \N__16423\
        );

    \I__1862\ : Odrv12
    port map (
            O => \N__16423\,
            I => \M_this_oam_ram_read_data_29\
        );

    \I__1861\ : InMux
    port map (
            O => \N__16420\,
            I => \N__16417\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__16417\,
            I => \N__16414\
        );

    \I__1859\ : Span4Mux_h
    port map (
            O => \N__16414\,
            I => \N__16411\
        );

    \I__1858\ : Odrv4
    port map (
            O => \N__16411\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_29\
        );

    \I__1857\ : InMux
    port map (
            O => \N__16408\,
            I => \N__16404\
        );

    \I__1856\ : InMux
    port map (
            O => \N__16407\,
            I => \N__16401\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__16404\,
            I => \N__16398\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__16401\,
            I => \N__16395\
        );

    \I__1853\ : Span4Mux_v
    port map (
            O => \N__16398\,
            I => \N__16392\
        );

    \I__1852\ : Span4Mux_h
    port map (
            O => \N__16395\,
            I => \N__16389\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__16392\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__16389\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__16384\,
            I => \N__16381\
        );

    \I__1848\ : InMux
    port map (
            O => \N__16381\,
            I => \N__16378\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__16378\,
            I => \M_this_oam_ram_read_data_i_21\
        );

    \I__1846\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16372\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__16372\,
            I => \N__16369\
        );

    \I__1844\ : Span4Mux_h
    port map (
            O => \N__16369\,
            I => \N__16366\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__16366\,
            I => \M_this_oam_ram_read_data_31\
        );

    \I__1842\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16360\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__16360\,
            I => \N__16357\
        );

    \I__1840\ : Span4Mux_h
    port map (
            O => \N__16357\,
            I => \N__16354\
        );

    \I__1839\ : Odrv4
    port map (
            O => \N__16354\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_31\
        );

    \I__1838\ : InMux
    port map (
            O => \N__16351\,
            I => \N__16348\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__16348\,
            I => \N__16345\
        );

    \I__1836\ : Span4Mux_h
    port map (
            O => \N__16345\,
            I => \N__16342\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__16342\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_19\
        );

    \I__1834\ : InMux
    port map (
            O => \N__16339\,
            I => \N__16333\
        );

    \I__1833\ : InMux
    port map (
            O => \N__16338\,
            I => \N__16333\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__16333\,
            I => \N__16330\
        );

    \I__1831\ : Span4Mux_v
    port map (
            O => \N__16330\,
            I => \N__16327\
        );

    \I__1830\ : Odrv4
    port map (
            O => \N__16327\,
            I => \M_this_oam_ram_read_data_19\
        );

    \I__1829\ : InMux
    port map (
            O => \N__16324\,
            I => \N__16321\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__16321\,
            I => \M_this_oam_ram_read_data_i_19\
        );

    \I__1827\ : InMux
    port map (
            O => \N__16318\,
            I => \N__16315\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__16315\,
            I => \N__16312\
        );

    \I__1825\ : Span4Mux_h
    port map (
            O => \N__16312\,
            I => \N__16309\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__16309\,
            I => \M_this_oam_ram_write_data_10\
        );

    \I__1823\ : IoInMux
    port map (
            O => \N__16306\,
            I => \N__16303\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__16303\,
            I => \N__16300\
        );

    \I__1821\ : Span12Mux_s8_v
    port map (
            O => \N__16300\,
            I => \N__16297\
        );

    \I__1820\ : Odrv12
    port map (
            O => \N__16297\,
            I => \N_260\
        );

    \I__1819\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16291\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__16291\,
            I => \N__16288\
        );

    \I__1817\ : Span4Mux_h
    port map (
            O => \N__16288\,
            I => \N__16285\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__16285\,
            I => \M_this_oam_ram_read_data_28\
        );

    \I__1815\ : InMux
    port map (
            O => \N__16282\,
            I => \N__16279\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__16279\,
            I => \N__16276\
        );

    \I__1813\ : Span12Mux_v
    port map (
            O => \N__16276\,
            I => \N__16273\
        );

    \I__1812\ : Odrv12
    port map (
            O => \N__16273\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_28\
        );

    \I__1811\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16267\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__16267\,
            I => \this_ppu.M_this_oam_ram_read_data_i_18\
        );

    \I__1809\ : InMux
    port map (
            O => \N__16264\,
            I => \this_ppu.un1_oam_data_1_cry_2\
        );

    \I__1808\ : InMux
    port map (
            O => \N__16261\,
            I => \this_ppu.un1_oam_data_1_cry_3\
        );

    \I__1807\ : InMux
    port map (
            O => \N__16258\,
            I => \N__16255\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__16255\,
            I => \N__16251\
        );

    \I__1805\ : InMux
    port map (
            O => \N__16254\,
            I => \N__16248\
        );

    \I__1804\ : Odrv12
    port map (
            O => \N__16251\,
            I => \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__16248\,
            I => \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0\
        );

    \I__1802\ : InMux
    port map (
            O => \N__16243\,
            I => \this_ppu.un1_oam_data_1_cry_4\
        );

    \I__1801\ : InMux
    port map (
            O => \N__16240\,
            I => \N__16237\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__16237\,
            I => \N__16234\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__16234\,
            I => \N__16230\
        );

    \I__1798\ : InMux
    port map (
            O => \N__16233\,
            I => \N__16227\
        );

    \I__1797\ : Odrv4
    port map (
            O => \N__16230\,
            I => \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__16227\,
            I => \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0\
        );

    \I__1795\ : InMux
    port map (
            O => \N__16222\,
            I => \this_ppu.un1_oam_data_1_cry_5\
        );

    \I__1794\ : InMux
    port map (
            O => \N__16219\,
            I => \N__16216\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__16216\,
            I => \this_ppu.un1_oam_data_1_cry_3_c_RNIT7IDZ0\
        );

    \I__1792\ : CascadeMux
    port map (
            O => \N__16213\,
            I => \N__16210\
        );

    \I__1791\ : InMux
    port map (
            O => \N__16210\,
            I => \N__16207\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__16207\,
            I => \this_ppu.un1_oam_data_1_cry_2_c_RNIR4HDZ0\
        );

    \I__1789\ : InMux
    port map (
            O => \N__16204\,
            I => \this_ppu.un1_oam_data_1_cry_6\
        );

    \I__1788\ : InMux
    port map (
            O => \N__16201\,
            I => \N__16198\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__16198\,
            I => \N__16195\
        );

    \I__1786\ : Span4Mux_v
    port map (
            O => \N__16195\,
            I => \N__16191\
        );

    \I__1785\ : InMux
    port map (
            O => \N__16194\,
            I => \N__16188\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__16191\,
            I => \this_ppu.m28_e_i_o3_2\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__16188\,
            I => \this_ppu.m28_e_i_o3_2\
        );

    \I__1782\ : InMux
    port map (
            O => \N__16183\,
            I => \N__16179\
        );

    \I__1781\ : InMux
    port map (
            O => \N__16182\,
            I => \N__16176\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__16179\,
            I => \N__16173\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__16176\,
            I => \N__16170\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__16173\,
            I => \N__16167\
        );

    \I__1777\ : Span4Mux_h
    port map (
            O => \N__16170\,
            I => \N__16164\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__16167\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__16164\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__1774\ : InMux
    port map (
            O => \N__16159\,
            I => \N__16156\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__16156\,
            I => \N__16153\
        );

    \I__1772\ : Span4Mux_h
    port map (
            O => \N__16153\,
            I => \N__16150\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__16150\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_18\
        );

    \I__1770\ : InMux
    port map (
            O => \N__16147\,
            I => \N__16144\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__16144\,
            I => \N__16141\
        );

    \I__1768\ : Span4Mux_h
    port map (
            O => \N__16141\,
            I => \N__16138\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__16138\,
            I => \M_this_oam_ram_write_data_5\
        );

    \I__1766\ : InMux
    port map (
            O => \N__16135\,
            I => \N__16131\
        );

    \I__1765\ : InMux
    port map (
            O => \N__16134\,
            I => \N__16128\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__16131\,
            I => \N__16125\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__16128\,
            I => \N__16122\
        );

    \I__1762\ : Span4Mux_v
    port map (
            O => \N__16125\,
            I => \N__16119\
        );

    \I__1761\ : Span4Mux_h
    port map (
            O => \N__16122\,
            I => \N__16116\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__16119\,
            I => \M_this_oam_ram_read_data_22\
        );

    \I__1759\ : Odrv4
    port map (
            O => \N__16116\,
            I => \M_this_oam_ram_read_data_22\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__16111\,
            I => \N__16108\
        );

    \I__1757\ : InMux
    port map (
            O => \N__16108\,
            I => \N__16105\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__16105\,
            I => \M_this_oam_ram_read_data_i_22\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__16102\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_cascade_\
        );

    \I__1754\ : InMux
    port map (
            O => \N__16099\,
            I => \N__16093\
        );

    \I__1753\ : InMux
    port map (
            O => \N__16098\,
            I => \N__16093\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__16093\,
            I => \this_vga_signals.if_m2\
        );

    \I__1751\ : InMux
    port map (
            O => \N__16090\,
            I => \N__16086\
        );

    \I__1750\ : InMux
    port map (
            O => \N__16089\,
            I => \N__16083\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__16086\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__16083\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__16078\,
            I => \N__16075\
        );

    \I__1746\ : InMux
    port map (
            O => \N__16075\,
            I => \N__16072\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__16072\,
            I => \N__16069\
        );

    \I__1744\ : Odrv12
    port map (
            O => \N__16069\,
            I => \M_this_vga_signals_address_1\
        );

    \I__1743\ : InMux
    port map (
            O => \N__16066\,
            I => \N__16063\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__16063\,
            I => \this_vga_signals.mult1_un75_sum_axb1\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__16060\,
            I => \N__16057\
        );

    \I__1740\ : CascadeBuf
    port map (
            O => \N__16057\,
            I => \N__16054\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__16054\,
            I => \N__16050\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__16053\,
            I => \N__16045\
        );

    \I__1737\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16042\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__16049\,
            I => \N__16039\
        );

    \I__1735\ : InMux
    port map (
            O => \N__16048\,
            I => \N__16036\
        );

    \I__1734\ : InMux
    port map (
            O => \N__16045\,
            I => \N__16033\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__16042\,
            I => \N__16030\
        );

    \I__1732\ : InMux
    port map (
            O => \N__16039\,
            I => \N__16027\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__16036\,
            I => \N__16022\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__16033\,
            I => \N__16022\
        );

    \I__1729\ : Span4Mux_h
    port map (
            O => \N__16030\,
            I => \N__16019\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__16027\,
            I => \this_ppu.M_oam_cache_cnt_qZ1Z_0\
        );

    \I__1727\ : Odrv12
    port map (
            O => \N__16022\,
            I => \this_ppu.M_oam_cache_cnt_qZ1Z_0\
        );

    \I__1726\ : Odrv4
    port map (
            O => \N__16019\,
            I => \this_ppu.M_oam_cache_cnt_qZ1Z_0\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__16012\,
            I => \N__16009\
        );

    \I__1724\ : InMux
    port map (
            O => \N__16009\,
            I => \N__16006\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__16006\,
            I => \N__16003\
        );

    \I__1722\ : Odrv4
    port map (
            O => \N__16003\,
            I => \M_this_vga_signals_address_3\
        );

    \I__1721\ : InMux
    port map (
            O => \N__16000\,
            I => \N__15996\
        );

    \I__1720\ : InMux
    port map (
            O => \N__15999\,
            I => \N__15993\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__15996\,
            I => \N__15990\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__15993\,
            I => \N__15987\
        );

    \I__1717\ : Span4Mux_h
    port map (
            O => \N__15990\,
            I => \N__15984\
        );

    \I__1716\ : Span12Mux_v
    port map (
            O => \N__15987\,
            I => \N__15981\
        );

    \I__1715\ : Span4Mux_v
    port map (
            O => \N__15984\,
            I => \N__15978\
        );

    \I__1714\ : Odrv12
    port map (
            O => \N__15981\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__1713\ : Odrv4
    port map (
            O => \N__15978\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__1712\ : InMux
    port map (
            O => \N__15973\,
            I => \N__15970\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__15970\,
            I => \this_ppu.M_this_oam_ram_read_data_i_16\
        );

    \I__1710\ : InMux
    port map (
            O => \N__15967\,
            I => \N__15964\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__15964\,
            I => \this_ppu.M_this_oam_ram_read_data_i_17\
        );

    \I__1708\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15958\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__15958\,
            I => \N__15955\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__15955\,
            I => \N__15952\
        );

    \I__1705\ : Span4Mux_v
    port map (
            O => \N__15952\,
            I => \N__15949\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__15949\,
            I => \M_this_oam_ram_read_data_24\
        );

    \I__1703\ : InMux
    port map (
            O => \N__15946\,
            I => \N__15943\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__15943\,
            I => \N__15940\
        );

    \I__1701\ : Odrv4
    port map (
            O => \N__15940\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_24\
        );

    \I__1700\ : InMux
    port map (
            O => \N__15937\,
            I => \N__15934\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__15934\,
            I => \N__15931\
        );

    \I__1698\ : Span4Mux_h
    port map (
            O => \N__15931\,
            I => \N__15928\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__15928\,
            I => \this_delay_clk.M_pipe_qZ0Z_1\
        );

    \I__1696\ : InMux
    port map (
            O => \N__15925\,
            I => \N__15921\
        );

    \I__1695\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15918\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__15921\,
            I => \N__15915\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__15918\,
            I => \N__15912\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__15915\,
            I => \N__15909\
        );

    \I__1691\ : Span4Mux_v
    port map (
            O => \N__15912\,
            I => \N__15906\
        );

    \I__1690\ : Span4Mux_v
    port map (
            O => \N__15909\,
            I => \N__15903\
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__15906\,
            I => \M_this_oam_ram_read_data_7\
        );

    \I__1688\ : Odrv4
    port map (
            O => \N__15903\,
            I => \M_this_oam_ram_read_data_7\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__15898\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__15895\,
            I => \this_vga_signals.mult1_un82_sum_axb1_cascade_\
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__15892\,
            I => \this_vga_signals.mult1_un89_sum_c3_cascade_\
        );

    \I__1684\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15886\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__15886\,
            I => \this_vga_signals.haddress_1_0\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__15883\,
            I => \N__15880\
        );

    \I__1681\ : InMux
    port map (
            O => \N__15880\,
            I => \N__15877\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__15877\,
            I => \N__15874\
        );

    \I__1679\ : Span4Mux_v
    port map (
            O => \N__15874\,
            I => \N__15871\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__15871\,
            I => \M_this_vga_signals_address_0\
        );

    \I__1677\ : InMux
    port map (
            O => \N__15868\,
            I => \N__15862\
        );

    \I__1676\ : InMux
    port map (
            O => \N__15867\,
            I => \N__15862\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__15862\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0_0\
        );

    \I__1674\ : InMux
    port map (
            O => \N__15859\,
            I => \N__15856\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__15856\,
            I => \this_ppu.un1_M_oam_curr_q_1_c4\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__15853\,
            I => \N__15848\
        );

    \I__1671\ : InMux
    port map (
            O => \N__15852\,
            I => \N__15836\
        );

    \I__1670\ : InMux
    port map (
            O => \N__15851\,
            I => \N__15836\
        );

    \I__1669\ : InMux
    port map (
            O => \N__15848\,
            I => \N__15836\
        );

    \I__1668\ : InMux
    port map (
            O => \N__15847\,
            I => \N__15836\
        );

    \I__1667\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15830\
        );

    \I__1666\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15830\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__15836\,
            I => \N__15827\
        );

    \I__1664\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15824\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__15830\,
            I => \this_ppu.M_oam_curr_qc_0_1\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__15827\,
            I => \this_ppu.M_oam_curr_qc_0_1\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__15824\,
            I => \this_ppu.M_oam_curr_qc_0_1\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__15817\,
            I => \N__15814\
        );

    \I__1659\ : InMux
    port map (
            O => \N__15814\,
            I => \N__15811\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__15811\,
            I => \N__15808\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__15808\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_CO\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__15805\,
            I => \N__15802\
        );

    \I__1655\ : CascadeBuf
    port map (
            O => \N__15802\,
            I => \N__15799\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__15799\,
            I => \N__15796\
        );

    \I__1653\ : InMux
    port map (
            O => \N__15796\,
            I => \N__15791\
        );

    \I__1652\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15787\
        );

    \I__1651\ : InMux
    port map (
            O => \N__15794\,
            I => \N__15784\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__15791\,
            I => \N__15781\
        );

    \I__1649\ : InMux
    port map (
            O => \N__15790\,
            I => \N__15778\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__15787\,
            I => \N__15775\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__15784\,
            I => \N__15770\
        );

    \I__1646\ : Span4Mux_h
    port map (
            O => \N__15781\,
            I => \N__15770\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__15778\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_1\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__15775\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_1\
        );

    \I__1643\ : Odrv4
    port map (
            O => \N__15770\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_1\
        );

    \I__1642\ : InMux
    port map (
            O => \N__15763\,
            I => \N__15760\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__15760\,
            I => \this_ppu.m62_0_a2_0_o2_1\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__15757\,
            I => \N__15754\
        );

    \I__1639\ : CascadeBuf
    port map (
            O => \N__15754\,
            I => \N__15751\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__15751\,
            I => \N__15748\
        );

    \I__1637\ : InMux
    port map (
            O => \N__15748\,
            I => \N__15743\
        );

    \I__1636\ : InMux
    port map (
            O => \N__15747\,
            I => \N__15738\
        );

    \I__1635\ : InMux
    port map (
            O => \N__15746\,
            I => \N__15738\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__15743\,
            I => \N__15734\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__15738\,
            I => \N__15729\
        );

    \I__1632\ : InMux
    port map (
            O => \N__15737\,
            I => \N__15725\
        );

    \I__1631\ : Span4Mux_h
    port map (
            O => \N__15734\,
            I => \N__15722\
        );

    \I__1630\ : InMux
    port map (
            O => \N__15733\,
            I => \N__15719\
        );

    \I__1629\ : InMux
    port map (
            O => \N__15732\,
            I => \N__15716\
        );

    \I__1628\ : Span4Mux_h
    port map (
            O => \N__15729\,
            I => \N__15713\
        );

    \I__1627\ : InMux
    port map (
            O => \N__15728\,
            I => \N__15710\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__15725\,
            I => \N__15705\
        );

    \I__1625\ : Span4Mux_v
    port map (
            O => \N__15722\,
            I => \N__15705\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__15719\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__15716\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__15713\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__15710\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__1620\ : Odrv4
    port map (
            O => \N__15705\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__15694\,
            I => \N__15691\
        );

    \I__1618\ : CascadeBuf
    port map (
            O => \N__15691\,
            I => \N__15688\
        );

    \I__1617\ : CascadeMux
    port map (
            O => \N__15688\,
            I => \N__15685\
        );

    \I__1616\ : InMux
    port map (
            O => \N__15685\,
            I => \N__15682\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__15682\,
            I => \N__15679\
        );

    \I__1614\ : Span4Mux_h
    port map (
            O => \N__15679\,
            I => \N__15668\
        );

    \I__1613\ : InMux
    port map (
            O => \N__15678\,
            I => \N__15665\
        );

    \I__1612\ : InMux
    port map (
            O => \N__15677\,
            I => \N__15662\
        );

    \I__1611\ : InMux
    port map (
            O => \N__15676\,
            I => \N__15657\
        );

    \I__1610\ : InMux
    port map (
            O => \N__15675\,
            I => \N__15657\
        );

    \I__1609\ : InMux
    port map (
            O => \N__15674\,
            I => \N__15650\
        );

    \I__1608\ : InMux
    port map (
            O => \N__15673\,
            I => \N__15650\
        );

    \I__1607\ : InMux
    port map (
            O => \N__15672\,
            I => \N__15650\
        );

    \I__1606\ : InMux
    port map (
            O => \N__15671\,
            I => \N__15647\
        );

    \I__1605\ : Span4Mux_v
    port map (
            O => \N__15668\,
            I => \N__15644\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__15665\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__15662\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__15657\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__15650\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__15647\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__1599\ : Odrv4
    port map (
            O => \N__15644\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__15631\,
            I => \N__15628\
        );

    \I__1597\ : CascadeBuf
    port map (
            O => \N__15628\,
            I => \N__15625\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__15625\,
            I => \N__15622\
        );

    \I__1595\ : InMux
    port map (
            O => \N__15622\,
            I => \N__15616\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__15621\,
            I => \N__15612\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__15620\,
            I => \N__15609\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__15619\,
            I => \N__15605\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__15616\,
            I => \N__15602\
        );

    \I__1590\ : InMux
    port map (
            O => \N__15615\,
            I => \N__15599\
        );

    \I__1589\ : InMux
    port map (
            O => \N__15612\,
            I => \N__15596\
        );

    \I__1588\ : InMux
    port map (
            O => \N__15609\,
            I => \N__15591\
        );

    \I__1587\ : InMux
    port map (
            O => \N__15608\,
            I => \N__15591\
        );

    \I__1586\ : InMux
    port map (
            O => \N__15605\,
            I => \N__15588\
        );

    \I__1585\ : Span4Mux_v
    port map (
            O => \N__15602\,
            I => \N__15585\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__15599\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__15596\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__15591\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__15588\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__15585\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__1579\ : InMux
    port map (
            O => \N__15574\,
            I => \N__15565\
        );

    \I__1578\ : InMux
    port map (
            O => \N__15573\,
            I => \N__15565\
        );

    \I__1577\ : InMux
    port map (
            O => \N__15572\,
            I => \N__15562\
        );

    \I__1576\ : InMux
    port map (
            O => \N__15571\,
            I => \N__15557\
        );

    \I__1575\ : InMux
    port map (
            O => \N__15570\,
            I => \N__15557\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__15565\,
            I => \this_ppu.un1_M_oam_curr_q_1_c2\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__15562\,
            I => \this_ppu.un1_M_oam_curr_q_1_c2\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__15557\,
            I => \this_ppu.un1_M_oam_curr_q_1_c2\
        );

    \I__1571\ : InMux
    port map (
            O => \N__15550\,
            I => \N__15547\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__15547\,
            I => \this_ppu.un1_M_oam_curr_q_1_c5\
        );

    \I__1569\ : InMux
    port map (
            O => \N__15544\,
            I => \N__15541\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__15541\,
            I => \N__15538\
        );

    \I__1567\ : Odrv12
    port map (
            O => \N__15538\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_CO\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__15535\,
            I => \N__15532\
        );

    \I__1565\ : CascadeBuf
    port map (
            O => \N__15532\,
            I => \N__15529\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__15529\,
            I => \N__15524\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__15528\,
            I => \N__15520\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__15527\,
            I => \N__15517\
        );

    \I__1561\ : InMux
    port map (
            O => \N__15524\,
            I => \N__15514\
        );

    \I__1560\ : InMux
    port map (
            O => \N__15523\,
            I => \N__15511\
        );

    \I__1559\ : InMux
    port map (
            O => \N__15520\,
            I => \N__15506\
        );

    \I__1558\ : InMux
    port map (
            O => \N__15517\,
            I => \N__15506\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__15514\,
            I => \N__15503\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__15511\,
            I => \N__15500\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__15506\,
            I => \N__15495\
        );

    \I__1554\ : Span4Mux_v
    port map (
            O => \N__15503\,
            I => \N__15495\
        );

    \I__1553\ : Odrv12
    port map (
            O => \N__15500\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_3\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__15495\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_3\
        );

    \I__1551\ : InMux
    port map (
            O => \N__15490\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_0\
        );

    \I__1550\ : InMux
    port map (
            O => \N__15487\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_1\
        );

    \I__1549\ : InMux
    port map (
            O => \N__15484\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_2\
        );

    \I__1548\ : InMux
    port map (
            O => \N__15481\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_3\
        );

    \I__1547\ : InMux
    port map (
            O => \N__15478\,
            I => \N__15475\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__15475\,
            I => \N__15472\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__15472\,
            I => \N__15469\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__15469\,
            I => \this_ppu.oam_cache.mem_7\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__15466\,
            I => \N__15463\
        );

    \I__1542\ : InMux
    port map (
            O => \N__15463\,
            I => \N__15460\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__15460\,
            I => \N__15457\
        );

    \I__1540\ : Span4Mux_v
    port map (
            O => \N__15457\,
            I => \N__15454\
        );

    \I__1539\ : Odrv4
    port map (
            O => \N__15454\,
            I => \N_41_0\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__15451\,
            I => \N__15448\
        );

    \I__1537\ : CascadeBuf
    port map (
            O => \N__15448\,
            I => \N__15445\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__15445\,
            I => \N__15442\
        );

    \I__1535\ : InMux
    port map (
            O => \N__15442\,
            I => \N__15436\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__15441\,
            I => \N__15432\
        );

    \I__1533\ : InMux
    port map (
            O => \N__15440\,
            I => \N__15428\
        );

    \I__1532\ : InMux
    port map (
            O => \N__15439\,
            I => \N__15425\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__15436\,
            I => \N__15422\
        );

    \I__1530\ : InMux
    port map (
            O => \N__15435\,
            I => \N__15419\
        );

    \I__1529\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15414\
        );

    \I__1528\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15414\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__15428\,
            I => \N__15411\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__15425\,
            I => \N__15408\
        );

    \I__1525\ : Span4Mux_v
    port map (
            O => \N__15422\,
            I => \N__15405\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__15419\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__15414\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__1522\ : Odrv4
    port map (
            O => \N__15411\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__1521\ : Odrv4
    port map (
            O => \N__15408\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__15405\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__1519\ : InMux
    port map (
            O => \N__15394\,
            I => \N__15390\
        );

    \I__1518\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15387\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__15390\,
            I => \N__15384\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__15387\,
            I => \N__15381\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__15384\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_4\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__15381\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_4\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__15376\,
            I => \this_ppu.m62_0_a2_0_o2_0_cascade_\
        );

    \I__1512\ : InMux
    port map (
            O => \N__15373\,
            I => \N__15370\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__15370\,
            I => \M_this_oam_ram_write_data_23\
        );

    \I__1510\ : InMux
    port map (
            O => \N__15367\,
            I => \N__15364\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__15364\,
            I => \M_this_oam_ram_write_data_20\
        );

    \I__1508\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15358\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__15358\,
            I => \M_this_oam_ram_write_data_19\
        );

    \I__1506\ : InMux
    port map (
            O => \N__15355\,
            I => \N__15352\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__15352\,
            I => \M_this_oam_ram_write_data_17\
        );

    \I__1504\ : IoInMux
    port map (
            O => \N__15349\,
            I => \N__15346\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__15346\,
            I => \N__15343\
        );

    \I__1502\ : IoSpan4Mux
    port map (
            O => \N__15343\,
            I => \N__15340\
        );

    \I__1501\ : Span4Mux_s3_h
    port map (
            O => \N__15340\,
            I => \N__15337\
        );

    \I__1500\ : Span4Mux_h
    port map (
            O => \N__15337\,
            I => \N__15334\
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__15334\,
            I => rgb_c_1
        );

    \I__1498\ : InMux
    port map (
            O => \N__15331\,
            I => \N__15328\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__15328\,
            I => \N__15325\
        );

    \I__1496\ : Span4Mux_h
    port map (
            O => \N__15325\,
            I => \N__15321\
        );

    \I__1495\ : InMux
    port map (
            O => \N__15324\,
            I => \N__15318\
        );

    \I__1494\ : Span4Mux_v
    port map (
            O => \N__15321\,
            I => \N__15315\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__15318\,
            I => \N__15312\
        );

    \I__1492\ : Span4Mux_v
    port map (
            O => \N__15315\,
            I => \N__15309\
        );

    \I__1491\ : Span4Mux_h
    port map (
            O => \N__15312\,
            I => \N__15306\
        );

    \I__1490\ : Odrv4
    port map (
            O => \N__15309\,
            I => \M_this_oam_ram_read_data_0\
        );

    \I__1489\ : Odrv4
    port map (
            O => \N__15306\,
            I => \M_this_oam_ram_read_data_0\
        );

    \I__1488\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15298\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__15298\,
            I => \N__15295\
        );

    \I__1486\ : Span4Mux_h
    port map (
            O => \N__15295\,
            I => \N__15292\
        );

    \I__1485\ : Odrv4
    port map (
            O => \N__15292\,
            I => \this_ppu.oam_cache.N_586_0\
        );

    \I__1484\ : InMux
    port map (
            O => \N__15289\,
            I => \N__15286\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__15286\,
            I => \N__15283\
        );

    \I__1482\ : Span4Mux_h
    port map (
            O => \N__15283\,
            I => \N__15280\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__15280\,
            I => \this_ppu.oam_cache.mem_10\
        );

    \I__1480\ : InMux
    port map (
            O => \N__15277\,
            I => \N__15274\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__15274\,
            I => \this_ppu.N_844_0\
        );

    \I__1478\ : InMux
    port map (
            O => \N__15271\,
            I => \N__15268\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__15268\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_10\
        );

    \I__1476\ : InMux
    port map (
            O => \N__15265\,
            I => \un1_M_this_warmup_d_cry_20\
        );

    \I__1475\ : InMux
    port map (
            O => \N__15262\,
            I => \N__15259\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__15259\,
            I => \M_this_warmup_qZ0Z_22\
        );

    \I__1473\ : InMux
    port map (
            O => \N__15256\,
            I => \un1_M_this_warmup_d_cry_21\
        );

    \I__1472\ : InMux
    port map (
            O => \N__15253\,
            I => \N__15250\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__15250\,
            I => \M_this_warmup_qZ0Z_23\
        );

    \I__1470\ : InMux
    port map (
            O => \N__15247\,
            I => \un1_M_this_warmup_d_cry_22\
        );

    \I__1469\ : InMux
    port map (
            O => \N__15244\,
            I => \N__15241\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__15241\,
            I => \M_this_warmup_qZ0Z_24\
        );

    \I__1467\ : InMux
    port map (
            O => \N__15238\,
            I => \un1_M_this_warmup_d_cry_23\
        );

    \I__1466\ : InMux
    port map (
            O => \N__15235\,
            I => \N__15232\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__15232\,
            I => \M_this_warmup_qZ0Z_25\
        );

    \I__1464\ : InMux
    port map (
            O => \N__15229\,
            I => \bfn_9_25_0_\
        );

    \I__1463\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15223\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__15223\,
            I => \M_this_warmup_qZ0Z_26\
        );

    \I__1461\ : InMux
    port map (
            O => \N__15220\,
            I => \un1_M_this_warmup_d_cry_25\
        );

    \I__1460\ : InMux
    port map (
            O => \N__15217\,
            I => \un1_M_this_warmup_d_cry_26\
        );

    \I__1459\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15208\
        );

    \I__1458\ : InMux
    port map (
            O => \N__15213\,
            I => \N__15208\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__15208\,
            I => \M_this_warmup_qZ0Z_27\
        );

    \I__1456\ : InMux
    port map (
            O => \N__15205\,
            I => \N__15202\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__15202\,
            I => \M_this_oam_ram_write_data_18\
        );

    \I__1454\ : InMux
    port map (
            O => \N__15199\,
            I => \N__15196\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__15196\,
            I => \M_this_warmup_qZ0Z_13\
        );

    \I__1452\ : InMux
    port map (
            O => \N__15193\,
            I => \un1_M_this_warmup_d_cry_12\
        );

    \I__1451\ : InMux
    port map (
            O => \N__15190\,
            I => \N__15187\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__15187\,
            I => \M_this_warmup_qZ0Z_14\
        );

    \I__1449\ : InMux
    port map (
            O => \N__15184\,
            I => \un1_M_this_warmup_d_cry_13\
        );

    \I__1448\ : InMux
    port map (
            O => \N__15181\,
            I => \N__15178\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__15178\,
            I => \M_this_warmup_qZ0Z_15\
        );

    \I__1446\ : InMux
    port map (
            O => \N__15175\,
            I => \un1_M_this_warmup_d_cry_14\
        );

    \I__1445\ : InMux
    port map (
            O => \N__15172\,
            I => \N__15169\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__15169\,
            I => \M_this_warmup_qZ0Z_16\
        );

    \I__1443\ : InMux
    port map (
            O => \N__15166\,
            I => \un1_M_this_warmup_d_cry_15\
        );

    \I__1442\ : InMux
    port map (
            O => \N__15163\,
            I => \N__15160\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__15160\,
            I => \M_this_warmup_qZ0Z_17\
        );

    \I__1440\ : InMux
    port map (
            O => \N__15157\,
            I => \bfn_9_24_0_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__15154\,
            I => \N__15151\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__15151\,
            I => \M_this_warmup_qZ0Z_18\
        );

    \I__1437\ : InMux
    port map (
            O => \N__15148\,
            I => \un1_M_this_warmup_d_cry_17\
        );

    \I__1436\ : InMux
    port map (
            O => \N__15145\,
            I => \N__15142\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__15142\,
            I => \M_this_warmup_qZ0Z_19\
        );

    \I__1434\ : InMux
    port map (
            O => \N__15139\,
            I => \un1_M_this_warmup_d_cry_18\
        );

    \I__1433\ : InMux
    port map (
            O => \N__15136\,
            I => \N__15133\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__15133\,
            I => \M_this_warmup_qZ0Z_20\
        );

    \I__1431\ : InMux
    port map (
            O => \N__15130\,
            I => \un1_M_this_warmup_d_cry_19\
        );

    \I__1430\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15124\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__15124\,
            I => \M_this_warmup_qZ0Z_21\
        );

    \I__1428\ : InMux
    port map (
            O => \N__15121\,
            I => \N__15118\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__15118\,
            I => \M_this_warmup_qZ0Z_5\
        );

    \I__1426\ : InMux
    port map (
            O => \N__15115\,
            I => \un1_M_this_warmup_d_cry_4\
        );

    \I__1425\ : InMux
    port map (
            O => \N__15112\,
            I => \N__15109\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__15109\,
            I => \M_this_warmup_qZ0Z_6\
        );

    \I__1423\ : InMux
    port map (
            O => \N__15106\,
            I => \un1_M_this_warmup_d_cry_5\
        );

    \I__1422\ : InMux
    port map (
            O => \N__15103\,
            I => \N__15100\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__15100\,
            I => \M_this_warmup_qZ0Z_7\
        );

    \I__1420\ : InMux
    port map (
            O => \N__15097\,
            I => \un1_M_this_warmup_d_cry_6\
        );

    \I__1419\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15091\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__15091\,
            I => \M_this_warmup_qZ0Z_8\
        );

    \I__1417\ : InMux
    port map (
            O => \N__15088\,
            I => \un1_M_this_warmup_d_cry_7\
        );

    \I__1416\ : InMux
    port map (
            O => \N__15085\,
            I => \N__15082\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__15082\,
            I => \M_this_warmup_qZ0Z_9\
        );

    \I__1414\ : InMux
    port map (
            O => \N__15079\,
            I => \bfn_9_23_0_\
        );

    \I__1413\ : InMux
    port map (
            O => \N__15076\,
            I => \N__15073\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__15073\,
            I => \M_this_warmup_qZ0Z_10\
        );

    \I__1411\ : InMux
    port map (
            O => \N__15070\,
            I => \un1_M_this_warmup_d_cry_9\
        );

    \I__1410\ : InMux
    port map (
            O => \N__15067\,
            I => \N__15064\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__15064\,
            I => \M_this_warmup_qZ0Z_11\
        );

    \I__1408\ : InMux
    port map (
            O => \N__15061\,
            I => \un1_M_this_warmup_d_cry_10\
        );

    \I__1407\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15055\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__15055\,
            I => \M_this_warmup_qZ0Z_12\
        );

    \I__1405\ : InMux
    port map (
            O => \N__15052\,
            I => \un1_M_this_warmup_d_cry_11\
        );

    \I__1404\ : InMux
    port map (
            O => \N__15049\,
            I => \N__15046\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__15046\,
            I => \N__15043\
        );

    \I__1402\ : Span4Mux_h
    port map (
            O => \N__15043\,
            I => \N__15040\
        );

    \I__1401\ : Odrv4
    port map (
            O => \N__15040\,
            I => \this_ppu.oam_cache.mem_2\
        );

    \I__1400\ : InMux
    port map (
            O => \N__15037\,
            I => \N__15034\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__15034\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_21\
        );

    \I__1398\ : InMux
    port map (
            O => \N__15031\,
            I => \N__15028\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__15028\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_22\
        );

    \I__1396\ : InMux
    port map (
            O => \N__15025\,
            I => \N__15022\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__15022\,
            I => \N__15018\
        );

    \I__1394\ : InMux
    port map (
            O => \N__15021\,
            I => \N__15015\
        );

    \I__1393\ : Span4Mux_v
    port map (
            O => \N__15018\,
            I => \N__15010\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__15015\,
            I => \N__15010\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__15010\,
            I => \M_this_oam_ram_read_data_3\
        );

    \I__1390\ : InMux
    port map (
            O => \N__15007\,
            I => \N__15003\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__15006\,
            I => \N__15000\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__15003\,
            I => \N__14997\
        );

    \I__1387\ : InMux
    port map (
            O => \N__15000\,
            I => \N__14994\
        );

    \I__1386\ : Span4Mux_v
    port map (
            O => \N__14997\,
            I => \N__14989\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__14994\,
            I => \N__14989\
        );

    \I__1384\ : Odrv4
    port map (
            O => \N__14989\,
            I => \M_this_oam_ram_read_data_6\
        );

    \I__1383\ : InMux
    port map (
            O => \N__14986\,
            I => \N__14983\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__14983\,
            I => \N__14980\
        );

    \I__1381\ : Span4Mux_v
    port map (
            O => \N__14980\,
            I => \N__14977\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__14977\,
            I => \M_this_oam_ram_read_data_25\
        );

    \I__1379\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14971\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__14971\,
            I => \N__14968\
        );

    \I__1377\ : Span4Mux_h
    port map (
            O => \N__14968\,
            I => \N__14965\
        );

    \I__1376\ : Odrv4
    port map (
            O => \N__14965\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_25\
        );

    \I__1375\ : InMux
    port map (
            O => \N__14962\,
            I => \N__14958\
        );

    \I__1374\ : InMux
    port map (
            O => \N__14961\,
            I => \N__14955\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__14958\,
            I => \N__14952\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__14955\,
            I => \M_this_warmup_qZ0Z_1\
        );

    \I__1371\ : Odrv4
    port map (
            O => \N__14952\,
            I => \M_this_warmup_qZ0Z_1\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__14947\,
            I => \N__14942\
        );

    \I__1369\ : InMux
    port map (
            O => \N__14946\,
            I => \N__14937\
        );

    \I__1368\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14937\
        );

    \I__1367\ : InMux
    port map (
            O => \N__14942\,
            I => \N__14934\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__14937\,
            I => \N__14929\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__14934\,
            I => \N__14929\
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__14929\,
            I => \M_this_warmup_qZ0Z_0\
        );

    \I__1363\ : InMux
    port map (
            O => \N__14926\,
            I => \N__14923\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__14923\,
            I => \M_this_warmup_qZ0Z_2\
        );

    \I__1361\ : InMux
    port map (
            O => \N__14920\,
            I => \un1_M_this_warmup_d_cry_1\
        );

    \I__1360\ : InMux
    port map (
            O => \N__14917\,
            I => \N__14914\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__14914\,
            I => \M_this_warmup_qZ0Z_3\
        );

    \I__1358\ : InMux
    port map (
            O => \N__14911\,
            I => \un1_M_this_warmup_d_cry_2\
        );

    \I__1357\ : InMux
    port map (
            O => \N__14908\,
            I => \N__14905\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__14905\,
            I => \M_this_warmup_qZ0Z_4\
        );

    \I__1355\ : InMux
    port map (
            O => \N__14902\,
            I => \un1_M_this_warmup_d_cry_3\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__14899\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_cascade_\
        );

    \I__1353\ : InMux
    port map (
            O => \N__14896\,
            I => \N__14891\
        );

    \I__1352\ : InMux
    port map (
            O => \N__14895\,
            I => \N__14886\
        );

    \I__1351\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14886\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__14891\,
            I => \N__14883\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__14886\,
            I => \this_ppu.N_841_0\
        );

    \I__1348\ : Odrv4
    port map (
            O => \N__14883\,
            I => \this_ppu.N_841_0\
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__14878\,
            I => \this_ppu.N_841_0_cascade_\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__14875\,
            I => \N__14872\
        );

    \I__1345\ : CascadeBuf
    port map (
            O => \N__14872\,
            I => \N__14869\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__14869\,
            I => \N__14866\
        );

    \I__1343\ : InMux
    port map (
            O => \N__14866\,
            I => \N__14863\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__14863\,
            I => \this_ppu.N_669_0\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__14860\,
            I => \this_ppu.m18_i_o2_1_cascade_\
        );

    \I__1340\ : InMux
    port map (
            O => \N__14857\,
            I => \N__14851\
        );

    \I__1339\ : InMux
    port map (
            O => \N__14856\,
            I => \N__14844\
        );

    \I__1338\ : InMux
    port map (
            O => \N__14855\,
            I => \N__14844\
        );

    \I__1337\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14844\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__14851\,
            I => \this_ppu.N_426_0\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__14844\,
            I => \this_ppu.N_426_0\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__14839\,
            I => \N__14836\
        );

    \I__1333\ : InMux
    port map (
            O => \N__14836\,
            I => \N__14833\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__14833\,
            I => \M_this_vga_signals_address_2\
        );

    \I__1331\ : InMux
    port map (
            O => \N__14830\,
            I => \N__14827\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__14827\,
            I => \this_ppu.oam_cache.mem_4\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__14824\,
            I => \N__14821\
        );

    \I__1328\ : CascadeBuf
    port map (
            O => \N__14821\,
            I => \N__14818\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__14818\,
            I => \N__14815\
        );

    \I__1326\ : InMux
    port map (
            O => \N__14815\,
            I => \N__14812\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__14812\,
            I => \this_ppu.N_985_0\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__14809\,
            I => \N__14806\
        );

    \I__1323\ : CascadeBuf
    port map (
            O => \N__14806\,
            I => \N__14803\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__14803\,
            I => \N__14800\
        );

    \I__1321\ : InMux
    port map (
            O => \N__14800\,
            I => \N__14797\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__14797\,
            I => \this_ppu.N_671_0\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__14794\,
            I => \this_ppu.N_426_0_cascade_\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__14791\,
            I => \this_ppu.un1_M_oam_curr_q_1_c2_cascade_\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__14788\,
            I => \N__14785\
        );

    \I__1316\ : CascadeBuf
    port map (
            O => \N__14785\,
            I => \N__14782\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__14782\,
            I => \N__14779\
        );

    \I__1314\ : InMux
    port map (
            O => \N__14779\,
            I => \N__14776\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__14776\,
            I => \this_ppu.N_986_0\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__14773\,
            I => \this_ppu.un1_M_oam_curr_q_1_c4_cascade_\
        );

    \I__1311\ : IoInMux
    port map (
            O => \N__14770\,
            I => \N__14767\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__14767\,
            I => \N__14764\
        );

    \I__1309\ : IoSpan4Mux
    port map (
            O => \N__14764\,
            I => \N__14761\
        );

    \I__1308\ : Span4Mux_s2_h
    port map (
            O => \N__14761\,
            I => \N__14758\
        );

    \I__1307\ : Sp12to4
    port map (
            O => \N__14758\,
            I => \N__14755\
        );

    \I__1306\ : Span12Mux_s8_h
    port map (
            O => \N__14755\,
            I => \N__14752\
        );

    \I__1305\ : Odrv12
    port map (
            O => \N__14752\,
            I => rgb_c_0
        );

    \I__1304\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14746\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__14746\,
            I => \N__14743\
        );

    \I__1302\ : Span4Mux_v
    port map (
            O => \N__14743\,
            I => \N__14740\
        );

    \I__1301\ : Odrv4
    port map (
            O => \N__14740\,
            I => \M_this_oam_ram_read_data_15\
        );

    \I__1300\ : InMux
    port map (
            O => \N__14737\,
            I => \N__14734\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__14734\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_15\
        );

    \I__1298\ : InMux
    port map (
            O => \N__14731\,
            I => \N__14728\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__14728\,
            I => \this_ppu.oam_cache.N_577_0\
        );

    \I__1296\ : InMux
    port map (
            O => \N__14725\,
            I => \N__14722\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__14722\,
            I => \this_ppu.oam_cache.N_567_0\
        );

    \I__1294\ : InMux
    port map (
            O => \N__14719\,
            I => \N__14716\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__14716\,
            I => \N__14713\
        );

    \I__1292\ : Span4Mux_v
    port map (
            O => \N__14713\,
            I => \N__14710\
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__14710\,
            I => \M_this_oam_ram_read_data_8\
        );

    \I__1290\ : InMux
    port map (
            O => \N__14707\,
            I => \N__14704\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__14704\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_8\
        );

    \I__1288\ : InMux
    port map (
            O => \N__14701\,
            I => \N__14698\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__14698\,
            I => \N__14695\
        );

    \I__1286\ : Span12Mux_h
    port map (
            O => \N__14695\,
            I => \N__14692\
        );

    \I__1285\ : Odrv12
    port map (
            O => \N__14692\,
            I => \M_this_oam_ram_read_data_9\
        );

    \I__1284\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14686\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__14686\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_9\
        );

    \I__1282\ : InMux
    port map (
            O => \N__14683\,
            I => \N__14680\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__14680\,
            I => \N__14677\
        );

    \I__1280\ : Span4Mux_h
    port map (
            O => \N__14677\,
            I => \N__14674\
        );

    \I__1279\ : Span4Mux_v
    port map (
            O => \N__14674\,
            I => \N__14671\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__14671\,
            I => \M_this_oam_ram_read_data_10\
        );

    \I__1277\ : InMux
    port map (
            O => \N__14668\,
            I => \N__14665\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__14665\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_10\
        );

    \I__1275\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14659\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__14659\,
            I => \N__14656\
        );

    \I__1273\ : Span4Mux_h
    port map (
            O => \N__14656\,
            I => \N__14653\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__14653\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_16\
        );

    \I__1271\ : InMux
    port map (
            O => \N__14650\,
            I => \N__14647\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__14647\,
            I => \this_ppu.oam_cache.mem_18\
        );

    \I__1269\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14641\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__14641\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_18\
        );

    \I__1267\ : InMux
    port map (
            O => \N__14638\,
            I => \N__14635\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__14635\,
            I => \N__14632\
        );

    \I__1265\ : Odrv12
    port map (
            O => \N__14632\,
            I => port_clk_c
        );

    \I__1264\ : InMux
    port map (
            O => \N__14629\,
            I => \N__14626\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__14626\,
            I => \this_delay_clk.M_pipe_qZ0Z_0\
        );

    \I__1262\ : InMux
    port map (
            O => \N__14623\,
            I => \N__14620\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__14620\,
            I => \N__14617\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__14617\,
            I => \M_this_oam_ram_read_data_12\
        );

    \I__1259\ : InMux
    port map (
            O => \N__14614\,
            I => \N__14611\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__14611\,
            I => \N__14608\
        );

    \I__1257\ : Span4Mux_h
    port map (
            O => \N__14608\,
            I => \N__14605\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__14605\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_12\
        );

    \I__1255\ : InMux
    port map (
            O => \N__14602\,
            I => \N__14599\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__14599\,
            I => \N__14596\
        );

    \I__1253\ : Span4Mux_h
    port map (
            O => \N__14596\,
            I => \N__14593\
        );

    \I__1252\ : Odrv4
    port map (
            O => \N__14593\,
            I => \this_ppu.oam_cache.N_579_0\
        );

    \I__1251\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14587\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__14587\,
            I => \N__14584\
        );

    \I__1249\ : Span4Mux_h
    port map (
            O => \N__14584\,
            I => \N__14581\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__14581\,
            I => \M_this_oam_ram_read_data_26\
        );

    \I__1247\ : InMux
    port map (
            O => \N__14578\,
            I => \N__14575\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__14575\,
            I => \N__14572\
        );

    \I__1245\ : Odrv4
    port map (
            O => \N__14572\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_26\
        );

    \I__1244\ : IoInMux
    port map (
            O => \N__14569\,
            I => \N__14566\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__14566\,
            I => \N__14563\
        );

    \I__1242\ : IoSpan4Mux
    port map (
            O => \N__14563\,
            I => \N__14560\
        );

    \I__1241\ : Span4Mux_s1_v
    port map (
            O => \N__14560\,
            I => \N__14557\
        );

    \I__1240\ : Span4Mux_v
    port map (
            O => \N__14557\,
            I => \N__14554\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__14554\,
            I => \N_84\
        );

    \I__1238\ : IoInMux
    port map (
            O => \N__14551\,
            I => \N__14548\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__14548\,
            I => \N__14545\
        );

    \I__1236\ : Span4Mux_s2_h
    port map (
            O => \N__14545\,
            I => \N__14542\
        );

    \I__1235\ : Span4Mux_h
    port map (
            O => \N__14542\,
            I => \N__14539\
        );

    \I__1234\ : Span4Mux_v
    port map (
            O => \N__14539\,
            I => \N__14536\
        );

    \I__1233\ : Span4Mux_v
    port map (
            O => \N__14536\,
            I => \N__14533\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__14533\,
            I => rgb_c_5
        );

    \I__1231\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14527\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__14527\,
            I => \this_ppu.oam_cache.N_561_0\
        );

    \I__1229\ : InMux
    port map (
            O => \N__14524\,
            I => \N__14521\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__14521\,
            I => \N__14518\
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__14518\,
            I => \this_ppu.oam_cache.mem_17\
        );

    \I__1226\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14512\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__14512\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_17\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__14509\,
            I => \N__14506\
        );

    \I__1223\ : InMux
    port map (
            O => \N__14506\,
            I => \N__14503\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__14503\,
            I => \this_ppu.M_oam_cache_read_data_i_16\
        );

    \I__1221\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14497\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__14497\,
            I => \this_ppu.M_oam_cache_read_data_i_17\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__14494\,
            I => \N__14491\
        );

    \I__1218\ : InMux
    port map (
            O => \N__14491\,
            I => \N__14487\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__14490\,
            I => \N__14484\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__14487\,
            I => \N__14477\
        );

    \I__1215\ : InMux
    port map (
            O => \N__14484\,
            I => \N__14474\
        );

    \I__1214\ : CascadeMux
    port map (
            O => \N__14483\,
            I => \N__14471\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__14482\,
            I => \N__14467\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__14481\,
            I => \N__14463\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__14480\,
            I => \N__14460\
        );

    \I__1210\ : Span4Mux_v
    port map (
            O => \N__14477\,
            I => \N__14453\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__14474\,
            I => \N__14453\
        );

    \I__1208\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14450\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__14470\,
            I => \N__14447\
        );

    \I__1206\ : InMux
    port map (
            O => \N__14467\,
            I => \N__14443\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__14466\,
            I => \N__14440\
        );

    \I__1204\ : InMux
    port map (
            O => \N__14463\,
            I => \N__14437\
        );

    \I__1203\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14434\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__14459\,
            I => \N__14431\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__14458\,
            I => \N__14428\
        );

    \I__1200\ : Span4Mux_h
    port map (
            O => \N__14453\,
            I => \N__14423\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__14450\,
            I => \N__14423\
        );

    \I__1198\ : InMux
    port map (
            O => \N__14447\,
            I => \N__14420\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__14446\,
            I => \N__14417\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__14443\,
            I => \N__14413\
        );

    \I__1195\ : InMux
    port map (
            O => \N__14440\,
            I => \N__14410\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__14437\,
            I => \N__14404\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__14434\,
            I => \N__14404\
        );

    \I__1192\ : InMux
    port map (
            O => \N__14431\,
            I => \N__14401\
        );

    \I__1191\ : InMux
    port map (
            O => \N__14428\,
            I => \N__14398\
        );

    \I__1190\ : Span4Mux_v
    port map (
            O => \N__14423\,
            I => \N__14393\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__14420\,
            I => \N__14393\
        );

    \I__1188\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14390\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__14416\,
            I => \N__14387\
        );

    \I__1186\ : Span4Mux_s2_v
    port map (
            O => \N__14413\,
            I => \N__14380\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__14410\,
            I => \N__14380\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__14409\,
            I => \N__14377\
        );

    \I__1183\ : Span4Mux_v
    port map (
            O => \N__14404\,
            I => \N__14370\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__14401\,
            I => \N__14370\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__14398\,
            I => \N__14370\
        );

    \I__1180\ : Span4Mux_h
    port map (
            O => \N__14393\,
            I => \N__14365\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__14390\,
            I => \N__14365\
        );

    \I__1178\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14361\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__14386\,
            I => \N__14358\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__14385\,
            I => \N__14355\
        );

    \I__1175\ : Span4Mux_v
    port map (
            O => \N__14380\,
            I => \N__14352\
        );

    \I__1174\ : InMux
    port map (
            O => \N__14377\,
            I => \N__14349\
        );

    \I__1173\ : Span4Mux_v
    port map (
            O => \N__14370\,
            I => \N__14344\
        );

    \I__1172\ : Span4Mux_v
    port map (
            O => \N__14365\,
            I => \N__14344\
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__14364\,
            I => \N__14341\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__14361\,
            I => \N__14338\
        );

    \I__1169\ : InMux
    port map (
            O => \N__14358\,
            I => \N__14335\
        );

    \I__1168\ : InMux
    port map (
            O => \N__14355\,
            I => \N__14332\
        );

    \I__1167\ : Sp12to4
    port map (
            O => \N__14352\,
            I => \N__14327\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__14349\,
            I => \N__14327\
        );

    \I__1165\ : Sp12to4
    port map (
            O => \N__14344\,
            I => \N__14324\
        );

    \I__1164\ : InMux
    port map (
            O => \N__14341\,
            I => \N__14321\
        );

    \I__1163\ : Span4Mux_s3_v
    port map (
            O => \N__14338\,
            I => \N__14314\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__14335\,
            I => \N__14314\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__14332\,
            I => \N__14314\
        );

    \I__1160\ : Span12Mux_h
    port map (
            O => \N__14327\,
            I => \N__14311\
        );

    \I__1159\ : Span12Mux_s6_h
    port map (
            O => \N__14324\,
            I => \N__14306\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__14321\,
            I => \N__14306\
        );

    \I__1157\ : Span4Mux_v
    port map (
            O => \N__14314\,
            I => \N__14303\
        );

    \I__1156\ : Span12Mux_v
    port map (
            O => \N__14311\,
            I => \N__14298\
        );

    \I__1155\ : Span12Mux_h
    port map (
            O => \N__14306\,
            I => \N__14298\
        );

    \I__1154\ : Span4Mux_v
    port map (
            O => \N__14303\,
            I => \N__14295\
        );

    \I__1153\ : Odrv12
    port map (
            O => \N__14298\,
            I => \M_this_ppu_spr_addr_4\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__14295\,
            I => \M_this_ppu_spr_addr_4\
        );

    \I__1151\ : InMux
    port map (
            O => \N__14290\,
            I => \this_ppu.offset_y_cry_0\
        );

    \I__1150\ : InMux
    port map (
            O => \N__14287\,
            I => \this_ppu.offset_y_cry_1\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__14284\,
            I => \N__14277\
        );

    \I__1148\ : CascadeMux
    port map (
            O => \N__14283\,
            I => \N__14273\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__14282\,
            I => \N__14270\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__14281\,
            I => \N__14259\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__14280\,
            I => \N__14254\
        );

    \I__1144\ : InMux
    port map (
            O => \N__14277\,
            I => \N__14251\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__14276\,
            I => \N__14248\
        );

    \I__1142\ : InMux
    port map (
            O => \N__14273\,
            I => \N__14245\
        );

    \I__1141\ : InMux
    port map (
            O => \N__14270\,
            I => \N__14242\
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__14269\,
            I => \N__14239\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__14268\,
            I => \N__14236\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__14267\,
            I => \N__14233\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__14266\,
            I => \N__14230\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__14265\,
            I => \N__14227\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__14264\,
            I => \N__14224\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__14263\,
            I => \N__14221\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__14262\,
            I => \N__14218\
        );

    \I__1132\ : InMux
    port map (
            O => \N__14259\,
            I => \N__14215\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__14258\,
            I => \N__14212\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__14257\,
            I => \N__14209\
        );

    \I__1129\ : InMux
    port map (
            O => \N__14254\,
            I => \N__14206\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__14251\,
            I => \N__14203\
        );

    \I__1127\ : InMux
    port map (
            O => \N__14248\,
            I => \N__14200\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__14245\,
            I => \N__14197\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__14242\,
            I => \N__14194\
        );

    \I__1124\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14191\
        );

    \I__1123\ : InMux
    port map (
            O => \N__14236\,
            I => \N__14188\
        );

    \I__1122\ : InMux
    port map (
            O => \N__14233\,
            I => \N__14185\
        );

    \I__1121\ : InMux
    port map (
            O => \N__14230\,
            I => \N__14182\
        );

    \I__1120\ : InMux
    port map (
            O => \N__14227\,
            I => \N__14179\
        );

    \I__1119\ : InMux
    port map (
            O => \N__14224\,
            I => \N__14176\
        );

    \I__1118\ : InMux
    port map (
            O => \N__14221\,
            I => \N__14173\
        );

    \I__1117\ : InMux
    port map (
            O => \N__14218\,
            I => \N__14170\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__14215\,
            I => \N__14167\
        );

    \I__1115\ : InMux
    port map (
            O => \N__14212\,
            I => \N__14164\
        );

    \I__1114\ : InMux
    port map (
            O => \N__14209\,
            I => \N__14161\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__14206\,
            I => \N__14158\
        );

    \I__1112\ : Span12Mux_h
    port map (
            O => \N__14203\,
            I => \N__14155\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__14200\,
            I => \N__14152\
        );

    \I__1110\ : Span12Mux_s6_v
    port map (
            O => \N__14197\,
            I => \N__14147\
        );

    \I__1109\ : Span12Mux_s7_h
    port map (
            O => \N__14194\,
            I => \N__14147\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__14191\,
            I => \N__14140\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__14188\,
            I => \N__14140\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__14185\,
            I => \N__14140\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__14182\,
            I => \N__14131\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__14179\,
            I => \N__14131\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__14176\,
            I => \N__14131\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__14173\,
            I => \N__14131\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__14170\,
            I => \N__14128\
        );

    \I__1100\ : Span4Mux_s2_v
    port map (
            O => \N__14167\,
            I => \N__14121\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__14164\,
            I => \N__14121\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__14161\,
            I => \N__14121\
        );

    \I__1097\ : Span12Mux_h
    port map (
            O => \N__14158\,
            I => \N__14118\
        );

    \I__1096\ : Span12Mux_h
    port map (
            O => \N__14155\,
            I => \N__14115\
        );

    \I__1095\ : Span12Mux_h
    port map (
            O => \N__14152\,
            I => \N__14112\
        );

    \I__1094\ : Span12Mux_h
    port map (
            O => \N__14147\,
            I => \N__14109\
        );

    \I__1093\ : Span12Mux_v
    port map (
            O => \N__14140\,
            I => \N__14102\
        );

    \I__1092\ : Span12Mux_v
    port map (
            O => \N__14131\,
            I => \N__14102\
        );

    \I__1091\ : Span12Mux_s7_h
    port map (
            O => \N__14128\,
            I => \N__14102\
        );

    \I__1090\ : Span4Mux_v
    port map (
            O => \N__14121\,
            I => \N__14099\
        );

    \I__1089\ : Span12Mux_h
    port map (
            O => \N__14118\,
            I => \N__14096\
        );

    \I__1088\ : Span12Mux_v
    port map (
            O => \N__14115\,
            I => \N__14091\
        );

    \I__1087\ : Span12Mux_h
    port map (
            O => \N__14112\,
            I => \N__14091\
        );

    \I__1086\ : Span12Mux_v
    port map (
            O => \N__14109\,
            I => \N__14086\
        );

    \I__1085\ : Span12Mux_h
    port map (
            O => \N__14102\,
            I => \N__14086\
        );

    \I__1084\ : Span4Mux_v
    port map (
            O => \N__14099\,
            I => \N__14083\
        );

    \I__1083\ : Odrv12
    port map (
            O => \N__14096\,
            I => \M_this_ppu_spr_addr_5\
        );

    \I__1082\ : Odrv12
    port map (
            O => \N__14091\,
            I => \M_this_ppu_spr_addr_5\
        );

    \I__1081\ : Odrv12
    port map (
            O => \N__14086\,
            I => \M_this_ppu_spr_addr_5\
        );

    \I__1080\ : Odrv4
    port map (
            O => \N__14083\,
            I => \M_this_ppu_spr_addr_5\
        );

    \I__1079\ : InMux
    port map (
            O => \N__14074\,
            I => \N__14071\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__14071\,
            I => \this_ppu.oam_cache.mem_16\
        );

    \I__1077\ : IoInMux
    port map (
            O => \N__14068\,
            I => \N__14065\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__14065\,
            I => \this_vga_signals.N_1307_0\
        );

    \I__1075\ : IoInMux
    port map (
            O => \N__14062\,
            I => \N__14059\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__14059\,
            I => \N_428\
        );

    \I__1073\ : IoInMux
    port map (
            O => \N__14056\,
            I => \N__14053\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__14053\,
            I => \N__14050\
        );

    \I__1071\ : Span12Mux_s1_v
    port map (
            O => \N__14050\,
            I => \N__14047\
        );

    \I__1070\ : Odrv12
    port map (
            O => \N__14047\,
            I => \N_842\
        );

    \I__1069\ : IoInMux
    port map (
            O => \N__14044\,
            I => \N__14041\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__14041\,
            I => \N__14038\
        );

    \I__1067\ : IoSpan4Mux
    port map (
            O => \N__14038\,
            I => \N__14035\
        );

    \I__1066\ : Span4Mux_s3_v
    port map (
            O => \N__14035\,
            I => \N__14032\
        );

    \I__1065\ : Span4Mux_v
    port map (
            O => \N__14032\,
            I => \N__14029\
        );

    \I__1064\ : Span4Mux_v
    port map (
            O => \N__14029\,
            I => \N__14026\
        );

    \I__1063\ : Span4Mux_v
    port map (
            O => \N__14026\,
            I => \N__14023\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__14023\,
            I => rgb_c_4
        );

    \I__1061\ : IoInMux
    port map (
            O => \N__14020\,
            I => \N__14017\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__14017\,
            I => \N__14014\
        );

    \I__1059\ : IoSpan4Mux
    port map (
            O => \N__14014\,
            I => \N__14011\
        );

    \I__1058\ : IoSpan4Mux
    port map (
            O => \N__14011\,
            I => \N__14008\
        );

    \I__1057\ : Span4Mux_s3_h
    port map (
            O => \N__14008\,
            I => \N__14005\
        );

    \I__1056\ : Odrv4
    port map (
            O => \N__14005\,
            I => \M_vcounter_q_esr_RNIQ82H7_9\
        );

    \I__1055\ : InMux
    port map (
            O => \N__14002\,
            I => \N__13999\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__13999\,
            I => \N__13996\
        );

    \I__1053\ : Span4Mux_v
    port map (
            O => \N__13996\,
            I => \N__13993\
        );

    \I__1052\ : Odrv4
    port map (
            O => \N__13993\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__1051\ : InMux
    port map (
            O => \N__13990\,
            I => \N__13987\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__13987\,
            I => \N__13984\
        );

    \I__1049\ : Span4Mux_h
    port map (
            O => \N__13984\,
            I => \N__13981\
        );

    \I__1048\ : Odrv4
    port map (
            O => \N__13981\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_13\
        );

    \I__1047\ : IoInMux
    port map (
            O => \N__13978\,
            I => \N__13975\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__13975\,
            I => \N__13972\
        );

    \I__1045\ : IoSpan4Mux
    port map (
            O => \N__13972\,
            I => \N__13969\
        );

    \I__1044\ : Span4Mux_s3_h
    port map (
            O => \N__13969\,
            I => \N__13966\
        );

    \I__1043\ : Odrv4
    port map (
            O => \N__13966\,
            I => rgb_c_2
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_surface_y_d_cry_6\,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_warmup_d_cry_8\,
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_warmup_d_cry_16\,
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_warmup_d_cry_24\,
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_24_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_23_0_\
        );

    \IN_MUX_bfv_24_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_map_address_q_cry_7\,
            carryinitout => \bfn_24_24_0_\
        );

    \IN_MUX_bfv_26_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_26_21_0_\
        );

    \IN_MUX_bfv_26_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_ext_address_q_cry_7\,
            carryinitout => \bfn_26_22_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_14_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \M_this_data_count_q_cry_7\,
            carryinitout => \bfn_14_25_0_\
        );

    \IN_MUX_bfv_18_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_21_0_\
        );

    \IN_MUX_bfv_18_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            carryinitout => \bfn_18_22_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.offset_x_cry_6_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_22_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_14_0_\
        );

    \IN_MUX_bfv_22_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_spr_address_q_cry_7\,
            carryinitout => \bfn_22_15_0_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIFLF77_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14068\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_1307_0_g\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI01JU6_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__25600\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_1637_g\
        );

    \this_reset_cond.M_stage_q_RNI6VB7_3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__26116\,
            GLOBALBUFFEROUTPUT => \M_this_reset_cond_out_g_0\
        );

    \this_reset_cond.M_stage_q_RNI6VB7_0_3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21778\,
            GLOBALBUFFEROUTPUT => \N_620_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIFLF77_9_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27343\,
            in2 => \_gnd_net_\,
            in3 => \N__34225\,
            lcout => \this_vga_signals.N_1307_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.port_data_rw_i_i_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37755\,
            in2 => \_gnd_net_\,
            in3 => \N__32877\,
            lcout => \N_428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIA65T2_0_9_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39506\,
            lcout => \N_842\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__17218\,
            in1 => \N__18526\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIQ82H7_9_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__39505\,
            in1 => \N__37735\,
            in2 => \_gnd_net_\,
            in3 => \N__37813\,
            lcout => \M_vcounter_q_esr_RNIQ82H7_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24136\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14002\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18127\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17216\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17217\,
            in2 => \_gnd_net_\,
            in3 => \N__20272\,
            lcout => rgb_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24081\,
            in2 => \_gnd_net_\,
            in3 => \N__15924\,
            lcout => \this_ppu.oam_cache.N_561_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_17_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNID8M7_17_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14515\,
            lcout => \this_ppu.M_oam_cache_read_data_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_y_cry_0_c_inv_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21586\,
            in2 => \N__14509\,
            in3 => \N__20151\,
            lcout => \this_ppu.M_oam_cache_read_data_i_16\,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \this_ppu.offset_y_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_y_cry_0_c_RNIVBJT1_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000110110100"
        )
    port map (
            in0 => \N__38187\,
            in1 => \N__14500\,
            in2 => \N__21541\,
            in3 => \N__14290\,
            lcout => \M_this_ppu_spr_addr_4\,
            ltout => OPEN,
            carryin => \this_ppu.offset_y_cry_0\,
            carryout => \this_ppu.offset_y_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI2GKT1_18_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001011100001"
        )
    port map (
            in0 => \N__14644\,
            in1 => \N__38188\,
            in2 => \N__21508\,
            in3 => \N__14287\,
            lcout => \M_this_ppu_spr_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_16_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14074\,
            lcout => \this_ppu.M_oam_cache_read_data_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_18_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14650\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_0_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14638\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42102\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_1_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14629\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42102\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14623\,
            in2 => \_gnd_net_\,
            in3 => \N__24137\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16860\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24139\,
            lcout => \this_ppu.oam_cache.N_579_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14590\,
            in2 => \_gnd_net_\,
            in3 => \N__24138\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_warmup_q_0_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14945\,
            lcout => \M_this_warmup_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42116\,
            ce => 'H',
            sr => \N__43129\
        );

    \M_this_warmup_q_1_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__14946\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14961\,
            lcout => \M_this_warmup_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42116\,
            ce => 'H',
            sr => \N__43129\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__17941\,
            in1 => \N__17806\,
            in2 => \_gnd_net_\,
            in3 => \N__17874\,
            lcout => \N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17194\,
            in2 => \_gnd_net_\,
            in3 => \N__18148\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_3_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__23254\,
            in1 => \N__15277\,
            in2 => \_gnd_net_\,
            in3 => \N__17515\,
            lcout => \this_ppu.M_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42049\,
            ce => 'H',
            sr => \N__43112\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14749\,
            in2 => \_gnd_net_\,
            in3 => \N__24016\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24008\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15025\,
            lcout => \this_ppu.oam_cache.N_577_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24011\,
            in2 => \_gnd_net_\,
            in3 => \N__15007\,
            lcout => \this_ppu.oam_cache.N_567_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24009\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14719\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14701\,
            in2 => \_gnd_net_\,
            in3 => \N__24017\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24010\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14683\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24007\,
            in2 => \_gnd_net_\,
            in3 => \N__15999\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_1_3_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15728\,
            in1 => \N__15671\,
            in2 => \N__15619\,
            in3 => \N__15439\,
            lcout => \this_ppu.m35_i_0_a3_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100100101"
        )
    port map (
            in0 => \N__18342\,
            in1 => \N__18294\,
            in2 => \N__18394\,
            in3 => \N__18428\,
            lcout => \this_vga_ramdac.i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_4_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14830\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNI61SIV_1_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000101000"
        )
    port map (
            in0 => \N__14894\,
            in1 => \N__16609\,
            in2 => \N__15441\,
            in3 => \N__14857\,
            lcout => \this_ppu.N_985_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNIU85NV_2_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__15571\,
            in1 => \N__15678\,
            in2 => \_gnd_net_\,
            in3 => \N__14895\,
            lcout => \this_ppu.N_671_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIK7UCK_3_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__16566\,
            in1 => \N__22117\,
            in2 => \N__24164\,
            in3 => \N__17497\,
            lcout => \this_ppu.N_426_0\,
            ltout => \this_ppu.N_426_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNI1KGLK_1_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__16608\,
            in1 => \_gnd_net_\,
            in2 => \N__14794\,
            in3 => \N__15431\,
            lcout => \this_ppu.un1_M_oam_curr_q_1_c2\,
            ltout => \this_ppu.un1_M_oam_curr_q_1_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNINHERV_3_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100010001000"
        )
    port map (
            in0 => \N__15747\,
            in1 => \N__14896\,
            in2 => \N__14791\,
            in3 => \N__15676\,
            lcout => \this_ppu.N_986_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNII43UK_3_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15746\,
            in1 => \N__15675\,
            in2 => \_gnd_net_\,
            in3 => \N__15570\,
            lcout => \this_ppu.un1_M_oam_curr_q_1_c4\,
            ltout => \this_ppu.un1_M_oam_curr_q_1_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_4_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15615\,
            in2 => \N__14773\,
            in3 => \N__15835\,
            lcout => \M_this_ppu_oam_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42073\,
            ce => 'H',
            sr => \N__41651\
        );

    \this_ppu.M_oam_curr_q_0_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__14855\,
            in1 => \N__16624\,
            in2 => \_gnd_net_\,
            in3 => \N__15845\,
            lcout => \M_this_ppu_oam_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42086\,
            ce => 'H',
            sr => \N__41648\
        );

    \this_ppu.M_state_q_ns_11_0__m13_0_i_a3_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__23112\,
            in1 => \N__24318\,
            in2 => \_gnd_net_\,
            in3 => \N__25906\,
            lcout => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0\,
            ltout => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIVDVLA_4_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22185\,
            in2 => \N__14899\,
            in3 => \N__24429\,
            lcout => \this_ppu.M_oam_curr_qc_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI5DBTA_4_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__24428\,
            in1 => \N__43223\,
            in2 => \N__22186\,
            in3 => \N__24569\,
            lcout => \this_ppu.N_841_0\,
            ltout => \this_ppu.N_841_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNIFQIEV_0_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001010000"
        )
    port map (
            in0 => \N__14854\,
            in1 => \_gnd_net_\,
            in2 => \N__14878\,
            in3 => \N__16623\,
            lcout => \this_ppu.N_669_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m18_i_o2_1_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000101010"
        )
    port map (
            in0 => \N__29791\,
            in1 => \N__35014\,
            in2 => \N__26236\,
            in3 => \N__30699\,
            lcout => OPEN,
            ltout => \this_ppu.m18_i_o2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m18_i_o2_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__30700\,
            in1 => \N__26200\,
            in2 => \N__14860\,
            in3 => \N__34751\,
            lcout => \N_792_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_1_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000101000"
        )
    port map (
            in0 => \N__15846\,
            in1 => \N__15435\,
            in2 => \N__16632\,
            in3 => \N__14856\,
            lcout => \M_this_ppu_oam_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42086\,
            ce => 'H',
            sr => \N__41648\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIK68L03_9_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18105\,
            in2 => \_gnd_net_\,
            in3 => \N__16090\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_2_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15049\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42098\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24114\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16408\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24115\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16135\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_4_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15021\,
            in1 => \N__21636\,
            in2 => \N__15006\,
            in3 => \N__15324\,
            lcout => \this_ppu.m28_e_i_a3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14986\,
            in2 => \_gnd_net_\,
            in3 => \N__24113\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_warmup_d_cry_1_c_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14962\,
            in2 => \N__14947\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \un1_M_this_warmup_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_warmup_q_2_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14926\,
            in2 => \_gnd_net_\,
            in3 => \N__14920\,
            lcout => \M_this_warmup_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_1\,
            carryout => \un1_M_this_warmup_d_cry_2\,
            clk => \N__42105\,
            ce => 'H',
            sr => \N__43123\
        );

    \M_this_warmup_q_3_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14917\,
            in2 => \_gnd_net_\,
            in3 => \N__14911\,
            lcout => \M_this_warmup_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_2\,
            carryout => \un1_M_this_warmup_d_cry_3\,
            clk => \N__42105\,
            ce => 'H',
            sr => \N__43123\
        );

    \M_this_warmup_q_4_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14908\,
            in2 => \_gnd_net_\,
            in3 => \N__14902\,
            lcout => \M_this_warmup_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_3\,
            carryout => \un1_M_this_warmup_d_cry_4\,
            clk => \N__42105\,
            ce => 'H',
            sr => \N__43123\
        );

    \M_this_warmup_q_5_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15121\,
            in2 => \_gnd_net_\,
            in3 => \N__15115\,
            lcout => \M_this_warmup_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_4\,
            carryout => \un1_M_this_warmup_d_cry_5\,
            clk => \N__42105\,
            ce => 'H',
            sr => \N__43123\
        );

    \M_this_warmup_q_6_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15112\,
            in2 => \_gnd_net_\,
            in3 => \N__15106\,
            lcout => \M_this_warmup_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_5\,
            carryout => \un1_M_this_warmup_d_cry_6\,
            clk => \N__42105\,
            ce => 'H',
            sr => \N__43123\
        );

    \M_this_warmup_q_7_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15103\,
            in2 => \_gnd_net_\,
            in3 => \N__15097\,
            lcout => \M_this_warmup_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_6\,
            carryout => \un1_M_this_warmup_d_cry_7\,
            clk => \N__42105\,
            ce => 'H',
            sr => \N__43123\
        );

    \M_this_warmup_q_8_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15094\,
            in2 => \_gnd_net_\,
            in3 => \N__15088\,
            lcout => \M_this_warmup_qZ0Z_8\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_7\,
            carryout => \un1_M_this_warmup_d_cry_8\,
            clk => \N__42105\,
            ce => 'H',
            sr => \N__43123\
        );

    \M_this_warmup_q_9_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15085\,
            in2 => \_gnd_net_\,
            in3 => \N__15079\,
            lcout => \M_this_warmup_qZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \un1_M_this_warmup_d_cry_9\,
            clk => \N__42112\,
            ce => 'H',
            sr => \N__43126\
        );

    \M_this_warmup_q_10_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15076\,
            in2 => \_gnd_net_\,
            in3 => \N__15070\,
            lcout => \M_this_warmup_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_9\,
            carryout => \un1_M_this_warmup_d_cry_10\,
            clk => \N__42112\,
            ce => 'H',
            sr => \N__43126\
        );

    \M_this_warmup_q_11_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15067\,
            in2 => \_gnd_net_\,
            in3 => \N__15061\,
            lcout => \M_this_warmup_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_10\,
            carryout => \un1_M_this_warmup_d_cry_11\,
            clk => \N__42112\,
            ce => 'H',
            sr => \N__43126\
        );

    \M_this_warmup_q_12_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15058\,
            in2 => \_gnd_net_\,
            in3 => \N__15052\,
            lcout => \M_this_warmup_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_11\,
            carryout => \un1_M_this_warmup_d_cry_12\,
            clk => \N__42112\,
            ce => 'H',
            sr => \N__43126\
        );

    \M_this_warmup_q_13_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15199\,
            in2 => \_gnd_net_\,
            in3 => \N__15193\,
            lcout => \M_this_warmup_qZ0Z_13\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_12\,
            carryout => \un1_M_this_warmup_d_cry_13\,
            clk => \N__42112\,
            ce => 'H',
            sr => \N__43126\
        );

    \M_this_warmup_q_14_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15190\,
            in2 => \_gnd_net_\,
            in3 => \N__15184\,
            lcout => \M_this_warmup_qZ0Z_14\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_13\,
            carryout => \un1_M_this_warmup_d_cry_14\,
            clk => \N__42112\,
            ce => 'H',
            sr => \N__43126\
        );

    \M_this_warmup_q_15_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15181\,
            in2 => \_gnd_net_\,
            in3 => \N__15175\,
            lcout => \M_this_warmup_qZ0Z_15\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_14\,
            carryout => \un1_M_this_warmup_d_cry_15\,
            clk => \N__42112\,
            ce => 'H',
            sr => \N__43126\
        );

    \M_this_warmup_q_16_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15172\,
            in2 => \_gnd_net_\,
            in3 => \N__15166\,
            lcout => \M_this_warmup_qZ0Z_16\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_15\,
            carryout => \un1_M_this_warmup_d_cry_16\,
            clk => \N__42112\,
            ce => 'H',
            sr => \N__43126\
        );

    \M_this_warmup_q_17_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15163\,
            in2 => \_gnd_net_\,
            in3 => \N__15157\,
            lcout => \M_this_warmup_qZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \un1_M_this_warmup_d_cry_17\,
            clk => \N__42119\,
            ce => 'H',
            sr => \N__43130\
        );

    \M_this_warmup_q_18_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15154\,
            in2 => \_gnd_net_\,
            in3 => \N__15148\,
            lcout => \M_this_warmup_qZ0Z_18\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_17\,
            carryout => \un1_M_this_warmup_d_cry_18\,
            clk => \N__42119\,
            ce => 'H',
            sr => \N__43130\
        );

    \M_this_warmup_q_19_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15145\,
            in2 => \_gnd_net_\,
            in3 => \N__15139\,
            lcout => \M_this_warmup_qZ0Z_19\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_18\,
            carryout => \un1_M_this_warmup_d_cry_19\,
            clk => \N__42119\,
            ce => 'H',
            sr => \N__43130\
        );

    \M_this_warmup_q_20_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15136\,
            in2 => \_gnd_net_\,
            in3 => \N__15130\,
            lcout => \M_this_warmup_qZ0Z_20\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_19\,
            carryout => \un1_M_this_warmup_d_cry_20\,
            clk => \N__42119\,
            ce => 'H',
            sr => \N__43130\
        );

    \M_this_warmup_q_21_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15127\,
            in2 => \_gnd_net_\,
            in3 => \N__15265\,
            lcout => \M_this_warmup_qZ0Z_21\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_20\,
            carryout => \un1_M_this_warmup_d_cry_21\,
            clk => \N__42119\,
            ce => 'H',
            sr => \N__43130\
        );

    \M_this_warmup_q_22_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15262\,
            in2 => \_gnd_net_\,
            in3 => \N__15256\,
            lcout => \M_this_warmup_qZ0Z_22\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_21\,
            carryout => \un1_M_this_warmup_d_cry_22\,
            clk => \N__42119\,
            ce => 'H',
            sr => \N__43130\
        );

    \M_this_warmup_q_23_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15253\,
            in2 => \_gnd_net_\,
            in3 => \N__15247\,
            lcout => \M_this_warmup_qZ0Z_23\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_22\,
            carryout => \un1_M_this_warmup_d_cry_23\,
            clk => \N__42119\,
            ce => 'H',
            sr => \N__43130\
        );

    \M_this_warmup_q_24_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15244\,
            in2 => \_gnd_net_\,
            in3 => \N__15238\,
            lcout => \M_this_warmup_qZ0Z_24\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_23\,
            carryout => \un1_M_this_warmup_d_cry_24\,
            clk => \N__42119\,
            ce => 'H',
            sr => \N__43130\
        );

    \M_this_warmup_q_25_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15235\,
            in2 => \_gnd_net_\,
            in3 => \N__15229\,
            lcout => \M_this_warmup_qZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_9_25_0_\,
            carryout => \un1_M_this_warmup_d_cry_25\,
            clk => \N__42123\,
            ce => 'H',
            sr => \N__43131\
        );

    \M_this_warmup_q_26_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15226\,
            in2 => \_gnd_net_\,
            in3 => \N__15220\,
            lcout => \M_this_warmup_qZ0Z_26\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_25\,
            carryout => \un1_M_this_warmup_d_cry_26\,
            clk => \N__42123\,
            ce => 'H',
            sr => \N__43131\
        );

    \M_this_warmup_q_27_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15213\,
            in2 => \_gnd_net_\,
            in3 => \N__15217\,
            lcout => \M_this_warmup_qZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42123\,
            ce => 'H',
            sr => \N__43131\
        );

    \M_this_status_flags_q_0_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__15214\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21856\,
            lcout => \M_this_status_flags_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42123\,
            ce => 'H',
            sr => \N__43131\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_18_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26731\,
            in2 => \_gnd_net_\,
            in3 => \N__17239\,
            lcout => \M_this_oam_ram_write_data_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_23_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26734\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18163\,
            lcout => \M_this_oam_ram_write_data_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_20_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26733\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17248\,
            lcout => \M_this_oam_ram_write_data_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_19_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26732\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17068\,
            lcout => \M_this_oam_ram_write_data_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_17_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17080\,
            in2 => \_gnd_net_\,
            in3 => \N__26643\,
            lcout => \M_this_oam_ram_write_data_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18253\,
            in2 => \_gnd_net_\,
            in3 => \N__17206\,
            lcout => rgb_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24012\,
            in2 => \_gnd_net_\,
            in3 => \N__15331\,
            lcout => \this_ppu.oam_cache.N_586_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_10_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15289\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42024\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m28_e_i_o3_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__16258\,
            in1 => \N__16240\,
            in2 => \_gnd_net_\,
            in3 => \N__16201\,
            lcout => \this_ppu.N_844_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI61M7_10_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15271\,
            lcout => \this_ppu.M_oam_cache_read_data_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_cnt_q_cry_0_c_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23993\,
            in2 => \N__16053\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \this_ppu.un1_M_oam_cache_cnt_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_LUT4_0_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15794\,
            in2 => \_gnd_net_\,
            in3 => \N__15490\,
            lcout => \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_cnt_q_cry_0\,
            carryout => \this_ppu.un1_M_oam_cache_cnt_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_LUT4_0_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22643\,
            in3 => \N__15487\,
            lcout => \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_cnt_q_cry_1\,
            carryout => \this_ppu.un1_M_oam_cache_cnt_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_LUT4_0_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15523\,
            in2 => \_gnd_net_\,
            in3 => \N__15484\,
            lcout => \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_cnt_q_cry_2\,
            carryout => \this_ppu.un1_M_oam_cache_cnt_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_cache_cnt_q_4_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__15394\,
            in1 => \N__43237\,
            in2 => \N__24679\,
            in3 => \N__15481\,
            lcout => \this_ppu.M_oam_cache_cnt_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_7_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15478\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIDR5V3_7_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__39508\,
            in1 => \N__17929\,
            in2 => \N__17716\,
            in3 => \N__16705\,
            lcout => \N_41_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_0_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__15795\,
            in1 => \N__15672\,
            in2 => \N__22653\,
            in3 => \N__15440\,
            lcout => OPEN,
            ltout => \this_ppu.m62_0_a2_0_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000000000"
        )
    port map (
            in0 => \N__15393\,
            in1 => \N__15608\,
            in2 => \N__15376\,
            in3 => \N__15763\,
            lcout => \this_ppu.N_762_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_3_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000011000000"
        )
    port map (
            in0 => \N__15574\,
            in1 => \N__15733\,
            in2 => \N__15853\,
            in3 => \N__15674\,
            lcout => \M_this_ppu_oam_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42040\,
            ce => 'H',
            sr => \N__41649\
        );

    \this_ppu.M_oam_curr_q_2_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__15673\,
            in1 => \N__15847\,
            in2 => \_gnd_net_\,
            in3 => \N__15573\,
            lcout => \M_this_ppu_oam_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42040\,
            ce => 'H',
            sr => \N__41649\
        );

    \this_ppu.M_oam_curr_q_5_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__15851\,
            in1 => \N__16662\,
            in2 => \N__15620\,
            in3 => \N__15859\,
            lcout => \M_this_ppu_oam_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42040\,
            ce => 'H',
            sr => \N__41649\
        );

    \this_ppu.M_oam_curr_q_6_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100011000000"
        )
    port map (
            in0 => \N__16661\,
            in1 => \N__15852\,
            in2 => \N__18713\,
            in3 => \N__15550\,
            lcout => \this_ppu.M_oam_curr_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42040\,
            ce => 'H',
            sr => \N__41649\
        );

    \this_ppu.M_surface_x_q_RNO_0_7_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22904\,
            in1 => \N__21243\,
            in2 => \N__23004\,
            in3 => \N__23271\,
            lcout => \this_ppu.un1_M_surface_x_q_ac0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_cache_cnt_q_1_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__15790\,
            in1 => \N__43238\,
            in2 => \N__15817\,
            in3 => \N__24581\,
            lcout => \this_ppu.M_oam_cache_cnt_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m62_0_a2_0_o2_1_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__15737\,
            in1 => \N__16607\,
            in2 => \N__15527\,
            in3 => \N__16048\,
            lcout => \this_ppu.m62_0_a2_0_o2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNO_0_6_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15732\,
            in1 => \N__15677\,
            in2 => \N__15621\,
            in3 => \N__15572\,
            lcout => \this_ppu.un1_M_oam_curr_q_1_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_cache_cnt_q_3_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__15544\,
            in1 => \N__43239\,
            in2 => \N__15528\,
            in3 => \N__24582\,
            lcout => \this_ppu.M_oam_cache_cnt_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__24134\,
            in1 => \N__15961\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_2_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15937\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_3_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15925\,
            in2 => \_gnd_net_\,
            in3 => \N__16752\,
            lcout => \this_ppu.m28_e_i_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010010001011"
        )
    port map (
            in0 => \N__17317\,
            in1 => \N__16098\,
            in2 => \N__18996\,
            in3 => \N__15867\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI8I4KS3_1_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111010000001"
        )
    port map (
            in0 => \N__17379\,
            in1 => \N__17319\,
            in2 => \N__15898\,
            in3 => \N__16066\,
            lcout => \this_vga_signals.haddress_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m1_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000111011110"
        )
    port map (
            in0 => \N__17318\,
            in1 => \N__16099\,
            in2 => \N__18997\,
            in3 => \N__15868\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_m2_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110100110100"
        )
    port map (
            in0 => \N__16921\,
            in1 => \N__17383\,
            in2 => \N__15895\,
            in3 => \N__17425\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un89_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI4NUA8C_1_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__18091\,
            in1 => \N__16809\,
            in2 => \N__15892\,
            in3 => \N__15889\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17605\,
            in2 => \_gnd_net_\,
            in3 => \N__16955\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000000000"
        )
    port map (
            in0 => \N__18553\,
            in1 => \N__19042\,
            in2 => \N__18061\,
            in3 => \N__16966\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un68_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m2_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16102\,
            in3 => \N__19120\,
            lcout => \this_vga_signals.if_m2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m18_i_a2_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__16233\,
            in1 => \N__16254\,
            in2 => \N__23249\,
            in3 => \N__16194\,
            lcout => \this_ppu.N_1394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIDPGC47_9_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18096\,
            in1 => \N__16089\,
            in2 => \_gnd_net_\,
            in3 => \N__16813\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19126\,
            in2 => \_gnd_net_\,
            in3 => \N__16958\,
            lcout => \this_vga_signals.mult1_un75_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_cache_cnt_q_0_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__24135\,
            in1 => \N__43240\,
            in2 => \N__16049\,
            in3 => \N__24580\,
            lcout => \this_ppu.M_oam_cache_cnt_qZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI1INF21_9_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18097\,
            in2 => \_gnd_net_\,
            in3 => \N__16959\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_0_c_inv_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15973\,
            in2 => \N__21585\,
            in3 => \N__16000\,
            lcout => \this_ppu.M_this_oam_ram_read_data_i_16\,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => \this_ppu.un1_oam_data_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_1_c_inv_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15967\,
            in2 => \N__21540\,
            in3 => \N__17010\,
            lcout => \this_ppu.M_this_oam_ram_read_data_i_17\,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_0\,
            carryout => \this_ppu.un1_oam_data_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_2_c_inv_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16270\,
            in2 => \N__21504\,
            in3 => \N__16182\,
            lcout => \this_ppu.M_this_oam_ram_read_data_i_18\,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_1\,
            carryout => \this_ppu.un1_oam_data_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_2_c_RNIR4HD_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16324\,
            in2 => \N__21468\,
            in3 => \N__16264\,
            lcout => \this_ppu.un1_oam_data_1_cry_2_c_RNIR4HDZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_2\,
            carryout => \this_ppu.un1_oam_data_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_3_c_RNIT7ID_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16537\,
            in2 => \N__21423\,
            in3 => \N__16261\,
            lcout => \this_ppu.un1_oam_data_1_cry_3_c_RNIT7IDZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_3\,
            carryout => \this_ppu.un1_oam_data_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJD_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21378\,
            in2 => \N__16384\,
            in3 => \N__16243\,
            lcout => \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_4\,
            carryout => \this_ppu.un1_oam_data_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKD_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21330\,
            in2 => \N__16111\,
            in3 => \N__16222\,
            lcout => \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_5\,
            carryout => \this_ppu.un1_oam_data_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m28_e_i_o3_2_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000001"
        )
    port map (
            in0 => \N__17059\,
            in1 => \N__16219\,
            in2 => \N__16213\,
            in3 => \N__16204\,
            lcout => \this_ppu.m28_e_i_o3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24172\,
            in2 => \_gnd_net_\,
            in3 => \N__16183\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_5_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26761\,
            in2 => \_gnd_net_\,
            in3 => \N__17992\,
            lcout => \M_this_oam_ram_write_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16134\,
            lcout => \M_this_oam_ram_read_data_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__24173\,
            in1 => \N__16432\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16407\,
            lcout => \M_this_oam_ram_read_data_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__24174\,
            in1 => \N__16375\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16339\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24175\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16338\,
            lcout => \M_this_oam_ram_read_data_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_10_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16975\,
            in2 => \_gnd_net_\,
            in3 => \N__26747\,
            lcout => \M_this_oam_ram_write_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIML464_9_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__17875\,
            in1 => \N__16477\,
            in2 => \N__17805\,
            in3 => \N__17937\,
            lcout => \N_260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16294\,
            in2 => \_gnd_net_\,
            in3 => \N__24171\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_9_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17137\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26748\,
            lcout => \M_this_oam_ram_write_data_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17583\,
            lcout => \M_this_oam_ram_read_data_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_28_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40783\,
            in2 => \_gnd_net_\,
            in3 => \N__26726\,
            lcout => \M_this_oam_ram_write_data_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_8_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17143\,
            in2 => \_gnd_net_\,
            in3 => \N__26728\,
            lcout => \M_this_oam_ram_write_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_31_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26727\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39870\,
            lcout => \M_this_oam_ram_write_data_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_16_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26730\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17086\,
            lcout => \M_this_oam_ram_write_data_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_24_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42416\,
            in2 => \_gnd_net_\,
            in3 => \N__26729\,
            lcout => \M_this_oam_ram_write_data_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIOC7D3_6_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110011"
        )
    port map (
            in0 => \N__17431\,
            in1 => \N__16438\,
            in2 => \N__19224\,
            in3 => \N__17707\,
            lcout => \this_vga_signals.hsync_1_i_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16465\,
            in2 => \_gnd_net_\,
            in3 => \N__24140\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI69GD1_0_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__17443\,
            in1 => \N__17358\,
            in2 => \N__18620\,
            in3 => \N__17417\,
            lcout => \this_vga_signals.hsync_1_i_0_0_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000110010111"
        )
    port map (
            in0 => \N__18353\,
            in1 => \N__18303\,
            in2 => \N__18404\,
            in3 => \N__18437\,
            lcout => \this_vga_ramdac.m16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110110100011"
        )
    port map (
            in0 => \N__18438\,
            in1 => \N__18354\,
            in2 => \N__18307\,
            in3 => \N__18398\,
            lcout => \this_vga_ramdac.m19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17773\,
            in2 => \_gnd_net_\,
            in3 => \N__17855\,
            lcout => \this_vga_signals.N_811_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18211\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17207\,
            lcout => rgb_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_1_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__16660\,
            in1 => \N__16631\,
            in2 => \_gnd_net_\,
            in3 => \N__16576\,
            lcout => \this_ppu.N_1196_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNITMA41_9_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__17854\,
            in1 => \N__17915\,
            in2 => \N__30472\,
            in3 => \N__17769\,
            lcout => \this_vga_signals.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_1_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010001"
        )
    port map (
            in0 => \N__26135\,
            in1 => \N__16819\,
            in2 => \N__24183\,
            in3 => \N__16567\,
            lcout => \this_ppu.M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42032\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIF4AR_5_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__17702\,
            in1 => \N__18594\,
            in2 => \_gnd_net_\,
            in3 => \N__17914\,
            lcout => \this_vga_signals.M_hcounter_d7_0_i_0_o3_0_o3_4_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101000101000"
        )
    port map (
            in0 => \N__17844\,
            in1 => \N__17905\,
            in2 => \N__17784\,
            in3 => \N__17701\,
            lcout => \this_vga_signals.N_291_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m28_e_i_a3_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__16864\,
            in1 => \N__16840\,
            in2 => \N__16786\,
            in3 => \N__16828\,
            lcout => \this_ppu.N_1184_7\,
            ltout => \this_ppu.N_1184_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m18_i_1_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100110011"
        )
    port map (
            in0 => \N__24270\,
            in1 => \N__16720\,
            in2 => \N__16822\,
            in3 => \N__23250\,
            lcout => \this_ppu.m18_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_2_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16711\,
            in1 => \N__16930\,
            in2 => \N__17956\,
            in3 => \N__16960\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_12_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16798\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42041\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16785\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24095\,
            lcout => \this_ppu.oam_cache.N_569_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24094\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16753\,
            lcout => \this_ppu.oam_cache.N_575_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m18_i_a3_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__23113\,
            in1 => \N__24319\,
            in2 => \N__21885\,
            in3 => \N__25916\,
            lcout => \this_ppu.N_1182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100101011"
        )
    port map (
            in0 => \N__17635\,
            in1 => \N__17305\,
            in2 => \N__17378\,
            in3 => \N__17604\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_9_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011010011111"
        )
    port map (
            in0 => \N__16957\,
            in1 => \N__19122\,
            in2 => \N__16714\,
            in3 => \N__17320\,
            lcout => \this_vga_signals.mult1_un82_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__19225\,
            in1 => \N__19149\,
            in2 => \_gnd_net_\,
            in3 => \N__19030\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_2\,
            ltout => \this_vga_signals.mult1_un68_sum_ac0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_1_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100111111"
        )
    port map (
            in0 => \N__19119\,
            in1 => \N__17616\,
            in2 => \N__16969\,
            in3 => \N__17634\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010111011"
        )
    port map (
            in0 => \N__19121\,
            in1 => \N__17306\,
            in2 => \_gnd_net_\,
            in3 => \N__16956\,
            lcout => \this_vga_signals.mult1_un75_sum_c2_0\,
            ltout => \this_vga_signals.mult1_un75_sum_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_x4_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17952\,
            in2 => \N__16924\,
            in3 => \N__19123\,
            lcout => \this_vga_signals.if_N_8_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_3_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16915\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42063\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI8F2M3_9_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__17787\,
            in1 => \N__17870\,
            in2 => \N__39507\,
            in3 => \N__17930\,
            lcout => \N_852_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16903\,
            in2 => \_gnd_net_\,
            in3 => \N__24163\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_0_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16876\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.IO_port_data_write_0_a2_i_o2_1_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__29248\,
            in1 => \N__27172\,
            in2 => \N__36358\,
            in3 => \N__29290\,
            lcout => \this_vga_signals.N_834_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_y_q_esr_RNICCL8_7_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21705\,
            in2 => \_gnd_net_\,
            in3 => \N__21672\,
            lcout => \this_ppu.un1_oam_data_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_6_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17035\,
            in2 => \_gnd_net_\,
            in3 => \N__26759\,
            lcout => \M_this_oam_ram_write_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_6_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40415\,
            lcout => \M_this_data_tmp_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42087\,
            ce => \N__25686\,
            sr => \N__43119\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_7_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17017\,
            in2 => \_gnd_net_\,
            in3 => \N__26760\,
            lcout => \M_this_oam_ram_write_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_7_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39926\,
            lcout => \M_this_data_tmp_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42087\,
            ce => \N__25686\,
            sr => \N__43119\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24177\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17011\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_11_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41513\,
            lcout => \M_this_data_tmp_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42099\,
            ce => \N__26563\,
            sr => \N__43122\
        );

    \M_this_data_tmp_q_esr_10_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__42796\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42099\,
            ce => \N__26563\,
            sr => \N__43122\
        );

    \M_this_data_tmp_q_esr_15_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39927\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42099\,
            ce => \N__26563\,
            sr => \N__43122\
        );

    \M_this_data_tmp_q_esr_8_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42429\,
            lcout => \M_this_data_tmp_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42099\,
            ce => \N__26563\,
            sr => \N__43122\
        );

    \M_this_data_tmp_q_esr_9_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39760\,
            lcout => \M_this_data_tmp_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42099\,
            ce => \N__26563\,
            sr => \N__43122\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_26_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__42792\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26722\,
            lcout => \M_this_oam_ram_write_data_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_27_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41512\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26723\,
            lcout => \M_this_oam_ram_write_data_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_30_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40435\,
            in2 => \_gnd_net_\,
            in3 => \N__26724\,
            lcout => \M_this_oam_ram_write_data_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_15_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26725\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17104\,
            lcout => \M_this_oam_ram_write_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_16_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42415\,
            lcout => \M_this_data_tmp_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42113\,
            ce => \N__25632\,
            sr => \N__43127\
        );

    \M_this_data_tmp_q_esr_17_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39728\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42113\,
            ce => \N__25632\,
            sr => \N__43127\
        );

    \M_this_data_tmp_q_esr_19_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__41511\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42113\,
            ce => \N__25632\,
            sr => \N__43127\
        );

    \M_this_data_tmp_q_esr_20_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40782\,
            lcout => \M_this_data_tmp_qZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42113\,
            ce => \N__25632\,
            sr => \N__43127\
        );

    \M_this_data_tmp_q_esr_18_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42791\,
            lcout => \M_this_data_tmp_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42113\,
            ce => \N__25632\,
            sr => \N__43127\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_0_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18154\,
            in2 => \_gnd_net_\,
            in3 => \N__26642\,
            lcout => \M_this_oam_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_q_ret_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__20307\,
            in1 => \N__18109\,
            in2 => \N__17193\,
            in3 => \N__26136\,
            lcout => \this_vga_ramdac.N_852_i_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41998\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17284\,
            in2 => \_gnd_net_\,
            in3 => \N__19072\,
            lcout => \this_vga_signals.N_298_0\,
            ltout => \this_vga_signals.N_298_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__17345\,
            in1 => \N__17408\,
            in2 => \N__17158\,
            in3 => \N__19209\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_1044_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__17155\,
            in1 => \N__17785\,
            in2 => \N__17146\,
            in3 => \N__17853\,
            lcout => \this_vga_signals.M_hcounter_d7_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_1_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__27296\,
            in1 => \_gnd_net_\,
            in2 => \N__17418\,
            in3 => \N__17346\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42005\,
            ce => 'H',
            sr => \N__18682\
        );

    \this_vga_signals.M_hcounter_q_0_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17409\,
            in2 => \_gnd_net_\,
            in3 => \N__27295\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42005\,
            ce => 'H',
            sr => \N__18682\
        );

    \this_vga_signals.M_hcounter_q_RNIADGD1_1_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__17347\,
            in1 => \N__17442\,
            in2 => \N__18619\,
            in3 => \N__19210\,
            lcout => \this_vga_signals.hsync_1_i_0_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17416\,
            in2 => \N__17368\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27291\,
            in1 => \N__17304\,
            in2 => \_gnd_net_\,
            in3 => \N__17269\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__42016\,
            ce => 'H',
            sr => \N__18681\
        );

    \this_vga_signals.M_hcounter_q_3_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27344\,
            in1 => \N__19118\,
            in2 => \_gnd_net_\,
            in3 => \N__17266\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__42016\,
            ce => 'H',
            sr => \N__18681\
        );

    \this_vga_signals.M_hcounter_q_4_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27292\,
            in1 => \N__19211\,
            in2 => \_gnd_net_\,
            in3 => \N__17263\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__42016\,
            ce => 'H',
            sr => \N__18681\
        );

    \this_vga_signals.M_hcounter_q_5_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27345\,
            in1 => \N__18603\,
            in2 => \_gnd_net_\,
            in3 => \N__17260\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \N__42016\,
            ce => 'H',
            sr => \N__18681\
        );

    \this_vga_signals.M_hcounter_q_6_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27293\,
            in1 => \N__17706\,
            in2 => \_gnd_net_\,
            in3 => \N__17257\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \N__42016\,
            ce => 'H',
            sr => \N__18681\
        );

    \this_vga_signals.M_hcounter_q_7_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27346\,
            in1 => \N__17916\,
            in2 => \_gnd_net_\,
            in3 => \N__17254\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \N__42016\,
            ce => 'H',
            sr => \N__18681\
        );

    \this_vga_signals.M_hcounter_q_8_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27294\,
            in1 => \N__17856\,
            in2 => \_gnd_net_\,
            in3 => \N__17251\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \N__42016\,
            ce => 'H',
            sr => \N__18681\
        );

    \this_vga_signals.M_hcounter_q_esr_9_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17774\,
            in2 => \_gnd_net_\,
            in3 => \N__17527\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42025\,
            ce => \N__18649\,
            sr => \N__18674\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_1_0_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111010011"
        )
    port map (
            in0 => \N__19216\,
            in1 => \N__17649\,
            in2 => \N__18621\,
            in3 => \N__17709\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17521\,
            in2 => \N__17524\,
            in3 => \N__17727\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_tz_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__18610\,
            in1 => \N__19215\,
            in2 => \_gnd_net_\,
            in3 => \N__17708\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_0_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI42MR5_6_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000111"
        )
    port map (
            in0 => \N__17508\,
            in1 => \N__23222\,
            in2 => \N__23836\,
            in3 => \N__23786\,
            lcout => \this_ppu.un1_M_state_q_7_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24096\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17488\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI83M7_12_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17464\,
            lcout => \this_ppu.M_oam_cache_read_data_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_15_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17458\,
            lcout => \this_ppu.M_oam_cache_read_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42033\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_0_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011101100"
        )
    port map (
            in0 => \N__17656\,
            in1 => \N__17728\,
            in2 => \N__18622\,
            in3 => \N__17712\,
            lcout => \this_vga_signals.mult1_un54_sum_c3\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb2_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__19028\,
            in1 => \N__18549\,
            in2 => \N__17959\,
            in3 => \N__19150\,
            lcout => \this_vga_signals.mult1_un68_sum_axb2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010000111"
        )
    port map (
            in0 => \N__19151\,
            in1 => \N__19029\,
            in2 => \N__19125\,
            in3 => \N__19222\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101100100100"
        )
    port map (
            in0 => \N__17920\,
            in1 => \N__17860\,
            in2 => \N__17786\,
            in3 => \N__17710\,
            lcout => \this_vga_signals.N_968\,
            ltout => \this_vga_signals.N_968_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111011111"
        )
    port map (
            in0 => \N__17711\,
            in1 => \N__18614\,
            in2 => \N__17659\,
            in3 => \N__17655\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19027\,
            in2 => \N__17638\,
            in3 => \N__19221\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1\,
            ltout => \this_vga_signals.mult1_un68_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001111101100"
        )
    port map (
            in0 => \N__19108\,
            in1 => \N__17626\,
            in2 => \N__17620\,
            in3 => \N__17617\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24181\,
            in2 => \_gnd_net_\,
            in3 => \N__17590\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_13_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17551\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNILTV6A_9_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__19041\,
            in1 => \_gnd_net_\,
            in2 => \N__18104\,
            in3 => \N__19153\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNINGAC6_9_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__18092\,
            in1 => \N__18057\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_0_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19256\,
            lcout => \this_pixel_clk_M_counter_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42064\,
            ce => 'H',
            sr => \N__43116\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_3_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18016\,
            in2 => \_gnd_net_\,
            in3 => \N__26739\,
            lcout => \M_this_oam_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_3_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__41515\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42076\,
            ce => \N__25685\,
            sr => \N__43117\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_4_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17998\,
            in2 => \_gnd_net_\,
            in3 => \N__26740\,
            lcout => \M_this_oam_ram_write_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_4_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40785\,
            lcout => \M_this_data_tmp_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42076\,
            ce => \N__25685\,
            sr => \N__43117\
        );

    \M_this_data_tmp_q_esr_5_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__40058\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42088\,
            ce => \N__25687\,
            sr => \N__43120\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_29_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40059\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26719\,
            lcout => \M_this_oam_ram_write_data_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_21_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18169\,
            in2 => \_gnd_net_\,
            in3 => \N__26721\,
            lcout => \M_this_oam_ram_write_data_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_1_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26720\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20227\,
            lcout => \M_this_oam_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_25_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39729\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26718\,
            lcout => \M_this_oam_ram_write_data_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_21_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40060\,
            lcout => \M_this_data_tmp_qZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42106\,
            ce => \N__25631\,
            sr => \N__43124\
        );

    \M_this_data_tmp_q_esr_23_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39931\,
            lcout => \M_this_data_tmp_qZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42106\,
            ce => \N__25631\,
            sr => \N__43124\
        );

    \M_this_data_tmp_q_esr_0_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42377\,
            lcout => \M_this_data_tmp_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42114\,
            ce => \N__25681\,
            sr => \N__43128\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__18454\,
            in1 => \N__20308\,
            in2 => \N__18147\,
            in3 => \N__26115\,
            lcout => \this_vga_ramdac.N_3856_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41992\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101100111"
        )
    port map (
            in0 => \N__18301\,
            in1 => \N__18349\,
            in2 => \N__18409\,
            in3 => \N__18447\,
            lcout => OPEN,
            ltout => \this_vga_ramdac.i2_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100000010"
        )
    port map (
            in0 => \N__20304\,
            in1 => \N__26075\,
            in2 => \N__18130\,
            in3 => \N__18120\,
            lcout => \this_vga_ramdac.N_3858_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41999\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.G_535_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__19240\,
            in1 => \N__19263\,
            in2 => \_gnd_net_\,
            in3 => \N__43217\,
            lcout => \G_535\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000100"
        )
    port map (
            in0 => \N__18300\,
            in1 => \N__18348\,
            in2 => \_gnd_net_\,
            in3 => \N__18446\,
            lcout => \this_vga_ramdac.N_24_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000111111"
        )
    port map (
            in0 => \N__18448\,
            in1 => \N__18408\,
            in2 => \N__18355\,
            in3 => \N__18302\,
            lcout => OPEN,
            ltout => \this_vga_ramdac.m6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000101110"
        )
    port map (
            in0 => \N__18249\,
            in1 => \N__20303\,
            in2 => \N__18256\,
            in3 => \N__26077\,
            lcout => \this_vga_ramdac.N_3857_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41999\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_9_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18238\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42006\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_RNIB85C3_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__22686\,
            in1 => \N__20341\,
            in2 => \_gnd_net_\,
            in3 => \N__27061\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_pcounter_q_ret_RNIB85CZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNILVU44_1_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__27280\,
            in1 => \_gnd_net_\,
            in2 => \N__18229\,
            in3 => \N__19327\,
            lcout => \this_vga_signals.N_3_0\,
            ltout => \this_vga_signals.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_RNIOILK7_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__20366\,
            in1 => \_gnd_net_\,
            in2 => \N__18226\,
            in3 => \N__18196\,
            lcout => \M_pcounter_q_ret_1_RNIOILK7\,
            ltout => \M_pcounter_q_ret_1_RNIOILK7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__18223\,
            in1 => \N__18207\,
            in2 => \N__18214\,
            in3 => \N__26074\,
            lcout => \this_vga_ramdac.N_3859_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42006\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_RNIAI4F3_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__20342\,
            in1 => \N__27279\,
            in2 => \N__20370\,
            in3 => \N__27062\,
            lcout => \this_vga_signals.N_2_0\,
            ltout => \this_vga_signals.N_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18538\,
            in3 => \N__22707\,
            lcout => \this_vga_signals.N_1417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42006\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__26073\,
            in1 => \N__18535\,
            in2 => \N__18525\,
            in3 => \N__20306\,
            lcout => \this_vga_ramdac.N_3860_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42006\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_14_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18508\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m35_i_0_a3_0_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18714\,
            in2 => \_gnd_net_\,
            in3 => \N__21916\,
            lcout => OPEN,
            ltout => \this_ppu.m35_i_0_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_4_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010110011"
        )
    port map (
            in0 => \N__18730\,
            in1 => \N__21967\,
            in2 => \N__18496\,
            in3 => \N__26086\,
            lcout => \this_ppu.M_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNIUU07_9_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18493\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.M_oam_cache_read_data_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_11_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18487\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_1_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18472\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNIA5M7_14_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18460\,
            lcout => \this_ppu.M_oam_cache_read_data_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_2_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__18729\,
            in1 => \N__18715\,
            in2 => \N__43252\,
            in3 => \N__21917\,
            lcout => \this_ppu.M_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI94M7_13_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18691\,
            lcout => \this_ppu.M_oam_cache_read_data_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIRSG13_9_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27082\,
            in2 => \_gnd_net_\,
            in3 => \N__27312\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNIRSG13Z0Z_9\,
            ltout => \this_vga_signals.M_hcounter_q_esr_RNIRSG13Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__27313\,
            in1 => \_gnd_net_\,
            in2 => \N__18652\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.N_1307_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_8_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18643\,
            lcout => \this_ppu.M_oam_cache_read_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42026\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI72M7_11_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18628\,
            lcout => \this_ppu.M_oam_cache_read_data_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m68_0_o2_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__21208\,
            in1 => \N__21145\,
            in2 => \N__21277\,
            in3 => \N__20437\,
            lcout => \this_ppu.N_82_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_0_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__21592\,
            in1 => \N__26118\,
            in2 => \_gnd_net_\,
            in3 => \N__24615\,
            lcout => \this_ppu.M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_0_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18618\,
            in2 => \_gnd_net_\,
            in3 => \N__19220\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_1_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__19239\,
            in1 => \N__19267\,
            in2 => \_gnd_net_\,
            in3 => \N__43248\,
            lcout => \this_pixel_clk_M_counter_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNII1437_3_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__19223\,
            in1 => \N__19152\,
            in2 => \N__19124\,
            in3 => \N__19034\,
            lcout => \this_vga_signals.M_hcounter_q_RNII1437Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m18_i_a3_1_0_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24250\,
            in2 => \_gnd_net_\,
            in3 => \N__30468\,
            lcout => \this_ppu.N_1182_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_ctle_7_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26117\,
            in2 => \_gnd_net_\,
            in3 => \N__24614\,
            lcout => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_1_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__24182\,
            in1 => \N__18979\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_3_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18949\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42042\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_RNI8FJF7_4_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__37330\,
            in1 => \N__39485\,
            in2 => \N__22474\,
            in3 => \N__37747\,
            lcout => \this_ppu.M_screen_y_q_RNI8FJF7Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_4_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__24678\,
            in1 => \N__22967\,
            in2 => \N__25822\,
            in3 => \N__23275\,
            lcout => \M_this_ppu_map_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42053\,
            ce => 'H',
            sr => \N__43114\
        );

    \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20200\,
            in1 => \N__38177\,
            in2 => \_gnd_net_\,
            in3 => \N__18934\,
            lcout => \read_data_RNI5QFJ1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI62LG1_16_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__38176\,
            in1 => \N__21572\,
            in2 => \_gnd_net_\,
            in3 => \N__20158\,
            lcout => \M_this_ppu_spr_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19951\,
            in1 => \N__38175\,
            in2 => \_gnd_net_\,
            in3 => \N__41374\,
            lcout => \read_data_RNI6RFJ1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__38178\,
            in1 => \N__19723\,
            in2 => \_gnd_net_\,
            in3 => \N__43612\,
            lcout => \read_data_RNI7SFJ1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19537\,
            in1 => \N__38174\,
            in2 => \_gnd_net_\,
            in3 => \N__43747\,
            lcout => \read_data_RNI9TFJ1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_1_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__22693\,
            in1 => \N__20350\,
            in2 => \_gnd_net_\,
            in3 => \N__27101\,
            lcout => \this_vga_signals.M_pcounter_q_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42065\,
            ce => \N__27335\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_11_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19315\,
            in2 => \_gnd_net_\,
            in3 => \N__26735\,
            lcout => \M_this_oam_ram_write_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_12_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26736\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20239\,
            lcout => \M_this_oam_ram_write_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_13_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21598\,
            in2 => \_gnd_net_\,
            in3 => \N__26737\,
            lcout => \M_this_oam_ram_write_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_14_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26738\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20233\,
            lcout => \M_this_oam_ram_write_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_12_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40763\,
            lcout => \M_this_data_tmp_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42077\,
            ce => \N__26559\,
            sr => \N__43118\
        );

    \M_this_data_tmp_q_esr_14_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40443\,
            lcout => \M_this_data_tmp_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42077\,
            ce => \N__26559\,
            sr => \N__43118\
        );

    \M_this_data_tmp_q_esr_1_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39686\,
            lcout => \M_this_data_tmp_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42089\,
            ce => \N__25668\,
            sr => \N__43121\
        );

    \M_this_data_tmp_q_esr_2_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42764\,
            lcout => \M_this_data_tmp_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42089\,
            ce => \N__25668\,
            sr => \N__43121\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_22_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20206\,
            in2 => \_gnd_net_\,
            in3 => \N__26641\,
            lcout => \M_this_oam_ram_write_data_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_22_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40444\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42107\,
            ce => \N__25633\,
            sr => \N__43125\
        );

    \this_vga_signals.IO_port_data_write_0_a2_i_1_LC_13_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43665\,
            in2 => \_gnd_net_\,
            in3 => \N__20199\,
            lcout => \N_724_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20420\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41993\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__20421\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20164\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41993\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20422\,
            in2 => \_gnd_net_\,
            in3 => \N__20428\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41993\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_8_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000011000100"
        )
    port map (
            in0 => \N__23081\,
            in1 => \N__22129\,
            in2 => \N__21991\,
            in3 => \N__24430\,
            lcout => \this_ppu.M_state_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__20412\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20380\,
            lcout => \M_this_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_0_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__20346\,
            in1 => \N__27297\,
            in2 => \N__20371\,
            in3 => \N__27103\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__20320\,
            in1 => \N__20305\,
            in2 => \N__20265\,
            in3 => \N__26076\,
            lcout => \this_vga_ramdac.N_3861_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNII6H51_6_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23818\,
            in1 => \N__23614\,
            in2 => \N__23083\,
            in3 => \N__22160\,
            lcout => \this_ppu.N_785_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_4_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110010001100"
        )
    port map (
            in0 => \N__37259\,
            in1 => \N__37318\,
            in2 => \N__24682\,
            in3 => \N__37289\,
            lcout => \this_ppu.M_screen_y_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42007\,
            ce => 'H',
            sr => \N__43107\
        );

    \this_ppu.M_screen_y_q_0_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__24677\,
            in1 => \N__22384\,
            in2 => \N__22401\,
            in3 => \N__37260\,
            lcout => \M_this_ppu_vram_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42007\,
            ce => 'H',
            sr => \N__43107\
        );

    \this_ppu.M_surface_x_q_7_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__24668\,
            in1 => \N__21167\,
            in2 => \N__25780\,
            in3 => \N__20248\,
            lcout => \M_this_ppu_map_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42007\,
            ce => 'H',
            sr => \N__43107\
        );

    \this_ppu.M_surface_x_q_1_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__25753\,
            in1 => \N__24669\,
            in2 => \N__23317\,
            in3 => \N__23425\,
            lcout => \this_ppu.M_surface_x_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42007\,
            ce => 'H',
            sr => \N__43107\
        );

    \this_ppu.M_surface_x_q_6_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__24667\,
            in1 => \N__21238\,
            in2 => \N__25795\,
            in3 => \N__21940\,
            lcout => \M_this_ppu_map_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42007\,
            ce => 'H',
            sr => \N__43107\
        );

    \this_ppu.M_surface_x_q_0_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010011001"
        )
    port map (
            in0 => \N__23455\,
            in1 => \N__21963\,
            in2 => \N__25765\,
            in3 => \N__24674\,
            lcout => \this_ppu.offset_x\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42007\,
            ce => 'H',
            sr => \N__43107\
        );

    \this_ppu.oam_cache.read_data_RNIB6J72_8_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000010100"
        )
    port map (
            in0 => \N__38151\,
            in1 => \N__23453\,
            in2 => \N__20905\,
            in3 => \N__23454\,
            lcout => \M_this_ppu_spr_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_3_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__21949\,
            in1 => \N__24670\,
            in2 => \N__23400\,
            in3 => \N__25831\,
            lcout => \M_this_ppu_map_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42007\,
            ce => 'H',
            sr => \N__43107\
        );

    \this_ppu.offset_x_cry_0_c_inv_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20890\,
            in2 => \N__23467\,
            in3 => \N__20901\,
            lcout => \this_ppu.M_oam_cache_read_data_i_8\,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \this_ppu.offset_x_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_0_c_RNI5N4U1_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000110110100"
        )
    port map (
            in0 => \N__38150\,
            in1 => \N__20884\,
            in2 => \N__23316\,
            in3 => \N__20680\,
            lcout => \M_this_ppu_spr_addr_1\,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_0\,
            carryout => \this_ppu.offset_x_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_1_c_RNIFSQU1_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000110110100"
        )
    port map (
            in0 => \N__38163\,
            in1 => \N__20677\,
            in2 => \N__23353\,
            in3 => \N__20446\,
            lcout => \M_this_ppu_spr_addr_2\,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_1\,
            carryout => \this_ppu.offset_x_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m68_0_o2_0_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010001000001"
        )
    port map (
            in0 => \N__21292\,
            in1 => \N__20443\,
            in2 => \N__23397\,
            in3 => \N__20431\,
            lcout => \this_ppu.m68_0_o2_0\,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_2\,
            carryout => \this_ppu.offset_x_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_3_c_RNI3UBP_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21301\,
            in2 => \N__22997\,
            in3 => \N__21286\,
            lcout => \this_ppu.offset_x_4\,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_3\,
            carryout => \this_ppu.offset_x_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_4_c_RNI62DP_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21283\,
            in2 => \N__22914\,
            in3 => \N__21268\,
            lcout => \this_ppu.offset_x_5\,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_4\,
            carryout => \this_ppu.offset_x_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_5_c_RNI96EP_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21265\,
            in2 => \N__21242\,
            in3 => \N__21202\,
            lcout => \this_ppu.offset_x_6\,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_5\,
            carryout => \this_ppu.offset_x_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_6_c_THRU_CRY_0_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24933\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_6\,
            carryout => \this_ppu.offset_x_cry_6_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_6_c_RNICAFP_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__21199\,
            in1 => \N__21171\,
            in2 => \_gnd_net_\,
            in3 => \N__21148\,
            lcout => \this_ppu.offset_x_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNI453Q6_1_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22079\,
            in2 => \_gnd_net_\,
            in3 => \N__37237\,
            lcout => \this_ppu.M_screen_y_q_esr_RNI453Q6Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNII6H51_1_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23064\,
            in1 => \N__21918\,
            in2 => \N__23671\,
            in3 => \N__23610\,
            lcout => \this_ppu.un30_0_a2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIJ1SE_10_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23200\,
            in2 => \_gnd_net_\,
            in3 => \N__22164\,
            lcout => \this_ppu.N_999_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m13_0_i_1_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011000010000"
        )
    port map (
            in0 => \N__22165\,
            in1 => \N__23202\,
            in2 => \N__24263\,
            in3 => \N__24422\,
            lcout => \this_ppu.m13_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CRY_0_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37238\,
            in2 => \N__37255\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_y_q_esr_0_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22345\,
            in2 => \N__22207\,
            in3 => \N__21550\,
            lcout => \this_ppu.offset_y\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_0\,
            clk => \N__42035\,
            ce => \N__37169\,
            sr => \N__43110\
        );

    \this_ppu.M_surface_y_q_esr_1_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21547\,
            in2 => \N__22198\,
            in3 => \N__21511\,
            lcout => \this_ppu.M_surface_y_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_0\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_1\,
            clk => \N__42035\,
            ce => \N__37169\,
            sr => \N__43110\
        );

    \this_ppu.M_surface_y_q_esr_2_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21685\,
            in2 => \N__22483\,
            in3 => \N__21478\,
            lcout => \this_ppu.M_surface_y_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_1\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_2\,
            clk => \N__42035\,
            ce => \N__37169\,
            sr => \N__43110\
        );

    \this_ppu.M_surface_y_q_esr_3_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23680\,
            in2 => \N__23697\,
            in3 => \N__21436\,
            lcout => \M_this_ppu_map_addr_5\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_2\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_3\,
            clk => \N__42035\,
            ce => \N__37169\,
            sr => \N__43110\
        );

    \this_ppu.M_surface_y_q_esr_4_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21433\,
            in2 => \N__22470\,
            in3 => \N__21391\,
            lcout => \M_this_ppu_map_addr_6\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_3\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_4\,
            clk => \N__42035\,
            ce => \N__37169\,
            sr => \N__43110\
        );

    \this_ppu.M_surface_y_q_esr_5_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37060\,
            in2 => \N__37086\,
            in3 => \N__21346\,
            lcout => \M_this_ppu_map_addr_7\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_4\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_5\,
            clk => \N__42035\,
            ce => \N__37169\,
            sr => \N__43110\
        );

    \this_ppu.M_surface_y_q_esr_6_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34597\,
            in2 => \N__34614\,
            in3 => \N__21304\,
            lcout => \M_this_ppu_map_addr_8\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_5\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_6\,
            clk => \N__42035\,
            ce => \N__37169\,
            sr => \N__43110\
        );

    \this_ppu.M_surface_y_q_esr_7_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__22447\,
            in1 => \N__37254\,
            in2 => \N__22102\,
            in3 => \N__21727\,
            lcout => \M_this_ppu_map_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42043\,
            ce => \N__37176\,
            sr => \N__43113\
        );

    \this_ppu.M_screen_y_q_esr_1_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__22080\,
            in1 => \N__22403\,
            in2 => \_gnd_net_\,
            in3 => \N__37253\,
            lcout => \this_ppu.M_screen_y_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42043\,
            ce => \N__37176\,
            sr => \N__43113\
        );

    \this_ppu.M_screen_y_q_esr_2_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010100000"
        )
    port map (
            in0 => \N__37251\,
            in1 => \N__22081\,
            in2 => \N__22030\,
            in3 => \N__22404\,
            lcout => \this_ppu.M_screen_y_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42043\,
            ce => \N__37176\,
            sr => \N__43113\
        );

    \this_ppu.M_screen_y_q_esr_RNI563Q6_2_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22025\,
            in2 => \_gnd_net_\,
            in3 => \N__37250\,
            lcout => \this_ppu.M_screen_y_q_esr_RNI563Q6Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_3_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__37252\,
            in1 => \N__23736\,
            in2 => \N__22009\,
            in3 => \N__22054\,
            lcout => \this_ppu.M_screen_y_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42043\,
            ce => \N__37176\,
            sr => \N__43113\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24179\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21676\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24178\,
            in2 => \_gnd_net_\,
            in3 => \N__21640\,
            lcout => \this_ppu.oam_cache.N_581_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_13_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40069\,
            lcout => \M_this_data_tmp_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42054\,
            ce => \N__26558\,
            sr => \N__43115\
        );

    \M_this_data_count_q_cry_c_0_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22426\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => \M_this_data_count_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_0_THRU_LUT4_0_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22588\,
            in2 => \N__25018\,
            in3 => \N__21754\,
            lcout => \M_this_data_count_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_0\,
            carryout => \M_this_data_count_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_1_THRU_LUT4_0_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24950\,
            in2 => \N__22567\,
            in3 => \N__21751\,
            lcout => \M_this_data_count_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_1\,
            carryout => \M_this_data_count_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_2_THRU_LUT4_0_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22541\,
            in2 => \N__25019\,
            in3 => \N__21748\,
            lcout => \M_this_data_count_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_2\,
            carryout => \M_this_data_count_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_3_THRU_LUT4_0_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24954\,
            in2 => \N__22747\,
            in3 => \N__21745\,
            lcout => \M_this_data_count_q_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_3\,
            carryout => \M_this_data_count_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_4_THRU_LUT4_0_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22764\,
            in2 => \N__25020\,
            in3 => \N__21742\,
            lcout => \M_this_data_count_q_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_4\,
            carryout => \M_this_data_count_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_5_THRU_LUT4_0_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24958\,
            in2 => \N__25717\,
            in3 => \N__21739\,
            lcout => \M_this_data_count_q_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_5\,
            carryout => \M_this_data_count_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_6_THRU_LUT4_0_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25741\,
            in2 => \N__25021\,
            in3 => \N__21736\,
            lcout => \M_this_data_count_q_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_6\,
            carryout => \M_this_data_count_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_8_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22777\,
            in2 => \N__24887\,
            in3 => \N__21733\,
            lcout => \M_this_data_count_q_s_8\,
            ltout => OPEN,
            carryin => \bfn_14_25_0_\,
            carryout => \M_this_data_count_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_8_THRU_LUT4_0_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25390\,
            in2 => \N__24890\,
            in3 => \N__21730\,
            lcout => \M_this_data_count_q_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_8\,
            carryout => \M_this_data_count_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_10_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22795\,
            in2 => \N__24886\,
            in3 => \N__21826\,
            lcout => \M_this_data_count_q_s_10\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_9\,
            carryout => \M_this_data_count_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_10_THRU_LUT4_0_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22825\,
            in2 => \N__24889\,
            in3 => \N__21823\,
            lcout => \M_this_data_count_q_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_10\,
            carryout => \M_this_data_count_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_11_THRU_LUT4_0_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22842\,
            in2 => \N__24888\,
            in3 => \N__21820\,
            lcout => \M_this_data_count_q_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_11\,
            carryout => \M_this_data_count_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_13_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22809\,
            in2 => \_gnd_net_\,
            in3 => \N__21817\,
            lcout => \M_this_data_count_q_s_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_7_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__26457\,
            in1 => \N__27489\,
            in2 => \N__21807\,
            in3 => \N__22726\,
            lcout => \M_this_oam_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42090\,
            ce => 'H',
            sr => \N__41640\
        );

    \this_vga_signals.IO_port_data_write_i_m2_i_m2_0_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__38233\,
            in1 => \N__43664\,
            in2 => \_gnd_net_\,
            in3 => \N__21878\,
            lcout => \IO_port_data_write_i_m2_i_m2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43218\,
            lcout => \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m48_i_0_a3_0_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__40479\,
            in1 => \N__22180\,
            in2 => \_gnd_net_\,
            in3 => \N__24423\,
            lcout => \this_ppu.N_1202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_9_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21760\,
            in2 => \_gnd_net_\,
            in3 => \N__43242\,
            lcout => \this_ppu.M_state_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41994\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNIU3I91_3_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__23172\,
            in1 => \N__23751\,
            in2 => \_gnd_net_\,
            in3 => \N__34454\,
            lcout => \this_ppu.N_1426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_6_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__21987\,
            in1 => \N__23074\,
            in2 => \_gnd_net_\,
            in3 => \N__43244\,
            lcout => \this_ppu.M_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42001\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m35_i_0_o3_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__23609\,
            in1 => \N__34368\,
            in2 => \_gnd_net_\,
            in3 => \N__23653\,
            lcout => \this_ppu.N_91_0\,
            ltout => \this_ppu.N_91_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_RNIN4DCD_1_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23346\,
            in1 => \N__23312\,
            in2 => \N__21952\,
            in3 => \N__23461\,
            lcout => \this_ppu.un1_M_surface_x_q_c3\,
            ltout => \this_ppu.un1_M_surface_x_q_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_RNO_0_6_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22887\,
            in1 => \N__22986\,
            in2 => \N__21943\,
            in3 => \N__23390\,
            lcout => \this_ppu.un1_M_surface_x_q_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_5_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__26129\,
            in1 => \N__21832\,
            in2 => \N__21934\,
            in3 => \N__22116\,
            lcout => \this_ppu.M_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42008\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIRJK11_1_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21922\,
            in1 => \N__23665\,
            in2 => \N__24176\,
            in3 => \N__24218\,
            lcout => \this_ppu.un1_M_pixel_cnt_d_1_sqmuxa_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_10_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100010"
        )
    port map (
            in0 => \N__24219\,
            in1 => \N__26130\,
            in2 => \N__21889\,
            in3 => \N__24681\,
            lcout => \this_ppu.M_state_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42008\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m48_i_0_a3_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23822\,
            in2 => \_gnd_net_\,
            in3 => \N__23793\,
            lcout => \this_ppu.N_1201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_8_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100110"
        )
    port map (
            in0 => \N__23073\,
            in1 => \N__22181\,
            in2 => \N__40480\,
            in3 => \N__43233\,
            lcout => \this_ppu.M_state_q_srsts_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNII1FQB_7_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23596\,
            in2 => \_gnd_net_\,
            in3 => \N__34374\,
            lcout => \this_ppu.N_1145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_7_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__37236\,
            in1 => \N__36594\,
            in2 => \N__22098\,
            in3 => \N__22039\,
            lcout => \this_ppu.M_screen_y_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42018\,
            ce => \N__37165\,
            sr => \N__43108\
        );

    \this_ppu.M_screen_y_q_esr_RNIQ8BT6_1_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22078\,
            in1 => \N__22394\,
            in2 => \_gnd_net_\,
            in3 => \N__37234\,
            lcout => \this_ppu.un3_M_screen_y_d_0_c2\,
            ltout => \this_ppu.un3_M_screen_y_d_0_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNI5MHHK_3_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37235\,
            in1 => \N__23750\,
            in2 => \N__22045\,
            in3 => \N__22002\,
            lcout => \this_ppu.un3_M_screen_y_d_0_c4\,
            ltout => \this_ppu.un3_M_screen_y_d_0_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNO_0_7_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37135\,
            in2 => \N__22042\,
            in3 => \N__37329\,
            lcout => \this_ppu.un3_M_screen_y_d_0_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI467N6_8_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__26368\,
            in1 => \N__37730\,
            in2 => \_gnd_net_\,
            in3 => \N__28038\,
            lcout => \N_861_0\,
            ltout => \N_861_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNI563Q6_0_2_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22033\,
            in3 => \N__22029\,
            lcout => \this_ppu.un3_M_screen_y_d_a_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_2_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__24665\,
            in1 => \N__26131\,
            in2 => \N__22233\,
            in3 => \N__23481\,
            lcout => \M_this_ppu_vram_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42027\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_RNIQ9FQ6_0_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22402\,
            in2 => \_gnd_net_\,
            in3 => \N__37233\,
            lcout => \this_ppu.M_screen_y_q_RNIQ9FQ6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_RNI5A3DD_2_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22224\,
            in1 => \N__23156\,
            in2 => \_gnd_net_\,
            in3 => \N__23479\,
            lcout => \this_ppu.un1_M_screen_x_q_c4\,
            ltout => \this_ppu.un1_M_screen_x_q_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_4_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22313\,
            in2 => \N__22339\,
            in3 => \N__23769\,
            lcout => \M_this_ppu_vram_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42027\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_5_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__23771\,
            in1 => \N__22281\,
            in2 => \N__22320\,
            in3 => \N__22336\,
            lcout => \M_this_ppu_vram_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42027\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_RNO_0_6_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23480\,
            in1 => \N__22225\,
            in2 => \N__23170\,
            in3 => \N__22312\,
            lcout => OPEN,
            ltout => \this_ppu.un1_M_screen_x_q_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_6_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__23772\,
            in1 => \N__22254\,
            in2 => \N__22297\,
            in3 => \N__22280\,
            lcout => \M_this_ppu_vram_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42027\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_3_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100000000000"
        )
    port map (
            in0 => \N__23482\,
            in1 => \N__22229\,
            in2 => \N__23171\,
            in3 => \N__23770\,
            lcout => \M_this_ppu_vram_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42027\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_scroll_q_esr_0_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42439\,
            lcout => \M_this_scroll_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42036\,
            ce => \N__26341\,
            sr => \N__43111\
        );

    \M_this_scroll_q_esr_1_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39753\,
            lcout => \M_this_scroll_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42036\,
            ce => \N__26341\,
            sr => \N__43111\
        );

    \M_this_scroll_q_esr_2_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42765\,
            lcout => \M_this_scroll_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42036\,
            ce => \N__26341\,
            sr => \N__43111\
        );

    \M_this_scroll_q_esr_3_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41514\,
            lcout => \M_this_scroll_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42036\,
            ce => \N__26341\,
            sr => \N__43111\
        );

    \M_this_scroll_q_esr_4_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__40784\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42036\,
            ce => \N__26341\,
            sr => \N__43111\
        );

    \M_this_scroll_q_esr_5_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40068\,
            lcout => \M_this_scroll_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42036\,
            ce => \N__26341\,
            sr => \N__43111\
        );

    \M_this_scroll_q_esr_6_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40411\,
            lcout => \M_this_scroll_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42036\,
            ce => \N__26341\,
            sr => \N__43111\
        );

    \M_this_scroll_q_esr_7_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39856\,
            lcout => \M_this_scroll_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42036\,
            ce => \N__26341\,
            sr => \N__43111\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__27853\,
            in1 => \N__27397\,
            in2 => \N__34768\,
            in3 => \N__35012\,
            lcout => this_vga_signals_vsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_o2_12_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43470\,
            in2 => \_gnd_net_\,
            in3 => \N__29285\,
            lcout => \N_1005_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_9_16_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22562\,
            in1 => \N__22586\,
            in2 => \N__22542\,
            in3 => \N__22424\,
            lcout => \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_0_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__22425\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27537\,
            lcout => \M_this_data_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42055\,
            ce => \N__25358\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_1_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__27538\,
            in1 => \N__22594\,
            in2 => \_gnd_net_\,
            in3 => \N__22587\,
            lcout => \M_this_data_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42055\,
            ce => \N__25358\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_2_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__22573\,
            in1 => \N__22563\,
            in2 => \_gnd_net_\,
            in3 => \N__27539\,
            lcout => \M_this_data_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42055\,
            ce => \N__25358\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_3_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000101"
        )
    port map (
            in0 => \N__27540\,
            in1 => \_gnd_net_\,
            in2 => \N__22543\,
            in3 => \N__22549\,
            lcout => \M_this_data_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42055\,
            ce => \N__25358\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_4_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__22522\,
            in1 => \N__27541\,
            in2 => \_gnd_net_\,
            in3 => \N__22746\,
            lcout => \M_this_data_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42055\,
            ce => \N__25358\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_5_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__27542\,
            in1 => \N__22516\,
            in2 => \_gnd_net_\,
            in3 => \N__22765\,
            lcout => \M_this_data_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42055\,
            ce => \N__25358\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_6_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__22510\,
            in1 => \N__25715\,
            in2 => \_gnd_net_\,
            in3 => \N__27543\,
            lcout => \M_this_data_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42055\,
            ce => \N__25358\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_11_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__27545\,
            in1 => \N__22504\,
            in2 => \_gnd_net_\,
            in3 => \N__22824\,
            lcout => \M_this_data_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42066\,
            ce => \N__25366\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_10_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22498\,
            in1 => \N__27544\,
            in2 => \N__43529\,
            in3 => \N__28138\,
            lcout => \M_this_data_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42066\,
            ce => \N__25366\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_12_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000101"
        )
    port map (
            in0 => \N__27546\,
            in1 => \_gnd_net_\,
            in2 => \N__22843\,
            in3 => \N__22489\,
            lcout => \M_this_data_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42066\,
            ce => \N__25366\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_13_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__22852\,
            in1 => \N__27547\,
            in2 => \N__33170\,
            in3 => \N__43249\,
            lcout => \M_this_data_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42066\,
            ce => \N__25366\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_8_16_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22838\,
            in1 => \N__22823\,
            in2 => \N__22810\,
            in3 => \N__22794\,
            lcout => \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_8_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__22783\,
            in1 => \N__27548\,
            in2 => \N__27490\,
            in3 => \N__43250\,
            lcout => \M_this_data_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42066\,
            ce => \N__25366\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_7_16_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22776\,
            in1 => \N__22763\,
            in2 => \N__25389\,
            in3 => \N__22742\,
            lcout => \this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNO_0_7_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26923\,
            in1 => \N__26988\,
            in2 => \N__26514\,
            in3 => \N__26943\,
            lcout => \un1_M_this_oam_address_q_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3SF72_9_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__30541\,
            in1 => \N__22720\,
            in2 => \_gnd_net_\,
            in3 => \N__30589\,
            lcout => \this_vga_signals.g0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22708\,
            lcout => \this_vga_signals.M_pcounter_q_i_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41990\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_cache_cnt_q_2_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__22669\,
            in1 => \N__43236\,
            in2 => \N__22636\,
            in3 => \N__24666\,
            lcout => \this_ppu.M_oam_cache_cnt_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41990\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNO_0_0_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000101"
        )
    port map (
            in0 => \N__30467\,
            in1 => \_gnd_net_\,
            in2 => \N__25891\,
            in3 => \N__25968\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_lcounter_q_e_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_0_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110001010101010"
        )
    port map (
            in0 => \N__25932\,
            in1 => \N__27334\,
            in2 => \N__23038\,
            in3 => \N__27102\,
            lcout => \this_vga_signals_M_lcounter_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41990\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m18_i_o2_2_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__25887\,
            in1 => \N__25931\,
            in2 => \_gnd_net_\,
            in3 => \N__25855\,
            lcout => \this_ppu.N_838_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNICH7OC_11_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__24220\,
            in1 => \N__23658\,
            in2 => \N__39952\,
            in3 => \N__23017\,
            lcout => \N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNII1FQB_0_7_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__23611\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34369\,
            lcout => \this_ppu.N_1198\,
            ltout => \this_ppu.N_1198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_RNINHSUC_1_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__23311\,
            in1 => \N__23657\,
            in2 => \N__23011\,
            in3 => \N__23466\,
            lcout => \this_ppu.un1_M_surface_x_q_c2\,
            ltout => \this_ppu.un1_M_surface_x_q_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_RNO_0_5_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23399\,
            in1 => \N__22987\,
            in2 => \N__22930\,
            in3 => \N__23344\,
            lcout => OPEN,
            ltout => \this_ppu.un1_M_surface_x_q_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_5_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__24675\,
            in1 => \N__25804\,
            in2 => \N__22927\,
            in3 => \N__22888\,
            lcout => \M_this_ppu_map_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41991\,
            ce => 'H',
            sr => \N__43105\
        );

    \this_ppu.M_surface_x_q_2_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__22858\,
            in1 => \N__24676\,
            in2 => \N__25840\,
            in3 => \N__23345\,
            lcout => \this_ppu.M_surface_x_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41991\,
            ce => 'H',
            sr => \N__43105\
        );

    \this_ppu.M_state_q_RNIOVBHC_9_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__34370\,
            in1 => \N__23612\,
            in2 => \N__23666\,
            in3 => \N__23465\,
            lcout => \this_ppu.un1_M_surface_x_q_c1\,
            ltout => \this_ppu.un1_M_surface_x_q_c1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_RNIOOTPD_1_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23398\,
            in1 => \N__23343\,
            in2 => \N__23320\,
            in3 => \N__23310\,
            lcout => \this_ppu.un1_M_surface_x_q_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_11_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__23203\,
            in1 => \N__24424\,
            in2 => \_gnd_net_\,
            in3 => \N__43243\,
            lcout => \this_ppu.M_state_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41997\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI41OT_10_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24142\,
            in1 => \N__23242\,
            in2 => \N__24223\,
            in3 => \N__23201\,
            lcout => \this_ppu.N_798_0\,
            ltout => \this_ppu.N_798_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNIDPQ54_3_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__23166\,
            in1 => \N__23752\,
            in2 => \N__23128\,
            in3 => \N__34306\,
            lcout => \M_this_ppu_vram_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_3_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000010010001000"
        )
    port map (
            in0 => \N__25310\,
            in1 => \N__25528\,
            in2 => \N__25288\,
            in3 => \N__25483\,
            lcout => \this_ppu.M_pixel_cnt_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41997\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_595_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__24311\,
            in1 => \N__23111\,
            in2 => \N__26141\,
            in3 => \N__25917\,
            lcout => \this_ppu.N_1659_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIPR8F3_5_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__24341\,
            in1 => \N__23602\,
            in2 => \N__23082\,
            in3 => \N__24401\,
            lcout => \this_ppu.M_pixel_cnt_q_600_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_m2_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111011"
        )
    port map (
            in0 => \N__26170\,
            in1 => \N__28483\,
            in2 => \N__25990\,
            in3 => \N__25975\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIKTRBBJ2_6_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__23866\,
            in1 => \N__28363\,
            in2 => \N__23857\,
            in3 => \N__27796\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_7_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__23835\,
            in1 => \N__26128\,
            in2 => \_gnd_net_\,
            in3 => \N__23797\,
            lcout => \this_ppu.M_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42004\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_0_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__23886\,
            in1 => \N__25508\,
            in2 => \_gnd_net_\,
            in3 => \N__25463\,
            lcout => \this_ppu.M_pixel_cnt_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42015\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_RNIF1DJ_7_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24693\,
            in2 => \_gnd_net_\,
            in3 => \N__23885\,
            lcout => \this_ppu.M_state_d30_i_i_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_0_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__23553\,
            in1 => \N__23498\,
            in2 => \N__26142\,
            in3 => \N__24664\,
            lcout => \M_this_ppu_vram_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42015\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_1_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100011000000"
        )
    port map (
            in0 => \N__23499\,
            in1 => \N__23773\,
            in2 => \N__23535\,
            in3 => \N__23554\,
            lcout => \M_this_ppu_vram_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42015\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNIF77F7_3_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23749\,
            in1 => \N__39459\,
            in2 => \N__23698\,
            in3 => \N__37740\,
            lcout => \this_ppu.M_screen_y_q_esr_RNIF77F7Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIB9B9C_11_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011111110"
        )
    port map (
            in0 => \N__23667\,
            in1 => \N__24221\,
            in2 => \N__23613\,
            in3 => \N__34375\,
            lcout => \this_ppu.N_61_0\,
            ltout => \this_ppu.N_61_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_RNIM77RC_1_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23528\,
            in2 => \N__23515\,
            in3 => \N__23497\,
            lcout => \this_ppu.un1_M_screen_x_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_RNIS5KD2_3_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__25311\,
            in1 => \N__24520\,
            in2 => \N__25441\,
            in3 => \N__24436\,
            lcout => \this_ppu.N_79_0\,
            ltout => \this_ppu.N_79_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_7_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101111"
        )
    port map (
            in0 => \N__24343\,
            in1 => \_gnd_net_\,
            in2 => \N__24367\,
            in3 => \N__24526\,
            lcout => \this_ppu.M_pixel_cnt_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42023\,
            ce => 'H',
            sr => \N__43109\
        );

    \this_ppu.M_state_q_RNIKF0ID_1_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__24364\,
            in1 => \N__24229\,
            in2 => \N__24355\,
            in3 => \N__26137\,
            lcout => \this_ppu.N_1730_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIQ0NP8_0_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010100000101"
        )
    port map (
            in0 => \N__24342\,
            in1 => \N__24301\,
            in2 => \N__24271\,
            in3 => \N__25585\,
            lcout => \this_ppu.N_1042_0\,
            ltout => \this_ppu.N_1042_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIV84EA_11_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24222\,
            in1 => \N__24180\,
            in2 => \N__23908\,
            in3 => \N__23905\,
            lcout => \this_ppu.N_677_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_c_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23890\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_THRU_LUT4_0_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24504\,
            in2 => \N__25073\,
            in3 => \N__23872\,
            lcout => \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_pixel_cnt_q_1_cry_0_s1\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1_THRU_LUT4_0_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25009\,
            in2 => \N__24478\,
            in3 => \N__23869\,
            lcout => \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_pixel_cnt_q_1_cry_1_s1\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1_THRU_LUT4_0_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25312\,
            in2 => \N__25074\,
            in3 => \N__25273\,
            lcout => \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_pixel_cnt_q_1_cry_2_s1\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1_THRU_LUT4_0_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25013\,
            in2 => \N__25439\,
            in3 => \N__25270\,
            lcout => \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_pixel_cnt_q_1_cry_3_s1\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1_THRU_LUT4_0_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24451\,
            in2 => \N__25075\,
            in3 => \N__25267\,
            lcout => \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_pixel_cnt_q_1_cry_4_s1\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1_THRU_LUT4_0_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25017\,
            in2 => \N__25555\,
            in3 => \N__24697\,
            lcout => \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_pixel_cnt_q_1_cry_5_s1\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_RNO_0_7_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001001"
        )
    port map (
            in0 => \N__24694\,
            in1 => \N__25462\,
            in2 => \N__24680\,
            in3 => \N__24529\,
            lcout => \this_ppu.N_1205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_RNIU2Q61_1_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24449\,
            in1 => \N__24473\,
            in2 => \N__25550\,
            in3 => \N__24500\,
            lcout => \this_ppu.M_state_d30_i_i_o2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_1_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000001010100000"
        )
    port map (
            in0 => \N__25523\,
            in1 => \N__24511\,
            in2 => \N__24505\,
            in3 => \N__25478\,
            lcout => \this_ppu.M_pixel_cnt_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_2_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100011000000000"
        )
    port map (
            in0 => \N__25479\,
            in1 => \N__24474\,
            in2 => \N__24487\,
            in3 => \N__25524\,
            lcout => \this_ppu.M_pixel_cnt_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_5_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000001010001000"
        )
    port map (
            in0 => \N__25526\,
            in1 => \N__24450\,
            in2 => \N__24460\,
            in3 => \N__25481\,
            lcout => \this_ppu.M_pixel_cnt_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_16_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__26265\,
            in1 => \N__26283\,
            in2 => \_gnd_net_\,
            in3 => \N__26253\,
            lcout => \this_ppu.N_1301\,
            ltout => \this_ppu.N_1301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_data_count_qlde_i_0_i_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111101"
        )
    port map (
            in0 => \N__27562\,
            in1 => \N__35785\,
            in2 => \N__25564\,
            in3 => \N__37438\,
            lcout => \N_231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_6_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001000000000"
        )
    port map (
            in0 => \N__25482\,
            in1 => \N__25561\,
            in2 => \N__25551\,
            in3 => \N__25527\,
            lcout => \this_ppu.M_pixel_cnt_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_4_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000001010100000"
        )
    port map (
            in0 => \N__25525\,
            in1 => \N__25492\,
            in2 => \N__25440\,
            in3 => \N__25480\,
            lcout => \this_ppu.M_pixel_cnt_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_7_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__25411\,
            in1 => \N__25737\,
            in2 => \_gnd_net_\,
            in3 => \N__27549\,
            lcout => \M_this_data_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42050\,
            ce => \N__25365\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_9_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__27550\,
            in1 => \N__25399\,
            in2 => \_gnd_net_\,
            in3 => \N__25388\,
            lcout => \M_this_data_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42050\,
            ce => \N__25365\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a3_0_a3_2_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26674\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25339\,
            lcout => \M_this_oam_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNIQFR31_2_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26876\,
            in1 => \N__26838\,
            in2 => \N__26403\,
            in3 => \N__26791\,
            lcout => \un1_M_this_oam_address_q_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_10_16_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__25733\,
            in1 => \N__25716\,
            in2 => \_gnd_net_\,
            in3 => \N__25693\,
            lcout => \this_ppu.M_this_state_q_srsts_i_a2_10Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI13IA1_1_1_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__26839\,
            in1 => \N__26792\,
            in2 => \N__26888\,
            in3 => \N__43226\,
            lcout => \N_1709_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI13IA1_1_LC_16_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__43227\,
            in1 => \N__26880\,
            in2 => \N__26797\,
            in3 => \N__26840\,
            lcout => \N_1693_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI01JU6_9_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27298\,
            in1 => \N__27074\,
            in2 => \N__25969\,
            in3 => \N__30466\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNI01JU6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un30_0_a2_i_a2_1_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35142\,
            in1 => \N__35004\,
            in2 => \N__26235\,
            in3 => \N__30687\,
            lcout => OPEN,
            ltout => \this_ppu.N_1269_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un30_0_a2_i_o2_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__26357\,
            in1 => \N__26199\,
            in2 => \N__25588\,
            in3 => \N__30588\,
            lcout => \this_ppu.N_1006_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_8_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__35141\,
            in1 => \N__30686\,
            in2 => \N__30451\,
            in3 => \N__30173\,
            lcout => \N_782_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_6_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011111"
        )
    port map (
            in0 => \N__29760\,
            in1 => \_gnd_net_\,
            in2 => \N__29718\,
            in3 => \N__28261\,
            lcout => \this_vga_signals.N_1264\,
            ltout => \this_vga_signals.N_1264_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_ns_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25846\,
            in2 => \N__25573\,
            in3 => \N__25570\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_4_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_x0_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__29706\,
            in1 => \N__29838\,
            in2 => \N__29766\,
            in3 => \N__29619\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_4_1_0_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_1_0_x1_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__29618\,
            in1 => \N__29756\,
            in2 => \N__29849\,
            in3 => \N__29707\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_4_1_0_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_scroll_q_esr_10_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42772\,
            lcout => \M_this_scroll_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42002\,
            ce => \N__26326\,
            sr => \N__43104\
        );

    \M_this_scroll_q_esr_11_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41474\,
            lcout => \M_this_scroll_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42002\,
            ce => \N__26326\,
            sr => \N__43104\
        );

    \M_this_scroll_q_esr_12_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40786\,
            lcout => \M_this_scroll_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42002\,
            ce => \N__26326\,
            sr => \N__43104\
        );

    \M_this_scroll_q_esr_13_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40039\,
            lcout => \M_this_scroll_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42002\,
            ce => \N__26326\,
            sr => \N__43104\
        );

    \M_this_scroll_q_esr_14_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40420\,
            lcout => \M_this_scroll_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42002\,
            ce => \N__26326\,
            sr => \N__43104\
        );

    \M_this_scroll_q_esr_15_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39906\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42002\,
            ce => \N__26326\,
            sr => \N__43104\
        );

    \M_this_scroll_q_esr_8_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__42449\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42002\,
            ce => \N__26326\,
            sr => \N__43104\
        );

    \M_this_scroll_q_esr_9_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39782\,
            lcout => \M_this_scroll_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42002\,
            ce => \N__26326\,
            sr => \N__43104\
        );

    \this_vga_signals.un5_vaddress_g0_14_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__29320\,
            in1 => \N__28524\,
            in2 => \N__27163\,
            in3 => \N__27151\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c3_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_7_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__25981\,
            in1 => \N__28664\,
            in2 => \N__25993\,
            in3 => \N__27817\,
            lcout => \this_vga_signals.N_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_x2_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28930\,
            in2 => \_gnd_net_\,
            in3 => \N__27433\,
            lcout => \this_vga_signals.g0_0_x2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m1_0_x2_1_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28931\,
            in1 => \N__27828\,
            in2 => \_gnd_net_\,
            in3 => \N__27004\,
            lcout => \this_vga_signals.if_m1_0_x2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_4_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__34973\,
            in1 => \N__35321\,
            in2 => \N__26228\,
            in3 => \N__30581\,
            lcout => \this_vga_signals.N_836_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_33_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110000111001"
        )
    port map (
            in0 => \N__28904\,
            in1 => \N__28957\,
            in2 => \N__35491\,
            in3 => \N__27124\,
            lcout => \this_vga_signals.r_N_2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNO_0_1_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100001011010"
        )
    port map (
            in0 => \N__27116\,
            in1 => \N__25961\,
            in2 => \N__25885\,
            in3 => \N__30453\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_1043_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_1_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011000100"
        )
    port map (
            in0 => \N__27333\,
            in1 => \N__25879\,
            in2 => \N__25942\,
            in3 => \N__25939\,
            lcout => \this_vga_signals_M_lcounter_q_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42019\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25938\,
            in1 => \N__25918\,
            in2 => \N__25886\,
            in3 => \N__30454\,
            lcout => \this_ppu.M_last_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42019\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__28903\,
            in1 => \N__27425\,
            in2 => \N__35490\,
            in3 => \N__27026\,
            lcout => \N_771_0\,
            ltout => \N_771_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m18_i_o2_3_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__35301\,
            in1 => \_gnd_net_\,
            in2 => \N__26203\,
            in3 => \N__34993\,
            lcout => \this_ppu.N_774_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__34994\,
            in1 => \N__35302\,
            in2 => \_gnd_net_\,
            in3 => \N__34750\,
            lcout => \this_vga_signals.g1_0_0\,
            ltout => \this_vga_signals.g1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_36_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100010111"
        )
    port map (
            in0 => \N__34995\,
            in1 => \N__27956\,
            in2 => \N__26173\,
            in3 => \N__35153\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_22_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27431\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27027\,
            lcout => \this_vga_signals.if_N_6_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIP1DV3_7_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001000101101"
        )
    port map (
            in0 => \N__27991\,
            in1 => \N__30328\,
            in2 => \N__26164\,
            in3 => \N__35150\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_27_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_35_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000001001100"
        )
    port map (
            in0 => \N__35000\,
            in1 => \N__28423\,
            in2 => \N__26155\,
            in3 => \N__26152\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_33_N_4L6_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26146\,
            in3 => \N__28525\,
            lcout => \this_vga_signals.g0_33_N_4L6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_1_12_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__35783\,
            in1 => \N__36534\,
            in2 => \N__26143\,
            in3 => \N__27145\,
            lcout => \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNI9A3Q6_6_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__26367\,
            in1 => \N__37696\,
            in2 => \N__36571\,
            in3 => \N__28039\,
            lcout => \this_ppu.N_753_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIO37G1_7_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__29053\,
            in1 => \N__30936\,
            in2 => \N__43251\,
            in3 => \N__43415\,
            lcout => \N_1725_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIKQ691_7_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__43416\,
            in1 => \N__43232\,
            in2 => \_gnd_net_\,
            in3 => \N__29052\,
            lcout => \N_1717_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_o2_0_13_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35763\,
            in2 => \_gnd_net_\,
            in3 => \N__29190\,
            lcout => \this_ppu.N_1002_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_12_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__36535\,
            in1 => \N__26314\,
            in2 => \N__33171\,
            in3 => \N__27384\,
            lcout => \M_this_state_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_4_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26305\,
            lcout => \M_this_delay_clk_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNIR3631_1_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28168\,
            in1 => \N__26843\,
            in2 => \N__26890\,
            in3 => \N__43371\,
            lcout => \un1_M_this_oam_address_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_0_o2_0_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__26290\,
            in1 => \N__37427\,
            in2 => \N__26272\,
            in3 => \N__26254\,
            lcout => \this_ppu.N_767_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27588\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27675\,
            lcout => \this_start_data_delay_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42056\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_data_tmp_d_1_sqmuxa_i_0_o3_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__27587\,
            in1 => \N__27615\,
            in2 => \N__27681\,
            in3 => \N__28167\,
            lcout => \N_778_0\,
            ltout => \N_778_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI13IA1_0_1_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__26887\,
            in1 => \N__26844\,
            in2 => \N__26566\,
            in3 => \N__43228\,
            lcout => \N_1701_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_0_LC_17_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27464\,
            in1 => \N__26841\,
            in2 => \_gnd_net_\,
            in3 => \N__26789\,
            lcout => \M_this_oam_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42067\,
            ce => 'H',
            sr => \N__41641\
        );

    \M_this_oam_address_q_5_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__26497\,
            in1 => \N__27463\,
            in2 => \_gnd_net_\,
            in3 => \N__26527\,
            lcout => \M_this_oam_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42067\,
            ce => 'H',
            sr => \N__41641\
        );

    \M_this_oam_address_q_RNIRA651_4_LC_17_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26970\,
            in1 => \N__26426\,
            in2 => \N__26924\,
            in3 => \N__26397\,
            lcout => \un1_M_this_oam_address_q_c5\,
            ltout => \un1_M_this_oam_address_q_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_6_LC_17_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__26498\,
            in1 => \N__26447\,
            in2 => \N__26473\,
            in3 => \N__27466\,
            lcout => \M_this_oam_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42067\,
            ce => 'H',
            sr => \N__41641\
        );

    \M_this_oam_address_q_3_LC_17_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__27465\,
            in1 => \N__26427\,
            in2 => \N__26981\,
            in3 => \N__26398\,
            lcout => \M_this_oam_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42067\,
            ce => 'H',
            sr => \N__41641\
        );

    \M_this_oam_address_q_1_LC_17_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__26842\,
            in1 => \N__27482\,
            in2 => \N__26889\,
            in3 => \N__26796\,
            lcout => \M_this_oam_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42078\,
            ce => 'H',
            sr => \N__41639\
        );

    \M_this_oam_address_q_2_LC_17_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__26399\,
            in1 => \N__27480\,
            in2 => \_gnd_net_\,
            in3 => \N__26431\,
            lcout => \M_this_oam_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42078\,
            ce => 'H',
            sr => \N__41639\
        );

    \M_this_oam_address_q_4_LC_17_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__27481\,
            in1 => \N__26977\,
            in2 => \N__26925\,
            in3 => \N__26944\,
            lcout => \M_this_oam_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42078\,
            ce => 'H',
            sr => \N__41639\
        );

    \this_ppu.M_this_oam_ram_write_data_0_sqmuxa_0_a3_0_a2_LC_17_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__26875\,
            in1 => \N__26845\,
            in2 => \_gnd_net_\,
            in3 => \N__26790\,
            lcout => \M_this_oam_ram_write_data_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011011101"
        )
    port map (
            in0 => \N__29929\,
            in1 => \N__29876\,
            in2 => \_gnd_net_\,
            in3 => \N__29842\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1\,
            ltout => \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110001"
        )
    port map (
            in0 => \N__30535\,
            in1 => \N__27763\,
            in2 => \N__26572\,
            in3 => \N__29626\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_0_1\,
            ltout => \this_vga_signals.mult1_un47_sum_ac0_3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__28702\,
            in1 => \_gnd_net_\,
            in2 => \N__26569\,
            in3 => \N__34990\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28293\,
            lcout => \this_vga_signals.M_vcounter_q_9_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42003\,
            ce => \N__34246\,
            sr => \N__34214\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30762\,
            lcout => \this_vga_signals.M_vcounter_q_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42003\,
            ce => \N__34246\,
            sr => \N__34214\
        );

    \this_vga_signals.un5_vaddress_g0_3_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__34991\,
            in1 => \N__28703\,
            in2 => \N__27187\,
            in3 => \N__28748\,
            lcout => \this_vga_signals.g0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30725\,
            lcout => \this_vga_signals.M_vcounter_q_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42003\,
            ce => \N__34246\,
            sr => \N__34214\
        );

    \this_vga_signals.un5_vaddress_g0_5_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__34992\,
            in1 => \N__28704\,
            in2 => \_gnd_net_\,
            in3 => \N__28749\,
            lcout => \this_vga_signals.mult1_un54_sum_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_4_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27708\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42009\,
            ce => \N__34248\,
            sr => \N__34215\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_5_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34277\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42009\,
            ce => \N__34248\,
            sr => \N__34215\
        );

    \this_vga_signals.M_vcounter_q_esr_9_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28292\,
            lcout => \this_vga_signals_M_vcounter_q_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42009\,
            ce => \N__34248\,
            sr => \N__34215\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28325\,
            lcout => \this_vga_signals.M_vcounter_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42009\,
            ce => \N__34248\,
            sr => \N__34215\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001111011"
        )
    port map (
            in0 => \N__35408\,
            in1 => \N__35515\,
            in2 => \N__28986\,
            in3 => \N__35248\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__28584\,
            in1 => \N__28977\,
            in2 => \_gnd_net_\,
            in3 => \N__35409\,
            lcout => \this_vga_signals.mult1_un61_sum_axb2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_0_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__29764\,
            in1 => \N__29714\,
            in2 => \_gnd_net_\,
            in3 => \N__29620\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI0FP_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__29715\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28196\,
            lcout => \this_vga_signals.vaddress_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__27949\,
            in1 => \N__34881\,
            in2 => \_gnd_net_\,
            in3 => \N__27910\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_33_N_3L4_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010100001111"
        )
    port map (
            in0 => \N__28705\,
            in1 => \_gnd_net_\,
            in2 => \N__34943\,
            in3 => \N__28768\,
            lcout => \this_vga_signals.g0_33_N_3L4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_24_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__34967\,
            in1 => \N__28711\,
            in2 => \_gnd_net_\,
            in3 => \N__28766\,
            lcout => \this_vga_signals.mult1_un54_sum_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_19_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000101010"
        )
    port map (
            in0 => \N__28424\,
            in1 => \N__27838\,
            in2 => \N__34999\,
            in3 => \N__28383\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_17_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__34966\,
            in1 => \N__28712\,
            in2 => \_gnd_net_\,
            in3 => \N__28767\,
            lcout => \this_vga_signals.mult1_un54_sum_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_16_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111000110"
        )
    port map (
            in0 => \N__29536\,
            in1 => \N__30112\,
            in2 => \N__29497\,
            in3 => \N__29572\,
            lcout => \this_vga_signals.mult1_un47_sum_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_a3_1_12_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__29201\,
            in1 => \N__36533\,
            in2 => \_gnd_net_\,
            in3 => \N__29289\,
            lcout => \this_ppu.N_1115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_33_N_5L8_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011001100"
        )
    port map (
            in0 => \N__29803\,
            in1 => \N__28666\,
            in2 => \N__27139\,
            in3 => \N__27130\,
            lcout => \this_vga_signals.g0_33_N_5L8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27326\,
            in1 => \N__27028\,
            in2 => \N__27118\,
            in3 => \N__27117\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_21_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            clk => \N__42037\,
            ce => 'H',
            sr => \N__34219\
        );

    \this_vga_signals.M_vcounter_q_1_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27328\,
            in1 => \N__27432\,
            in2 => \_gnd_net_\,
            in3 => \N__27010\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            clk => \N__42037\,
            ce => 'H',
            sr => \N__34219\
        );

    \this_vga_signals.M_vcounter_q_2_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27327\,
            in1 => \N__28928\,
            in2 => \_gnd_net_\,
            in3 => \N__27007\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            clk => \N__42037\,
            ce => 'H',
            sr => \N__34219\
        );

    \this_vga_signals.M_vcounter_q_3_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27329\,
            in1 => \N__35464\,
            in2 => \_gnd_net_\,
            in3 => \N__27208\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            clk => \N__42037\,
            ce => 'H',
            sr => \N__34219\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35318\,
            in2 => \_gnd_net_\,
            in3 => \N__27205\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34947\,
            in2 => \_gnd_net_\,
            in3 => \N__27202\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34758\,
            in2 => \_gnd_net_\,
            in3 => \N__27199\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35151\,
            in2 => \_gnd_net_\,
            in3 => \N__27196\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30692\,
            in2 => \_gnd_net_\,
            in3 => \N__27193\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\,
            ltout => OPEN,
            carryin => \bfn_18_22_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30452\,
            in2 => \_gnd_net_\,
            in3 => \N__27190\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27426\,
            in2 => \_gnd_net_\,
            in3 => \N__28905\,
            lcout => \this_vga_signals.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.IO_port_data_write_0_a2_i_o2_2_1_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__27874\,
            in1 => \N__30895\,
            in2 => \N__29155\,
            in3 => \N__36430\,
            lcout => \this_vga_signals.IO_port_data_write_0_a2_i_o2_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__27427\,
            in1 => \N__35465\,
            in2 => \N__28929\,
            in3 => \N__35319\,
            lcout => \this_vga_signals.vsync_1_0_a3_0_a3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_13_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__29082\,
            in1 => \N__27385\,
            in2 => \N__36442\,
            in3 => \N__31059\,
            lcout => \M_this_state_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_data_count_qlde_i_0_o2_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__27871\,
            in1 => \N__29144\,
            in2 => \_gnd_net_\,
            in3 => \N__27382\,
            lcout => \N_816_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_1_18_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100011"
        )
    port map (
            in0 => \N__27616\,
            in1 => \N__43221\,
            in2 => \N__27682\,
            in3 => \N__27592\,
            lcout => \this_ppu.N_430_1_0\,
            ltout => \this_ppu.N_430_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_fast_13_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__29081\,
            in1 => \N__27383\,
            in2 => \N__27364\,
            in3 => \N__27361\,
            lcout => \M_this_state_q_fastZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42057\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_18_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__28163\,
            in1 => \N__29080\,
            in2 => \N__31075\,
            in3 => \N__27872\,
            lcout => \M_this_state_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42057\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_38_i_0_a2_3_0_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27360\,
            in2 => \_gnd_net_\,
            in3 => \N__28162\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_38_i_0_a2_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_38_i_0_a2_3_x1_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__38588\,
            in1 => \N__29041\,
            in2 => \N__27352\,
            in3 => \N__37394\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_38_i_0_a2_3_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_38_i_0_a2_3_ns_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27349\,
            in3 => \N__30805\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_38_i_0_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_38_i_0_o3_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__37426\,
            in1 => \N__27688\,
            in2 => \N__27691\,
            in3 => \N__36518\,
            lcout => \N_38_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_38_i_0_a2_0_4_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__30918\,
            in1 => \N__27883\,
            in2 => \N__36443\,
            in3 => \N__41060\,
            lcout => \this_vga_signals.N_38_i_0_a2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_o2_0_15_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__27586\,
            in1 => \N__27679\,
            in2 => \_gnd_net_\,
            in3 => \N__27614\,
            lcout => \this_ppu.N_787_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_o2_15_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__27680\,
            in1 => \N__27613\,
            in2 => \_gnd_net_\,
            in3 => \N__27585\,
            lcout => \N_765_0\,
            ltout => \N_765_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_this_data_count_q4_i_0_366_i_0_1_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101111"
        )
    port map (
            in0 => \N__41061\,
            in1 => \_gnd_net_\,
            in2 => \N__27565\,
            in3 => \N__43219\,
            lcout => \this_ppu.N_229_1_0\,
            ltout => \this_ppu.N_229_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_this_data_count_q4_i_0_366_i_0_i_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27553\,
            in3 => \N__29194\,
            lcout => \N_229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_data_count_d_5_sqmuxa_0_a3_i_o3_i_a2_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43372\,
            in2 => \_gnd_net_\,
            in3 => \N__29240\,
            lcout => \N_1423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNI99C6_5_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000111"
        )
    port map (
            in0 => \N__29705\,
            in1 => \N__29755\,
            in2 => \N__29644\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.SUM_2_i_i_1_0_3\,
            ltout => \this_vga_signals.SUM_2_i_i_1_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI3GK81_8_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110100100011"
        )
    port map (
            in0 => \N__35137\,
            in1 => \N__30420\,
            in2 => \N__27436\,
            in3 => \N__30685\,
            lcout => \this_vga_signals.N_39_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_x1_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101111111"
        )
    port map (
            in0 => \N__29703\,
            in1 => \N__29753\,
            in2 => \N__29643\,
            in3 => \N__27733\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_1_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28229\,
            in2 => \N__28216\,
            in3 => \N__28253\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_1\,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_x0_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__29704\,
            in1 => \_gnd_net_\,
            in2 => \N__27727\,
            in3 => \N__29754\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_1_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_ns_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29658\,
            in2 => \N__27724\,
            in3 => \N__27721\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_6_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28332\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42010\,
            ce => \N__34247\,
            sr => \N__34216\
        );

    \this_vga_signals.M_vcounter_q_esr_4_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27715\,
            lcout => \this_vga_signals_M_vcounter_q_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42020\,
            ce => \N__34250\,
            sr => \N__34217\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIFI5N_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__28195\,
            in1 => \N__35219\,
            in2 => \_gnd_net_\,
            in3 => \N__34705\,
            lcout => \this_vga_signals.vaddress_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34284\,
            lcout => \this_vga_signals.M_vcounter_q_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42020\,
            ce => \N__34250\,
            sr => \N__34217\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_1_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__28194\,
            in1 => \N__29716\,
            in2 => \_gnd_net_\,
            in3 => \N__28237\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_0_ns_1_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001000101000"
        )
    port map (
            in0 => \N__29872\,
            in1 => \N__29831\,
            in2 => \N__29930\,
            in3 => \N__29621\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un47_sum_ac0_3_0_0_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_0_ns_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111110101111"
        )
    port map (
            in0 => \N__29622\,
            in1 => \N__29765\,
            in2 => \N__27781\,
            in3 => \N__29717\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\,
            ltout => \this_vga_signals.mult1_un47_sum_ac0_3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010110000"
        )
    port map (
            in0 => \N__27778\,
            in1 => \N__27772\,
            in2 => \N__27766\,
            in3 => \N__27762\,
            lcout => \this_vga_signals.mult1_un47_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m5_s_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001100000"
        )
    port map (
            in0 => \N__28937\,
            in1 => \N__35518\,
            in2 => \N__29008\,
            in3 => \N__28981\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m5_s_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m5_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__28856\,
            in1 => \N__28650\,
            in2 => \N__27751\,
            in3 => \N__27742\,
            lcout => \this_vga_signals.mult1_un68_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_21_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100110010000"
        )
    port map (
            in0 => \N__34735\,
            in1 => \N__34162\,
            in2 => \N__29988\,
            in3 => \N__34141\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_0_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001100000"
        )
    port map (
            in0 => \N__35516\,
            in1 => \N__28935\,
            in2 => \N__27748\,
            in3 => \N__29002\,
            lcout => \this_vga_signals.N_2840_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_ns_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35553\,
            in2 => \N__28435\,
            in3 => \N__28597\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m5_d_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110011000101"
        )
    port map (
            in0 => \N__35517\,
            in1 => \N__28936\,
            in2 => \N__27745\,
            in3 => \N__29003\,
            lcout => \this_vga_signals.if_m5_d\,
            ltout => \this_vga_signals.if_m5_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_18_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__28651\,
            in1 => \N__28855\,
            in2 => \N__27736\,
            in3 => \N__27844\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_1_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__27909\,
            in1 => \N__35684\,
            in2 => \_gnd_net_\,
            in3 => \N__27945\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIS9T25_0_9_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101001"
        )
    port map (
            in0 => \N__28030\,
            in1 => \N__27914\,
            in2 => \N__27990\,
            in3 => \N__28785\,
            lcout => \this_vga_signals.N_27_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_0_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__27787\,
            in1 => \N__28425\,
            in2 => \_gnd_net_\,
            in3 => \N__28516\,
            lcout => \this_vga_signals.g0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNICUI21_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100110011001"
        )
    port map (
            in0 => \N__34716\,
            in1 => \N__35146\,
            in2 => \N__35300\,
            in3 => \N__28201\,
            lcout => \this_vga_signals.vaddress_7\,
            ltout => \this_vga_signals.vaddress_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIS9T25_9_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001001011"
        )
    port map (
            in0 => \N__28784\,
            in1 => \N__27982\,
            in2 => \N__27832\,
            in3 => \N__28029\,
            lcout => \this_vga_signals.N_27_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_N_3_i_LC_19_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28456\,
            in1 => \N__27829\,
            in2 => \N__27816\,
            in3 => \N__28858\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_9_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011100101000"
        )
    port map (
            in0 => \N__28603\,
            in1 => \N__28792\,
            in2 => \N__27799\,
            in3 => \N__28828\,
            lcout => \this_vga_signals.if_m6_i_x2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIA65T2_9_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000001"
        )
    port map (
            in0 => \N__30429\,
            in1 => \N__28359\,
            in2 => \N__28031\,
            in3 => \_gnd_net_\,
            lcout => \N_842_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_3_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111010100110"
        )
    port map (
            in0 => \N__27964\,
            in1 => \N__27915\,
            in2 => \N__35013\,
            in3 => \N__27958\,
            lcout => \this_vga_signals.g1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_32_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35460\,
            in2 => \_gnd_net_\,
            in3 => \N__28909\,
            lcout => \this_vga_signals.g0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI65531_6_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001001"
        )
    port map (
            in0 => \N__30540\,
            in1 => \N__30670\,
            in2 => \N__35155\,
            in3 => \N__34745\,
            lcout => \this_vga_signals.vaddress_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_1_9_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__30571\,
            in1 => \N__30428\,
            in2 => \_gnd_net_\,
            in3 => \N__30539\,
            lcout => \this_vga_signals_CO0_0_i_i\,
            ltout => \this_vga_signals_CO0_0_i_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIGBA04_9_LC_19_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28786\,
            in2 => \N__27994\,
            in3 => \N__27989\,
            lcout => \this_vga_signals.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_3_LC_19_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__35286\,
            in1 => \N__27957\,
            in2 => \N__27919\,
            in3 => \N__34746\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_38_i_0_a2_0_4_1_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30833\,
            in2 => \_gnd_net_\,
            in3 => \N__28164\,
            lcout => \this_vga_signals.N_38_i_0_a2_0_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_1_17_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101110011"
        )
    port map (
            in0 => \N__29222\,
            in1 => \N__27873\,
            in2 => \N__29206\,
            in3 => \N__43355\,
            lcout => OPEN,
            ltout => \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_17_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000001100"
        )
    port map (
            in0 => \N__43356\,
            in1 => \N__29062\,
            in2 => \N__27877\,
            in3 => \N__28166\,
            lcout => \M_this_state_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42068\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIQ6821_8_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__30693\,
            in1 => \N__30457\,
            in2 => \_gnd_net_\,
            in3 => \N__35152\,
            lcout => \this_vga_signals.vsync_1_0_a3_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_1_7_5__m12_0_a3_0_a3_0_o2_LC_19_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__29221\,
            in1 => \N__36099\,
            in2 => \_gnd_net_\,
            in3 => \N__29271\,
            lcout => \N_773_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_a3_4_LC_19_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31034\,
            in2 => \_gnd_net_\,
            in3 => \N__38587\,
            lcout => \this_ppu.N_1162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_this_state_q_8_0_i_0_0_i_LC_19_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__28165\,
            in1 => \N__43354\,
            in2 => \N__36532\,
            in3 => \N__30836\,
            lcout => \N_247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_7_LC_19_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__30296\,
            in1 => \N__31054\,
            in2 => \N__29116\,
            in3 => \N__29046\,
            lcout => \M_this_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_8_LC_19_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__30297\,
            in1 => \N__31055\,
            in2 => \N__29101\,
            in3 => \N__30928\,
            lcout => \M_this_state_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_address_q_0_i_0_o2_1_LC_19_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__43365\,
            in1 => \N__36354\,
            in2 => \_gnd_net_\,
            in3 => \N__38586\,
            lcout => \N_794_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_address_d_4_sqmuxa_0_a3_i_o3_i_a3_0_LC_19_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43234\,
            in2 => \_gnd_net_\,
            in3 => \N__36113\,
            lcout => \this_ppu_M_this_map_address_d_4_sqmuxa_0_a3_i_o3_i_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_data_1_0_a2_3_LC_19_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__36513\,
            in1 => \N__43401\,
            in2 => \_gnd_net_\,
            in3 => \N__36444\,
            lcout => \this_ppu.N_1322\,
            ltout => \this_ppu.N_1322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_data_1_0_i_0_LC_19_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__42444\,
            in1 => \N__40751\,
            in2 => \N__28129\,
            in3 => \N__36514\,
            lcout => \M_this_spr_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI65531_0_6_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__30684\,
            in1 => \N__34704\,
            in2 => \N__35154\,
            in3 => \N__30502\,
            lcout => \this_vga_signals.N_1247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_0_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28270\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28231\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0\,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_2_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__30683\,
            in1 => \N__34703\,
            in2 => \N__28336\,
            in3 => \N__30501\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_6_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28333\,
            lcout => \this_vga_signals_M_vcounter_q_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42021\,
            ce => \N__34249\,
            sr => \N__34218\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_9_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28300\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42021\,
            ce => \N__34249\,
            sr => \N__34218\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_1_1_1_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100010000111"
        )
    port map (
            in0 => \N__28269\,
            in1 => \N__28230\,
            in2 => \N__28260\,
            in3 => \N__28215\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_0_1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_7_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30766\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42021\,
            ce => \N__34249\,
            sr => \N__34218\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_8_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30730\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42021\,
            ce => \N__34249\,
            sr => \N__34218\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010000111"
        )
    port map (
            in0 => \N__28693\,
            in1 => \N__28769\,
            in2 => \N__35293\,
            in3 => \N__28200\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1\,
            ltout => \this_vga_signals.mult1_un54_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011011001111"
        )
    port map (
            in0 => \N__34971\,
            in1 => \N__35240\,
            in2 => \N__28171\,
            in3 => \N__34123\,
            lcout => \this_vga_signals.mult1_un54_sum_c2_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_10_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101111010100"
        )
    port map (
            in0 => \N__34039\,
            in1 => \N__28444\,
            in2 => \N__28459\,
            in3 => \N__30037\,
            lcout => \this_vga_signals.g0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35602\,
            in2 => \_gnd_net_\,
            in3 => \N__34070\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_29_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101011010"
        )
    port map (
            in0 => \N__30073\,
            in1 => \N__29488\,
            in2 => \N__28447\,
            in3 => \N__29531\,
            lcout => \this_vga_signals.mult1_un47_sum_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110100101"
        )
    port map (
            in0 => \N__35663\,
            in1 => \N__35603\,
            in2 => \N__35705\,
            in3 => \N__34071\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc1\,
            ltout => \this_vga_signals.mult1_un47_sum_axbxc1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x1_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001010"
        )
    port map (
            in0 => \N__35241\,
            in1 => \N__34972\,
            in2 => \N__28438\,
            in3 => \N__34131\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_1_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__34132\,
            in1 => \N__30028\,
            in2 => \_gnd_net_\,
            in3 => \N__29987\,
            lcout => \this_vga_signals.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010111101"
        )
    port map (
            in0 => \N__30017\,
            in1 => \N__29982\,
            in2 => \N__34137\,
            in3 => \N__35384\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__35317\,
            in1 => \_gnd_net_\,
            in2 => \N__35405\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000100010"
        )
    port map (
            in0 => \N__28426\,
            in1 => \N__28387\,
            in2 => \N__34946\,
            in3 => \N__28369\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x0_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101100110011"
        )
    port map (
            in0 => \N__35315\,
            in1 => \N__30016\,
            in2 => \N__34944\,
            in3 => \N__34125\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_3_1_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100000011110"
        )
    port map (
            in0 => \N__34130\,
            in1 => \N__29983\,
            in2 => \N__28947\,
            in3 => \N__35566\,
            lcout => \this_vga_signals.g0_0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m3_i_m2_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000111100"
        )
    port map (
            in0 => \N__35316\,
            in1 => \N__34152\,
            in2 => \N__34945\,
            in3 => \N__34126\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m3_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__35514\,
            in1 => \N__35552\,
            in2 => \N__28591\,
            in3 => \N__35380\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_d\,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__28588\,
            in1 => \N__28539\,
            in2 => \N__28564\,
            in3 => \N__30079\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_15_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011001100011"
        )
    port map (
            in0 => \N__30031\,
            in1 => \N__35400\,
            in2 => \N__28561\,
            in3 => \N__29989\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__28549\,
            in1 => \N__28540\,
            in2 => \N__28528\,
            in3 => \N__28517\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30196\,
            in1 => \N__29014\,
            in2 => \N__28492\,
            in3 => \N__28489\,
            lcout => \this_vga_signals.N_3_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35399\,
            in1 => \N__28648\,
            in2 => \N__28474\,
            in3 => \N__28982\,
            lcout => \this_vga_signals.g0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_0_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__29007\,
            in1 => \_gnd_net_\,
            in2 => \N__28987\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_c2_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010001110001"
        )
    port map (
            in0 => \N__28948\,
            in1 => \N__28649\,
            in2 => \N__35521\,
            in3 => \N__28857\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_3_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35323\,
            in1 => \N__35401\,
            in2 => \N__28837\,
            in3 => \N__28834\,
            lcout => \this_vga_signals.g0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111100000000"
        )
    port map (
            in0 => \N__35410\,
            in1 => \N__28822\,
            in2 => \N__28813\,
            in3 => \N__28798\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_31_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28713\,
            in2 => \_gnd_net_\,
            in3 => \N__28770\,
            lcout => \this_vga_signals.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_9_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__30455\,
            in1 => \N__30567\,
            in2 => \_gnd_net_\,
            in3 => \N__30533\,
            lcout => \this_vga_signals.vaddress_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_x2_1_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__28771\,
            in1 => \_gnd_net_\,
            in2 => \N__28717\,
            in3 => \N__34986\,
            lcout => \this_vga_signals.N_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111101101111"
        )
    port map (
            in0 => \N__35489\,
            in1 => \N__28665\,
            in2 => \N__28618\,
            in3 => \N__30211\,
            lcout => \this_vga_signals.if_m5_i_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_1_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110010011"
        )
    port map (
            in0 => \N__35322\,
            in1 => \N__35099\,
            in2 => \N__35005\,
            in3 => \N__34747\,
            lcout => \this_vga_signals.g1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_0_a3_1_2_1_0_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__30929\,
            in1 => \N__30887\,
            in2 => \_gnd_net_\,
            in3 => \N__43224\,
            lcout => \this_ppu.M_this_state_q_srsts_0_0_a3_1_2_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_16_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__29143\,
            in1 => \N__29089\,
            in2 => \N__31090\,
            in3 => \N__30838\,
            lcout => \M_this_state_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_2_15_LC_20_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__43225\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35784\,
            lcout => \this_ppu.N_235_2_0\,
            ltout => \this_ppu.N_235_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_0_15_LC_20_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__29142\,
            in1 => \N__43471\,
            in2 => \N__29056\,
            in3 => \N__30837\,
            lcout => \this_ppu.M_this_state_q_srsts_i_i_0_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_1_LC_20_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__40862\,
            in1 => \N__31067\,
            in2 => \N__29449\,
            in3 => \N__30969\,
            lcout => \M_this_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_10_LC_20_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__31137\,
            in1 => \N__31065\,
            in2 => \N__36114\,
            in3 => \N__33015\,
            lcout => \M_this_state_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_1_7_5__m17_0_a3_0_a3_0_o2_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__40861\,
            in1 => \N__29042\,
            in2 => \_gnd_net_\,
            in3 => \N__37386\,
            lcout => \N_815_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_4_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__29020\,
            in1 => \N__36160\,
            in2 => \N__32866\,
            in3 => \N__30793\,
            lcout => \M_this_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_9_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__31068\,
            in1 => \N__31138\,
            in2 => \N__33022\,
            in3 => \N__29281\,
            lcout => \M_this_state_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_11_LC_20_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__29107\,
            in1 => \N__30792\,
            in2 => \N__29244\,
            in3 => \N__31066\,
            lcout => \M_this_state_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_15_LC_20_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000011001100"
        )
    port map (
            in0 => \N__29205\,
            in1 => \N__29161\,
            in2 => \N__29151\,
            in3 => \N__37455\,
            lcout => \M_this_state_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_7_LC_20_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__36154\,
            in1 => \N__36298\,
            in2 => \_gnd_net_\,
            in3 => \N__35846\,
            lcout => \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_0_a2_0_0_LC_20_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__42616\,
            in1 => \N__35777\,
            in2 => \N__29445\,
            in3 => \N__43235\,
            lcout => \this_ppu.N_1425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_11_LC_20_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__32927\,
            in1 => \N__33013\,
            in2 => \_gnd_net_\,
            in3 => \N__33088\,
            lcout => \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_8_LC_20_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__36155\,
            in1 => \N__36299\,
            in2 => \_gnd_net_\,
            in3 => \N__35847\,
            lcout => \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_o2_6_LC_20_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__33089\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32928\,
            lcout => \this_ppu.N_807_0\,
            ltout => \this_ppu.N_807_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_this_state_q_11_0_0_m3_LC_20_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__36300\,
            in1 => \N__33014\,
            in2 => \N__29092\,
            in3 => \N__36242\,
            lcout => \this_ppu.N_969\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_2_LC_20_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__32981\,
            in1 => \N__33091\,
            in2 => \_gnd_net_\,
            in3 => \N__32935\,
            lcout => \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_a2_0_1_LC_20_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32934\,
            in1 => \N__32980\,
            in2 => \N__36210\,
            in3 => \N__33090\,
            lcout => \this_ppu.N_1341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_data_1_0_i_2_LC_20_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__42773\,
            in1 => \N__35976\,
            in2 => \N__40436\,
            in3 => \N__36531\,
            lcout => \M_this_spr_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_5_LC_21_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29341\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42011\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_20_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010000101011"
        )
    port map (
            in0 => \N__30030\,
            in1 => \N__29980\,
            in2 => \N__29299\,
            in3 => \N__35407\,
            lcout => \this_vga_signals.mult1_un54_sum_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_a3_0_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35320\,
            in2 => \_gnd_net_\,
            in3 => \N__35548\,
            lcout => \this_vga_signals.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_11_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100110100110"
        )
    port map (
            in0 => \N__30108\,
            in1 => \N__29527\,
            in2 => \N__29490\,
            in3 => \N__29571\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un47_sum_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_8_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001100110000"
        )
    port map (
            in0 => \N__34186\,
            in1 => \N__34174\,
            in2 => \N__29308\,
            in3 => \N__29305\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_23_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101110110100"
        )
    port map (
            in0 => \N__29480\,
            in1 => \N__29523\,
            in2 => \N__29776\,
            in3 => \N__29569\,
            lcout => \this_vga_signals.mult1_un47_sum_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_28_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010110011010"
        )
    port map (
            in0 => \N__29570\,
            in1 => \N__29481\,
            in2 => \N__29532\,
            in3 => \N__30107\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un47_sum_3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_38_LC_21_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010000101011"
        )
    port map (
            in0 => \N__30029\,
            in1 => \N__29981\,
            in2 => \N__29806\,
            in3 => \N__35406\,
            lcout => \this_vga_signals.mult1_un54_sum_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_3_0_LC_21_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__29880\,
            in1 => \N__29843\,
            in2 => \N__29937\,
            in3 => \N__29642\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_0_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m18_i_o2_0_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100001"
        )
    port map (
            in0 => \N__30688\,
            in1 => \N__34706\,
            in2 => \N__35136\,
            in3 => \N__30520\,
            lcout => \this_ppu.m18_i_o2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_25_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__34069\,
            in1 => \_gnd_net_\,
            in2 => \N__35616\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_5_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29767\,
            in2 => \_gnd_net_\,
            in3 => \N__29719\,
            lcout => \N_814_0\,
            ltout => \N_814_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_1_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__29665\,
            in1 => \N__29659\,
            in2 => \N__29647\,
            in3 => \N__29635\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un47_sum_axbxc3_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_2_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001110000"
        )
    port map (
            in0 => \N__35100\,
            in1 => \N__30421\,
            in2 => \N__29578\,
            in3 => \N__30669\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_2_2\,
            ltout => \this_vga_signals.mult1_un47_sum_axbxc3_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_21_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29476\,
            in2 => \N__29575\,
            in3 => \N__29557\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_21_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100110100110"
        )
    port map (
            in0 => \N__29558\,
            in1 => \N__29522\,
            in2 => \N__29489\,
            in3 => \N__34068\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un47_sum_axbxc3_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_21_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35604\,
            in1 => \_gnd_net_\,
            in2 => \N__30133\,
            in3 => \N__30130\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000111110101"
        )
    port map (
            in0 => \N__35656\,
            in1 => \N__35609\,
            in2 => \N__35713\,
            in3 => \N__34072\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un47_sum_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_21_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__30124\,
            in1 => \N__30103\,
            in2 => \N__30085\,
            in3 => \N__34118\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1\,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_21_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010000101101"
        )
    port map (
            in0 => \N__34119\,
            in1 => \N__30018\,
            in2 => \N__30082\,
            in3 => \N__29978\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_1_LC_21_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30072\,
            in1 => \N__34880\,
            in2 => \N__30052\,
            in3 => \N__35386\,
            lcout => \this_vga_signals.g0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_x2_2_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100110011010"
        )
    port map (
            in0 => \N__35385\,
            in1 => \N__30019\,
            in2 => \N__34136\,
            in3 => \N__29979\,
            lcout => \this_vga_signals.N_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_4_LC_21_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001110011"
        )
    port map (
            in0 => \N__29851\,
            in1 => \N__29938\,
            in2 => \N__29902\,
            in3 => \N__29887\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_3_LC_21_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__29886\,
            in1 => \N__29850\,
            in2 => \N__30186\,
            in3 => \N__30156\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_3\,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb1_LC_21_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001011111"
        )
    port map (
            in0 => \N__35608\,
            in1 => \_gnd_net_\,
            in2 => \N__30280\,
            in3 => \N__35709\,
            lcout => \this_vga_signals.mult1_un47_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIPMQM_6_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__35089\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34748\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_8_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101010000"
        )
    port map (
            in0 => \N__30534\,
            in1 => \N__30459\,
            in2 => \N__30277\,
            in3 => \N__30651\,
            lcout => \this_vga_signals.N_5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI3GK81_0_8_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011011011"
        )
    port map (
            in0 => \N__30652\,
            in1 => \N__30274\,
            in2 => \N__35133\,
            in3 => \N__30458\,
            lcout => \this_vga_signals.N_39_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_26_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100011100111"
        )
    port map (
            in0 => \N__30240\,
            in1 => \N__34879\,
            in2 => \N__34633\,
            in3 => \N__30259\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_LC_21_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111111111"
        )
    port map (
            in0 => \N__30250\,
            in1 => \N__30241\,
            in2 => \N__30229\,
            in3 => \N__35304\,
            lcout => OPEN,
            ltout => \this_vga_signals.g3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_13_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__30226\,
            in1 => \N__35329\,
            in2 => \N__30220\,
            in3 => \N__30217\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__35305\,
            in1 => \N__35398\,
            in2 => \N__35520\,
            in3 => \N__30205\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_1_0_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011111111"
        )
    port map (
            in0 => \N__30638\,
            in1 => \N__30187\,
            in2 => \N__35135\,
            in3 => \N__30157\,
            lcout => \this_vga_signals.g2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_7_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30755\,
            lcout => \this_vga_signals_M_vcounter_q_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42070\,
            ce => \N__34252\,
            sr => \N__34221\
        );

    \this_vga_signals.M_vcounter_q_esr_8_LC_21_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30726\,
            lcout => \this_vga_signals_M_vcounter_q_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42070\,
            ce => \N__34252\,
            sr => \N__34221\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIN3821_6_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__35075\,
            in1 => \N__30637\,
            in2 => \_gnd_net_\,
            in3 => \N__34744\,
            lcout => \N_1001_0\,
            ltout => \N_1001_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_0_9_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30532\,
            in2 => \N__30475\,
            in3 => \N__30456\,
            lcout => \this_vga_signals.g4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_o2_3_15_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30835\,
            in2 => \_gnd_net_\,
            in3 => \N__36100\,
            lcout => \this_ppu.N_856_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_a2_3_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__36000\,
            in1 => \N__36307\,
            in2 => \N__36250\,
            in3 => \N__35840\,
            lcout => \this_ppu.N_1278\,
            ltout => \this_ppu.N_1278_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_3_LC_21_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__31129\,
            in1 => \N__31089\,
            in2 => \N__30319\,
            in3 => \N__36343\,
            lcout => \M_this_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_0_a3_0_LC_21_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__36001\,
            in1 => \N__36306\,
            in2 => \N__31123\,
            in3 => \N__30315\,
            lcout => OPEN,
            ltout => \this_ppu.N_1149_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_0_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001010"
        )
    port map (
            in0 => \N__30316\,
            in1 => \N__30301\,
            in2 => \N__30283\,
            in3 => \N__30943\,
            lcout => led_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_0_0_tz_0_LC_21_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100010101"
        )
    port map (
            in0 => \N__31088\,
            in1 => \N__35793\,
            in2 => \N__30955\,
            in3 => \N__35841\,
            lcout => \this_ppu.M_this_state_q_srsts_0_0_0_tz_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_1_7_5__m17_0_a3_0_a3_0_a3_LC_21_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000000"
        )
    port map (
            in0 => \N__30937\,
            in1 => \N__30888\,
            in2 => \N__35797\,
            in3 => \_gnd_net_\,
            lcout => led_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_6_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__30791\,
            in1 => \N__33020\,
            in2 => \N__30847\,
            in3 => \N__30775\,
            lcout => \M_this_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42091\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_0_sqmuxa_i_i_o3_0_a2_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30834\,
            in2 => \_gnd_net_\,
            in3 => \N__38275\,
            lcout => \N_1415\,
            ltout => \N_1415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_0_sqmuxa_i_i_o3_0_o3_LC_21_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30796\,
            in3 => \N__43460\,
            lcout => \N_296_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_5_LC_21_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__31064\,
            in1 => \N__30790\,
            in2 => \N__30994\,
            in3 => \N__37387\,
            lcout => \M_this_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42091\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_a3_6_LC_21_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__38276\,
            in1 => \N__31063\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.N_1166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_a2_1_LC_21_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__34486\,
            in1 => \N__43756\,
            in2 => \N__36287\,
            in3 => \N__35839\,
            lcout => \this_ppu.N_1263\,
            ltout => \this_ppu.N_1263_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_a3_0_1_10_LC_21_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__33052\,
            in1 => \N__36243\,
            in2 => \N__30769\,
            in3 => \N__32932\,
            lcout => \this_ppu.N_1176_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_a3_0_0_3_LC_21_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33021\,
            in1 => \N__33051\,
            in2 => \N__32942\,
            in3 => \N__36153\,
            lcout => \this_ppu.M_this_state_q_srsts_0_i_a3_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_0_m2_0_LC_21_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110000010"
        )
    port map (
            in0 => \N__33019\,
            in1 => \N__36226\,
            in2 => \N__33087\,
            in3 => \N__32933\,
            lcout => \this_ppu.N_893\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_this_state_q_11_0_0_LC_21_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__42615\,
            in1 => \N__31096\,
            in2 => \N__31111\,
            in3 => \N__35773\,
            lcout => OPEN,
            ltout => \un1_M_this_state_q_11_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_substate_q_LC_21_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__32856\,
            in1 => \N__36156\,
            in2 => \N__31102\,
            in3 => \N__36124\,
            lcout => \M_this_substate_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42100\,
            ce => 'H',
            sr => \N__43106\
        );

    \this_ppu.un1_M_this_state_q_11_0_0_0_LC_21_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000000"
        )
    port map (
            in0 => \N__32988\,
            in1 => \N__33074\,
            in2 => \N__32947\,
            in3 => \N__35845\,
            lcout => OPEN,
            ltout => \this_ppu.un1_M_this_state_q_11_0_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_this_state_q_11_0_0_1_LC_21_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__33075\,
            in1 => \N__32989\,
            in2 => \N__31099\,
            in3 => \N__36196\,
            lcout => \this_ppu.un1_M_this_state_q_11_0_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_a3_2_LC_21_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37781\,
            in2 => \_gnd_net_\,
            in3 => \N__31079\,
            lcout => OPEN,
            ltout => \this_ppu.N_1158_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_2_LC_21_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__36195\,
            in1 => \N__30990\,
            in2 => \N__30973\,
            in3 => \N__30970\,
            lcout => \M_this_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_substate_d_0_sqmuxa_3_0_a3_0_a2_LC_21_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000001"
        )
    port map (
            in0 => \N__33073\,
            in1 => \N__32987\,
            in2 => \N__32943\,
            in3 => \_gnd_net_\,
            lcout => \N_1422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_spr_address_q_0_LC_22_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33210\,
            in1 => \N__32661\,
            in2 => \N__36379\,
            in3 => \N__36378\,
            lcout => \M_this_spr_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_22_14_0_\,
            carryout => \un1_M_this_spr_address_q_cry_0\,
            clk => \N__42012\,
            ce => 'H',
            sr => \N__41653\
        );

    \M_this_spr_address_q_1_LC_22_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33214\,
            in1 => \N__32441\,
            in2 => \_gnd_net_\,
            in3 => \N__32398\,
            lcout => \M_this_spr_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_0\,
            carryout => \un1_M_this_spr_address_q_cry_1\,
            clk => \N__42012\,
            ce => 'H',
            sr => \N__41653\
        );

    \M_this_spr_address_q_2_LC_22_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33211\,
            in1 => \N__32211\,
            in2 => \_gnd_net_\,
            in3 => \N__32191\,
            lcout => \M_this_spr_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_1\,
            carryout => \un1_M_this_spr_address_q_cry_2\,
            clk => \N__42012\,
            ce => 'H',
            sr => \N__41653\
        );

    \M_this_spr_address_q_3_LC_22_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33215\,
            in1 => \N__31998\,
            in2 => \_gnd_net_\,
            in3 => \N__31975\,
            lcout => \M_this_spr_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_2\,
            carryout => \un1_M_this_spr_address_q_cry_3\,
            clk => \N__42012\,
            ce => 'H',
            sr => \N__41653\
        );

    \M_this_spr_address_q_4_LC_22_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33212\,
            in1 => \N__31779\,
            in2 => \_gnd_net_\,
            in3 => \N__31759\,
            lcout => \M_this_spr_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_3\,
            carryout => \un1_M_this_spr_address_q_cry_4\,
            clk => \N__42012\,
            ce => 'H',
            sr => \N__41653\
        );

    \M_this_spr_address_q_5_LC_22_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33216\,
            in1 => \N__31581\,
            in2 => \_gnd_net_\,
            in3 => \N__31549\,
            lcout => \M_this_spr_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_4\,
            carryout => \un1_M_this_spr_address_q_cry_5\,
            clk => \N__42012\,
            ce => 'H',
            sr => \N__41653\
        );

    \M_this_spr_address_q_6_LC_22_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33213\,
            in1 => \N__31371\,
            in2 => \_gnd_net_\,
            in3 => \N__31351\,
            lcout => \M_this_spr_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_5\,
            carryout => \un1_M_this_spr_address_q_cry_6\,
            clk => \N__42012\,
            ce => 'H',
            sr => \N__41653\
        );

    \M_this_spr_address_q_7_LC_22_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33217\,
            in1 => \N__31159\,
            in2 => \_gnd_net_\,
            in3 => \N__31141\,
            lcout => \M_this_spr_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_6\,
            carryout => \un1_M_this_spr_address_q_cry_7\,
            clk => \N__42012\,
            ce => 'H',
            sr => \N__41653\
        );

    \M_this_spr_address_q_8_LC_22_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33206\,
            in1 => \N__33700\,
            in2 => \_gnd_net_\,
            in3 => \N__33682\,
            lcout => \M_this_spr_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_22_15_0_\,
            carryout => \un1_M_this_spr_address_q_cry_8\,
            clk => \N__42022\,
            ce => 'H',
            sr => \N__41652\
        );

    \M_this_spr_address_q_9_LC_22_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33209\,
            in1 => \N__33482\,
            in2 => \_gnd_net_\,
            in3 => \N__33457\,
            lcout => \M_this_spr_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_8\,
            carryout => \un1_M_this_spr_address_q_cry_9\,
            clk => \N__42022\,
            ce => 'H',
            sr => \N__41652\
        );

    \M_this_spr_address_q_10_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33204\,
            in1 => \N__33264\,
            in2 => \_gnd_net_\,
            in3 => \N__33226\,
            lcout => \M_this_spr_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_9\,
            carryout => \un1_M_this_spr_address_q_cry_10\,
            clk => \N__42022\,
            ce => 'H',
            sr => \N__41652\
        );

    \M_this_spr_address_q_11_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33208\,
            in1 => \N__38846\,
            in2 => \_gnd_net_\,
            in3 => \N__33223\,
            lcout => \M_this_spr_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_10\,
            carryout => \un1_M_this_spr_address_q_cry_11\,
            clk => \N__42022\,
            ce => 'H',
            sr => \N__41652\
        );

    \M_this_spr_address_q_12_LC_22_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33205\,
            in1 => \N__38902\,
            in2 => \_gnd_net_\,
            in3 => \N__33220\,
            lcout => \M_this_spr_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_11\,
            carryout => \un1_M_this_spr_address_q_cry_12\,
            clk => \N__42022\,
            ce => 'H',
            sr => \N__41652\
        );

    \M_this_spr_address_q_13_LC_22_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__38755\,
            in1 => \N__33207\,
            in2 => \_gnd_net_\,
            in3 => \N__33118\,
            lcout => \M_this_spr_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42022\,
            ce => 'H',
            sr => \N__41652\
        );

    \this_spr_ram.mem_radreg_11_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33115\,
            in1 => \N__43935\,
            in2 => \_gnd_net_\,
            in3 => \N__38205\,
            lcout => \this_spr_ram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42028\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_12_LC_22_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34027\,
            in1 => \N__41602\,
            in2 => \_gnd_net_\,
            in3 => \N__38206\,
            lcout => \this_spr_ram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42028\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_6_LC_22_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33109\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42038\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_22_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39107\,
            in1 => \N__34021\,
            in2 => \_gnd_net_\,
            in3 => \N__34006\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_mem_0_1_RNIM6VFZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_22_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__37027\,
            in1 => \N__36978\,
            in2 => \N__33988\,
            in3 => \N__36628\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_22_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__36979\,
            in1 => \N__37861\,
            in2 => \N__33985\,
            in3 => \N__36754\,
            lcout => \M_this_spr_ram_read_data_2\,
            ltout => \M_this_spr_ram_read_data_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNITTE65_5_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__34476\,
            in1 => \N__37122\,
            in2 => \N__33982\,
            in3 => \N__34437\,
            lcout => \M_this_ppu_vram_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39106\,
            in1 => \N__33964\,
            in2 => \_gnd_net_\,
            in3 => \N__33949\,
            lcout => \this_spr_ram.mem_mem_1_0_RNIMA1GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39121\,
            in1 => \N__33931\,
            in2 => \_gnd_net_\,
            in3 => \N__33919\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__39019\,
            in1 => \N__36995\,
            in2 => \N__33898\,
            in3 => \N__37038\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_22_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__36999\,
            in1 => \N__36790\,
            in2 => \N__33895\,
            in3 => \N__36013\,
            lcout => \M_this_spr_ram_read_data_1\,
            ltout => \M_this_spr_ram_read_data_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.vram_en_iv_i_0_o2_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36945\,
            in1 => \N__34384\,
            in2 => \N__34378\,
            in3 => \N__34296\,
            lcout => \this_ppu.N_1000_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_RNIB2R65_4_LC_22_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__34477\,
            in1 => \N__34430\,
            in2 => \N__37345\,
            in3 => \N__34336\,
            lcout => \M_this_ppu_vram_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_22_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001100100011"
        )
    port map (
            in0 => \N__36826\,
            in1 => \N__36712\,
            in2 => \N__37003\,
            in3 => \N__34312\,
            lcout => \M_this_spr_ram_read_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_5_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34285\,
            lcout => \this_vga_signals_M_vcounter_q_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42058\,
            ce => \N__34251\,
            sr => \N__34220\
        );

    \this_vga_signals.un5_vaddress_g0_3_2_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34842\,
            in2 => \_gnd_net_\,
            in3 => \N__35306\,
            lcout => \this_vga_signals.N_5_i_0\,
            ltout => \this_vga_signals.N_5_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_12_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010000111"
        )
    port map (
            in0 => \N__34074\,
            in1 => \N__35610\,
            in2 => \N__34177\,
            in3 => \N__35710\,
            lcout => \this_vga_signals.mult1_un47_sum_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_21_1_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011111010"
        )
    port map (
            in0 => \N__35314\,
            in1 => \N__35611\,
            in2 => \N__34938\,
            in3 => \N__34073\,
            lcout => \this_vga_signals.g0_21_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_40_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000111100"
        )
    port map (
            in0 => \N__35307\,
            in1 => \N__34153\,
            in2 => \N__34897\,
            in3 => \N__34124\,
            lcout => \this_vga_signals.if_N_7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_30_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__34075\,
            in1 => \N__35712\,
            in2 => \N__35617\,
            in3 => \N__35665\,
            lcout => \this_vga_signals.mult1_un47_sum_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_43_LC_22_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010011001"
        )
    port map (
            in0 => \N__35711\,
            in1 => \N__35664\,
            in2 => \N__35629\,
            in3 => \N__35615\,
            lcout => \this_vga_signals.mult1_un47_sum_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_45_LC_22_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__35557\,
            in1 => \N__35527\,
            in2 => \N__35519\,
            in3 => \N__35392\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_d_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_6_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010010011"
        )
    port map (
            in0 => \N__35303\,
            in1 => \N__35134\,
            in2 => \N__34942\,
            in3 => \N__34749\,
            lcout => \this_vga_signals.vaddress_0_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNILD7F7_6_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__36560\,
            in1 => \N__39460\,
            in2 => \N__34624\,
            in3 => \N__37736\,
            lcout => \this_ppu.M_screen_y_q_esr_RNILD7F7Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_data_1_0_i_3_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__35992\,
            in1 => \N__41510\,
            in2 => \N__39898\,
            in3 => \N__36484\,
            lcout => \M_this_spr_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_0_a2_1_x_0_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__42649\,
            in1 => \N__35782\,
            in2 => \_gnd_net_\,
            in3 => \N__43222\,
            lcout => \this_ppu.M_this_state_q_srsts_0_0_a2_1_xZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNIUUE65_6_LC_22_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__34469\,
            in1 => \N__34438\,
            in2 => \N__36567\,
            in3 => \N__36949\,
            lcout => \M_this_ppu_vram_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_en_0_i_0_0_0_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__36477\,
            in1 => \N__36437\,
            in2 => \_gnd_net_\,
            in3 => \N__43431\,
            lcout => \M_this_spr_ram_write_en_0_i_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_0_a2_1_0_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__43799\,
            in1 => \N__42648\,
            in2 => \_gnd_net_\,
            in3 => \N__35719\,
            lcout => \this_ppu.N_1257\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_data_1_0_i_1_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__36478\,
            in1 => \N__39783\,
            in2 => \N__40052\,
            in3 => \N__35988\,
            lcout => \M_this_spr_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_14_LC_22_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__43432\,
            in1 => \N__36438\,
            in2 => \_gnd_net_\,
            in3 => \N__43241\,
            lcout => \M_this_state_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_address_q_0_i_0_a2_1_1_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36335\,
            in2 => \_gnd_net_\,
            in3 => \N__38595\,
            lcout => \N_1258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_1_7_5__m17_0_a3_0_a3_0_a2_LC_22_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35830\,
            in2 => \_gnd_net_\,
            in3 => \N__37785\,
            lcout => \N_1416\,
            ltout => \N_1416_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_1_7_5__m17_0_a3_0_a3_0_a3_2_LC_22_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42240\,
            in2 => \N__35800\,
            in3 => \N__38287\,
            lcout => \N_1151_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_address_q_0_i_0_a3_1_4_LC_22_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__43489\,
            in1 => \N__40747\,
            in2 => \_gnd_net_\,
            in3 => \N__38597\,
            lcout => \N_1066\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_0_a2_1_sx_0_LC_22_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__43855\,
            in1 => \N__35781\,
            in2 => \N__43894\,
            in3 => \N__43220\,
            lcout => \this_ppu.M_this_state_q_srsts_0_0_a2_1_sxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_address_q_0_i_0_a2_0_5_LC_22_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__43488\,
            in1 => \N__36336\,
            in2 => \_gnd_net_\,
            in3 => \N__38596\,
            lcout => \N_1276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_en_0_i_0_0_i_0_LC_22_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__36476\,
            in1 => \N__36445\,
            in2 => \_gnd_net_\,
            in3 => \N__43487\,
            lcout => \M_this_spr_ram_write_en_0_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_address_q_0_i_0_o2_5_LC_22_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__36350\,
            in1 => \N__43502\,
            in2 => \_gnd_net_\,
            in3 => \N__38605\,
            lcout => \N_801_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_substate_d_0_sqmuxa_3_0_a3_0_a3_1_LC_22_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__42614\,
            in1 => \N__36272\,
            in2 => \N__36235\,
            in3 => \N__36152\,
            lcout => \this_ppu_M_this_substate_d_0_sqmuxa_3_0_a3_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_1_1_LC_22_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__39381\,
            in1 => \N__42499\,
            in2 => \_gnd_net_\,
            in3 => \N__38534\,
            lcout => OPEN,
            ltout => \M_this_map_address_qc_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_0_1_LC_22_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__39781\,
            in1 => \N__43503\,
            in2 => \N__36118\,
            in3 => \N__38606\,
            lcout => \M_this_map_address_qc_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_address_q_0_i_0_a2_1_LC_22_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__42262\,
            in1 => \N__43501\,
            in2 => \_gnd_net_\,
            in3 => \N__36115\,
            lcout => \N_1242\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_i_0_0_LC_22_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42443\,
            in2 => \_gnd_net_\,
            in3 => \N__40122\,
            lcout => \N_169_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_1_7_5__N_1048_i_LC_23_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38482\,
            lcout => \N_1048_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_23_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36043\,
            in1 => \N__36028\,
            in2 => \_gnd_net_\,
            in3 => \N__39117\,
            lcout => \this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_23_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36784\,
            in1 => \N__36769\,
            in2 => \_gnd_net_\,
            in3 => \N__39105\,
            lcout => \this_spr_ram.mem_mem_1_1_RNIOA1GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39100\,
            in1 => \N__36748\,
            in2 => \_gnd_net_\,
            in3 => \N__36730\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__37037\,
            in1 => \N__37002\,
            in2 => \N__36715\,
            in3 => \N__39139\,
            lcout => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_7_0_wclke_3_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__38923\,
            in1 => \N__38847\,
            in2 => \N__38795\,
            in3 => \N__38709\,
            lcout => \this_spr_ram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_13_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36676\,
            in1 => \N__39006\,
            in2 => \_gnd_net_\,
            in3 => \N__38204\,
            lcout => \this_spr_ram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39099\,
            in1 => \N__36661\,
            in2 => \_gnd_net_\,
            in3 => \N__36640\,
            lcout => \this_spr_ram.mem_mem_2_1_RNIQE3GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_23_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39098\,
            in1 => \N__36622\,
            in2 => \_gnd_net_\,
            in3 => \N__36610\,
            lcout => \this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_6_LC_23_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__37344\,
            in1 => \N__37290\,
            in2 => \N__37134\,
            in3 => \N__36595\,
            lcout => \this_ppu.M_screen_y_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42059\,
            ce => \N__37177\,
            sr => \N__43098\
        );

    \this_ppu.M_screen_y_q_esr_5_LC_23_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100000000000"
        )
    port map (
            in0 => \N__37343\,
            in1 => \N__37291\,
            in2 => \N__37133\,
            in3 => \N__37264\,
            lcout => \this_ppu.M_screen_y_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42059\,
            ce => \N__37177\,
            sr => \N__43098\
        );

    \this_ppu.M_screen_y_q_esr_RNIJB7F7_5_LC_23_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__37123\,
            in1 => \N__39492\,
            in2 => \N__37093\,
            in3 => \N__37734\,
            lcout => \this_ppu.M_screen_y_q_esr_RNIJB7F7Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNITCNI1_12_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__37000\,
            in1 => \N__36865\,
            in2 => \N__37042\,
            in3 => \N__37009\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNINL8S2_11_LC_23_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__36901\,
            in1 => \N__37001\,
            in2 => \N__36952\,
            in3 => \N__37819\,
            lcout => \M_this_spr_ram_read_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36934\,
            in1 => \N__36919\,
            in2 => \_gnd_net_\,
            in3 => \N__39110\,
            lcout => \this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_23_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39109\,
            in1 => \N__36895\,
            in2 => \_gnd_net_\,
            in3 => \N__36880\,
            lcout => \this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_23_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36859\,
            in1 => \N__36838\,
            in2 => \_gnd_net_\,
            in3 => \N__39112\,
            lcout => \this_spr_ram.mem_mem_3_0_RNIQI5GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_23_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39113\,
            in1 => \N__36820\,
            in2 => \_gnd_net_\,
            in3 => \N__36802\,
            lcout => \this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_1_RNISI5G_LC_23_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37891\,
            in1 => \N__37873\,
            in2 => \_gnd_net_\,
            in3 => \N__39108\,
            lcout => \this_spr_ram.mem_mem_3_1_RNISI5GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_23_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__39111\,
            in1 => \_gnd_net_\,
            in2 => \N__37849\,
            in3 => \N__37831\,
            lcout => \this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_ext_address_q_9_LC_23_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__40606\,
            in1 => \N__43543\,
            in2 => \N__41153\,
            in3 => \N__39784\,
            lcout => \M_this_ext_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42082\,
            ce => 'H',
            sr => \N__43100\
        );

    \M_this_ctrl_flags_q_7_LC_23_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__37800\,
            in1 => \N__40880\,
            in2 => \N__39897\,
            in3 => \N__43544\,
            lcout => \M_this_ctrl_flags_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42093\,
            ce => 'H',
            sr => \N__43103\
        );

    \led_1_7_5__m5_i_a2_i_o3_i_a3_LC_23_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__37399\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37789\,
            lcout => m5_i_a2_i_o3_i_a3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \N_38_i_0_sbtinv_LC_23_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37748\,
            lcout => \N_38_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_this_state_q_7_i_0_0_0_LC_23_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111001001110"
        )
    port map (
            in0 => \N__37459\,
            in1 => \N__43485\,
            in2 => \N__42261\,
            in3 => \N__38285\,
            lcout => \this_ppu_un1_M_this_state_q_7_i_0_0_0\,
            ltout => \this_ppu_un1_M_this_state_q_7_i_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_0_c_RNO_LC_23_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39563\,
            in2 => \N__37441\,
            in3 => \N__39198\,
            lcout => \un1_M_this_map_address_q_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_1_7_5__m12_0_a3_0_a3_0_a3_LC_23_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__37437\,
            in1 => \N__37405\,
            in2 => \N__41130\,
            in3 => \N__37395\,
            lcout => led_c_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_address_q_0_i_0_a3_1_2_LC_23_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__43486\,
            in1 => \N__42774\,
            in2 => \_gnd_net_\,
            in3 => \N__38598\,
            lcout => \N_1058\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_this_state_q_7_i_0_a3_0_0_LC_23_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__40840\,
            in1 => \N__43484\,
            in2 => \_gnd_net_\,
            in3 => \N__38286\,
            lcout => \un1_M_this_state_q_7_i_0_a3_0_0\,
            ltout => \un1_M_this_state_q_7_i_0_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_1_0_LC_23_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100001010"
        )
    port map (
            in0 => \N__38260\,
            in1 => \_gnd_net_\,
            in2 => \N__38254\,
            in3 => \N__39562\,
            lcout => \un1_M_this_map_address_q_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_23_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38251\,
            in1 => \N__38226\,
            in2 => \_gnd_net_\,
            in3 => \N__38198\,
            lcout => \read_data_RNI4PFJ1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_2_LC_23_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__38503\,
            in1 => \N__39298\,
            in2 => \N__37912\,
            in3 => \N__42259\,
            lcout => \M_this_map_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42115\,
            ce => 'H',
            sr => \N__41643\
        );

    \this_ppu.M_this_map_address_q_0_i_0_a3_1_3_LC_23_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__41509\,
            in1 => \N__43499\,
            in2 => \_gnd_net_\,
            in3 => \N__38608\,
            lcout => OPEN,
            ltout => \N_1062_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_3_LC_23_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__37897\,
            in1 => \N__39253\,
            in2 => \N__37900\,
            in3 => \N__42260\,
            lcout => \M_this_map_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42115\,
            ce => 'H',
            sr => \N__41643\
        );

    \M_this_map_address_q_RNO_0_3_LC_23_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__39273\,
            in1 => \N__42529\,
            in2 => \_gnd_net_\,
            in3 => \N__38532\,
            lcout => \M_this_map_address_qc_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_0_4_LC_23_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__38533\,
            in1 => \_gnd_net_\,
            in2 => \N__42542\,
            in3 => \N__39228\,
            lcout => OPEN,
            ltout => \M_this_map_address_qc_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_4_LC_23_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__42258\,
            in1 => \N__38617\,
            in2 => \N__38611\,
            in3 => \N__39208\,
            lcout => \M_this_map_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42115\,
            ce => 'H',
            sr => \N__41643\
        );

    \this_ppu.M_this_map_address_q_0_i_0_a3_1_0_LC_23_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__42445\,
            in1 => \N__43500\,
            in2 => \_gnd_net_\,
            in3 => \N__38607\,
            lcout => \N_1097\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_0_0_LC_23_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__39547\,
            in1 => \N__42507\,
            in2 => \_gnd_net_\,
            in3 => \N__38535\,
            lcout => \M_this_map_address_qc_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_0_2_LC_23_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__38536\,
            in1 => \N__39318\,
            in2 => \_gnd_net_\,
            in3 => \N__42508\,
            lcout => \M_this_map_address_qc_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_i_0_1_LC_23_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39761\,
            in2 => \_gnd_net_\,
            in3 => \N__40150\,
            lcout => \N_918_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \N_1048_sbtinv_LC_23_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38478\,
            lcout => \N_1048_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_0_wclke_3_LC_24_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__38921\,
            in1 => \N__38859\,
            in2 => \N__38793\,
            in3 => \N__38719\,
            lcout => \this_spr_ram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_0_wclke_3_LC_24_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__38717\,
            in1 => \N__38904\,
            in2 => \N__38858\,
            in3 => \N__38759\,
            lcout => \this_spr_ram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_0_wclke_3_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38903\,
            in1 => \N__38839\,
            in2 => \N__38776\,
            in3 => \N__38716\,
            lcout => \this_spr_ram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_0_wclke_3_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__38922\,
            in1 => \N__38865\,
            in2 => \N__38794\,
            in3 => \N__38718\,
            lcout => \this_spr_ram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39163\,
            in1 => \N__39097\,
            in2 => \_gnd_net_\,
            in3 => \N__39154\,
            lcout => \this_spr_ram.mem_mem_0_0_RNIK6VFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_24_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39133\,
            in1 => \N__39104\,
            in2 => \_gnd_net_\,
            in3 => \N__39034\,
            lcout => \this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.IO_port_data_write_i_m2_i_m2_7_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39415\,
            in1 => \N__43681\,
            in2 => \_gnd_net_\,
            in3 => \N__39010\,
            lcout => \IO_port_data_write_i_m2_i_m2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_4_0_wclke_3_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__38924\,
            in1 => \N__38861\,
            in2 => \N__38796\,
            in3 => \N__38701\,
            lcout => \this_spr_ram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_5_0_wclke_3_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__38702\,
            in1 => \N__38789\,
            in2 => \N__38866\,
            in3 => \N__38925\,
            lcout => \this_spr_ram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_6_0_wclke_3_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__38926\,
            in1 => \N__38860\,
            in2 => \N__38797\,
            in3 => \N__38703\,
            lcout => \this_spr_ram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_ext_address_q_0_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000010010"
        )
    port map (
            in0 => \N__40312\,
            in1 => \N__43528\,
            in2 => \N__40281\,
            in3 => \N__41145\,
            lcout => \M_this_ext_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42101\,
            ce => 'H',
            sr => \N__43101\
        );

    \M_this_status_flags_q_7_LC_24_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39461\,
            lcout => \M_this_status_flags_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42101\,
            ce => 'H',
            sr => \N__43101\
        );

    \M_this_map_address_q_1_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011000100"
        )
    port map (
            in0 => \N__42288\,
            in1 => \N__39406\,
            in2 => \N__39377\,
            in3 => \N__39340\,
            lcout => \M_this_map_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42109\,
            ce => 'H',
            sr => \N__41647\
        );

    \un1_M_this_map_address_q_cry_0_c_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39394\,
            in2 => \N__39564\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_24_23_0_\,
            carryout => \un1_M_this_map_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_0_THRU_LUT4_0_LC_24_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39364\,
            in2 => \_gnd_net_\,
            in3 => \N__39334\,
            lcout => \un1_M_this_map_address_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_0\,
            carryout => \un1_M_this_map_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_1_2_LC_24_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39317\,
            in2 => \_gnd_net_\,
            in3 => \N__39292\,
            lcout => \M_this_map_address_q_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_1\,
            carryout => \un1_M_this_map_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_1_3_LC_24_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39272\,
            in2 => \_gnd_net_\,
            in3 => \N__39247\,
            lcout => \M_this_map_address_q_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_2\,
            carryout => \un1_M_this_map_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_1_4_LC_24_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39227\,
            in2 => \_gnd_net_\,
            in3 => \N__39202\,
            lcout => \M_this_map_address_q_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_3\,
            carryout => \un1_M_this_map_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_1_5_LC_24_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39199\,
            in2 => \N__42183\,
            in3 => \N__39187\,
            lcout => \M_this_map_address_q_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_4\,
            carryout => \un1_M_this_map_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_5_THRU_LUT4_0_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39632\,
            in2 => \_gnd_net_\,
            in3 => \N__39805\,
            lcout => \un1_M_this_map_address_q_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_5\,
            carryout => \un1_M_this_map_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_6_THRU_LUT4_0_LC_24_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42869\,
            in2 => \_gnd_net_\,
            in3 => \N__39802\,
            lcout => \un1_M_this_map_address_q_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_6\,
            carryout => \un1_M_this_map_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_map_address_q_cry_7_THRU_LUT4_0_LC_24_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41542\,
            in2 => \_gnd_net_\,
            in3 => \N__39799\,
            lcout => \un1_M_this_map_address_q_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_24_24_0_\,
            carryout => \un1_M_this_map_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_9_LC_24_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110010001100"
        )
    port map (
            in0 => \N__40808\,
            in1 => \N__40651\,
            in2 => \N__42295\,
            in3 => \N__39796\,
            lcout => \M_this_map_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42120\,
            ce => 'H',
            sr => \N__41645\
        );

    \M_this_map_address_q_RNO_0_6_LC_24_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010100001101"
        )
    port map (
            in0 => \N__42834\,
            in1 => \N__42283\,
            in2 => \N__39633\,
            in3 => \N__39793\,
            lcout => OPEN,
            ltout => \M_this_map_address_qc_8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_6_LC_24_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__39777\,
            in1 => \N__42588\,
            in2 => \N__39649\,
            in3 => \N__42541\,
            lcout => \M_this_map_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42124\,
            ce => 'H',
            sr => \N__41644\
        );

    \M_this_map_address_q_8_LC_24_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100000000"
        )
    port map (
            in0 => \N__42284\,
            in1 => \N__39604\,
            in2 => \N__41550\,
            in3 => \N__41383\,
            lcout => \M_this_map_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42124\,
            ce => 'H',
            sr => \N__41644\
        );

    \M_this_map_address_q_0_LC_24_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__39598\,
            in1 => \N__39589\,
            in2 => \N__39583\,
            in3 => \N__42289\,
            lcout => \M_this_map_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42129\,
            ce => 'H',
            sr => \N__41642\
        );

    \this_ppu.M_this_map_ram_write_data_i_0_4_LC_24_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40685\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40129\,
            lcout => \N_921_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_i_0_2_LC_24_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__42750\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40151\,
            lcout => \N_919_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_i_0_6_LC_24_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40153\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40397\,
            lcout => \N_923_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_i_0_3_LC_24_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41466\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40152\,
            lcout => \N_920_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_i_0_5_LC_24_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40154\,
            in2 => \_gnd_net_\,
            in3 => \N__40061\,
            lcout => \N_922_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_i_0_7_LC_24_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40155\,
            in2 => \_gnd_net_\,
            in3 => \N__39905\,
            lcout => \N_924_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_ext_address_q_13_LC_26_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__40555\,
            in1 => \N__43566\,
            in2 => \N__41160\,
            in3 => \N__40012\,
            lcout => \M_this_ext_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42096\,
            ce => 'H',
            sr => \N__43097\
        );

    \M_this_ctrl_flags_q_5_LC_26_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__43564\,
            in1 => \N__39945\,
            in2 => \N__40032\,
            in3 => \N__40890\,
            lcout => \M_this_ctrl_flags_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42096\,
            ce => 'H',
            sr => \N__43097\
        );

    \M_this_ext_address_q_2_LC_26_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000010010"
        )
    port map (
            in0 => \N__40210\,
            in1 => \N__43568\,
            in2 => \N__40236\,
            in3 => \N__41152\,
            lcout => \M_this_ext_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42096\,
            ce => 'H',
            sr => \N__43097\
        );

    \M_this_ext_address_q_15_LC_26_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__41151\,
            in1 => \N__39838\,
            in2 => \N__43576\,
            in3 => \N__41035\,
            lcout => \M_this_ext_address_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42096\,
            ce => 'H',
            sr => \N__43097\
        );

    \M_this_ctrl_flags_q_6_LC_26_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__43565\,
            in1 => \N__40458\,
            in2 => \N__40419\,
            in3 => \N__40891\,
            lcout => \M_this_ctrl_flags_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42096\,
            ce => 'H',
            sr => \N__43097\
        );

    \M_this_ext_address_q_14_LC_26_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__40519\,
            in1 => \N__43567\,
            in2 => \N__41161\,
            in3 => \N__40404\,
            lcout => \M_this_ext_address_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42096\,
            ce => 'H',
            sr => \N__43097\
        );

    \un1_M_this_ext_address_q_cry_0_c_LC_26_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40311\,
            in2 => \N__40280\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_26_21_0_\,
            carryout => \un1_M_this_ext_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_0_THRU_LUT4_0_LC_26_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41288\,
            in2 => \_gnd_net_\,
            in3 => \N__40249\,
            lcout => \un1_M_this_ext_address_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_0\,
            carryout => \un1_M_this_ext_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_1_THRU_LUT4_0_LC_26_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40232\,
            in2 => \_gnd_net_\,
            in3 => \N__40201\,
            lcout => \un1_M_this_ext_address_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_1\,
            carryout => \un1_M_this_ext_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_2_THRU_LUT4_0_LC_26_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41249\,
            in2 => \_gnd_net_\,
            in3 => \N__40198\,
            lcout => \un1_M_this_ext_address_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_2\,
            carryout => \un1_M_this_ext_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_3_THRU_LUT4_0_LC_26_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41213\,
            in2 => \_gnd_net_\,
            in3 => \N__40195\,
            lcout => \un1_M_this_ext_address_q_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_3\,
            carryout => \un1_M_this_ext_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_4_THRU_LUT4_0_LC_26_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41177\,
            in2 => \_gnd_net_\,
            in3 => \N__40192\,
            lcout => \un1_M_this_ext_address_q_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_4\,
            carryout => \un1_M_this_ext_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_5_THRU_LUT4_0_LC_26_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43275\,
            in3 => \N__40189\,
            lcout => \un1_M_this_ext_address_q_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_5\,
            carryout => \un1_M_this_ext_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_6_THRU_LUT4_0_LC_26_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40971\,
            in2 => \_gnd_net_\,
            in3 => \N__40642\,
            lcout => \un1_M_this_ext_address_q_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_6\,
            carryout => \un1_M_this_ext_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_7_c_RNIQ14F_LC_26_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41322\,
            in2 => \_gnd_net_\,
            in3 => \N__40639\,
            lcout => \un1_M_this_ext_address_q_cry_7_c_RNIQ14FZ0\,
            ltout => OPEN,
            carryin => \bfn_26_22_0_\,
            carryout => \un1_M_this_ext_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_8_c_RNIS45F_LC_26_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40626\,
            in2 => \_gnd_net_\,
            in3 => \N__40594\,
            lcout => \un1_M_this_ext_address_q_cry_8_c_RNIS45FZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_8\,
            carryout => \un1_M_this_ext_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_9_c_RNI55NH_LC_26_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41004\,
            in2 => \_gnd_net_\,
            in3 => \N__40591\,
            lcout => \un1_M_this_ext_address_q_cry_9_c_RNI55NHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_9\,
            carryout => \un1_M_this_ext_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_10_c_RNIEGOA_LC_26_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40929\,
            in2 => \_gnd_net_\,
            in3 => \N__40588\,
            lcout => \un1_M_this_ext_address_q_cry_10_c_RNIEGOAZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_10\,
            carryout => \un1_M_this_ext_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_11_c_RNIGJPA_LC_26_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40902\,
            in2 => \_gnd_net_\,
            in3 => \N__40585\,
            lcout => \un1_M_this_ext_address_q_cry_11_c_RNIGJPAZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_11\,
            carryout => \un1_M_this_ext_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_12_c_RNIIMQA_LC_26_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40572\,
            in2 => \_gnd_net_\,
            in3 => \N__40546\,
            lcout => \un1_M_this_ext_address_q_cry_12_c_RNIIMQAZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_12\,
            carryout => \un1_M_this_ext_address_q_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_13_c_RNIKPRA_LC_26_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40536\,
            in2 => \_gnd_net_\,
            in3 => \N__40510\,
            lcout => \un1_M_this_ext_address_q_cry_13_c_RNIKPRAZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_13\,
            carryout => \un1_M_this_ext_address_q_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_14_c_RNIMSSA_LC_26_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40503\,
            in2 => \_gnd_net_\,
            in3 => \N__41038\,
            lcout => \un1_M_this_ext_address_q_cry_14_c_RNIMSSAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_ext_address_q_10_LC_26_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__41026\,
            in1 => \N__41097\,
            in2 => \N__42757\,
            in3 => \N__43561\,
            lcout => \M_this_ext_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42125\,
            ce => 'H',
            sr => \N__43102\
        );

    \M_this_ext_address_q_7_LC_26_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001110001100"
        )
    port map (
            in0 => \N__41096\,
            in1 => \N__40967\,
            in2 => \N__43575\,
            in3 => \N__40993\,
            lcout => \M_this_ext_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42125\,
            ce => 'H',
            sr => \N__43102\
        );

    \M_this_ext_address_q_11_LC_26_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__40948\,
            in1 => \N__41454\,
            in2 => \N__41129\,
            in3 => \N__43562\,
            lcout => \M_this_ext_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42125\,
            ce => 'H',
            sr => \N__43102\
        );

    \M_this_ext_address_q_12_LC_26_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__41095\,
            in1 => \N__40709\,
            in2 => \N__43574\,
            in3 => \N__40918\,
            lcout => \M_this_ext_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42125\,
            ce => 'H',
            sr => \N__43102\
        );

    \M_this_ctrl_flags_q_4_LC_26_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__40881\,
            in1 => \N__40839\,
            in2 => \N__40726\,
            in3 => \N__43563\,
            lcout => \M_this_ctrl_flags_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42125\,
            ce => 'H',
            sr => \N__43102\
        );

    \this_ppu.M_this_map_address_q_0_i_0_a3_9_LC_26_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40812\,
            in2 => \_gnd_net_\,
            in3 => \N__42828\,
            lcout => OPEN,
            ltout => \N_1081_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_0_9_LC_26_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__40705\,
            in1 => \N__42593\,
            in2 => \N__40654\,
            in3 => \N__42543\,
            lcout => \M_this_map_address_qc_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_address_q_0_i_0_a3_5_LC_26_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42167\,
            in2 => \_gnd_net_\,
            in3 => \N__42829\,
            lcout => \N_1068\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_address_q_0_i_0_a3_8_LC_26_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__42830\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41549\,
            lcout => OPEN,
            ltout => \N_1078_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_0_8_LC_26_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__41470\,
            in1 => \N__42540\,
            in2 => \N__41386\,
            in3 => \N__42594\,
            lcout => \M_this_map_address_qc_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.IO_port_data_write_0_a2_i_2_LC_26_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__43703\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41364\,
            lcout => \N_726_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_ext_address_q_8_LC_27_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__41341\,
            in1 => \N__41133\,
            in2 => \N__42463\,
            in3 => \N__43545\,
            lcout => \M_this_ext_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42126\,
            ce => 'H',
            sr => \N__43099\
        );

    \M_this_ext_address_q_1_LC_27_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100001011010"
        )
    port map (
            in0 => \N__41311\,
            in1 => \N__41134\,
            in2 => \N__41295\,
            in3 => \N__43546\,
            lcout => \M_this_ext_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42126\,
            ce => 'H',
            sr => \N__43099\
        );

    \M_this_ext_address_q_3_LC_27_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100001011010"
        )
    port map (
            in0 => \N__41272\,
            in1 => \N__41135\,
            in2 => \N__41256\,
            in3 => \N__43547\,
            lcout => \M_this_ext_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42126\,
            ce => 'H',
            sr => \N__43099\
        );

    \M_this_ext_address_q_4_LC_27_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001110001100"
        )
    port map (
            in0 => \N__41131\,
            in1 => \N__41214\,
            in2 => \N__43572\,
            in3 => \N__41233\,
            lcout => \M_this_ext_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42126\,
            ce => 'H',
            sr => \N__43099\
        );

    \M_this_ext_address_q_5_LC_27_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100001011010"
        )
    port map (
            in0 => \N__41197\,
            in1 => \N__41136\,
            in2 => \N__41184\,
            in3 => \N__43548\,
            lcout => \M_this_ext_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42126\,
            ce => 'H',
            sr => \N__43099\
        );

    \M_this_ext_address_q_6_LC_27_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001110001100"
        )
    port map (
            in0 => \N__41132\,
            in1 => \N__43271\,
            in2 => \N__43573\,
            in3 => \N__43285\,
            lcout => \M_this_ext_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42126\,
            ce => 'H',
            sr => \N__43099\
        );

    \M_this_map_address_q_7_LC_27_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010101010"
        )
    port map (
            in0 => \N__42655\,
            in1 => \N__42895\,
            in2 => \N__42870\,
            in3 => \N__42293\,
            lcout => \M_this_map_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42132\,
            ce => 'H',
            sr => \N__41650\
        );

    \this_ppu.M_this_map_address_q_0_i_0_a3_7_LC_27_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42859\,
            in2 => \_gnd_net_\,
            in3 => \N__42835\,
            lcout => OPEN,
            ltout => \N_1075_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_0_7_LC_27_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__42710\,
            in1 => \N__42595\,
            in2 => \N__42658\,
            in3 => \N__42544\,
            lcout => \M_this_map_address_qc_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_substate_d_0_sqmuxa_3_0_o2_LC_27_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43854\,
            in1 => \N__42636\,
            in2 => \N__43887\,
            in3 => \N__43813\,
            lcout => \N_459_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_RNO_0_5_LC_27_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__42592\,
            in1 => \N__42539\,
            in2 => \N__42459\,
            in3 => \N__42319\,
            lcout => \M_this_map_address_qc_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_5_LC_27_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__42313\,
            in1 => \N__42307\,
            in2 => \_gnd_net_\,
            in3 => \N__42294\,
            lcout => \M_this_map_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42137\,
            ce => 'H',
            sr => \N__41646\
        );

    \this_vga_signals.IO_port_data_write_0_a2_i_6_LC_28_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__43696\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41601\,
            lcout => \N_734_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.IO_port_data_write_0_a2_i_5_LC_28_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__43936\,
            in1 => \N__43695\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_996_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_substate_d_0_sqmuxa_3_0_o2_x_LC_28_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__43874\,
            in1 => \N__43847\,
            in2 => \_gnd_net_\,
            in3 => \N__43806\,
            lcout => \M_this_substate_d_0_sqmuxa_3_0_o2_x\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.IO_port_data_write_0_a2_i_4_LC_28_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__43704\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43746\,
            lcout => \N_730_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.IO_port_data_write_0_a2_i_3_LC_28_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__43705\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43608\,
            lcout => \N_728_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
