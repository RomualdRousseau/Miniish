-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     May 27 2022 09:13:54

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : inout std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    debug : out std_logic_vector(1 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    led : out std_logic_vector(7 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : inout std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__33435\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal port_nmib_0_i : std_logic;
signal this_vga_signals_vvisibility_i : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_1\ : std_logic;
signal rgb_c_2 : std_logic;
signal port_clk_c : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_0\ : std_logic;
signal \M_this_oam_address_qZ0Z_0\ : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal \M_this_oam_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_oam_address_q_cry_0\ : std_logic;
signal \M_this_oam_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_oam_address_q_cry_1\ : std_logic;
signal \M_this_oam_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_oam_address_q_cry_2\ : std_logic;
signal \M_this_oam_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_oam_address_q_cry_3\ : std_logic;
signal \un1_M_this_oam_address_q_cry_4\ : std_logic;
signal \M_this_oam_address_qZ0Z_5\ : std_logic;
signal \this_oam_ram.M_this_oam_ram_read_data_19\ : std_logic;
signal \M_this_data_tmp_qZ0Z_26\ : std_logic;
signal \M_this_oam_ram_write_data_26\ : std_logic;
signal \M_this_oam_ram_write_data_20\ : std_logic;
signal \N_892_0\ : std_logic;
signal rgb_c_0 : std_logic;
signal rgb_c_3 : std_logic;
signal rgb_c_4 : std_logic;
signal \N_834_0\ : std_logic;
signal \N_818_0\ : std_logic;
signal \N_837_0\ : std_logic;
signal \M_this_oam_ram_write_data_5\ : std_logic;
signal \M_this_oam_ram_write_data_8\ : std_logic;
signal \N_836_0\ : std_logic;
signal \N_896_0\ : std_logic;
signal \M_this_oam_ram_write_data_4\ : std_logic;
signal \N_895_0\ : std_logic;
signal \N_891_0\ : std_logic;
signal \this_oam_ram.M_this_oam_ram_read_data_10\ : std_logic;
signal \this_oam_ram.M_this_oam_ram_read_data_11\ : std_logic;
signal \M_this_oam_ram_write_data_28\ : std_logic;
signal \N_894_0\ : std_logic;
signal \N_889_0\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_i_16\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_0\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_1\ : std_logic;
signal \M_this_oam_ram_read_data_i_19\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_2\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_3\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_4\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_5\ : std_logic;
signal \M_this_oam_ram_read_data_23\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_6\ : std_logic;
signal \this_oam_ram.M_this_oam_ram_read_data_21\ : std_logic;
signal \M_this_oam_ram_read_data_i_21\ : std_logic;
signal \M_this_oam_ram_write_data_0\ : std_logic;
signal \this_oam_ram.M_this_oam_ram_read_data_12\ : std_logic;
signal \this_oam_ram.M_this_oam_ram_read_data_17\ : std_logic;
signal \M_this_oam_ram_read_data_i_17\ : std_logic;
signal \this_oam_ram.M_this_oam_ram_read_data_18\ : std_logic;
signal \M_this_oam_ram_read_data_i_18\ : std_logic;
signal \this_oam_ram.M_this_oam_ram_read_data_20\ : std_logic;
signal \M_this_oam_ram_read_data_i_20\ : std_logic;
signal \this_pixel_clk_M_counter_q_i_1\ : std_logic;
signal \this_pixel_clk_M_counter_q_0\ : std_logic;
signal rgb_c_1 : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal \N_816_0\ : std_logic;
signal \this_vga_ramdac.N_2612_reto\ : std_logic;
signal \M_this_map_address_qZ0Z_0\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \M_this_map_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_map_address_q_cry_0\ : std_logic;
signal \M_this_map_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_map_address_q_cry_1\ : std_logic;
signal \M_this_map_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_map_address_q_cry_2\ : std_logic;
signal \M_this_map_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_map_address_q_cry_3\ : std_logic;
signal \M_this_map_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_map_address_q_cry_4\ : std_logic;
signal \M_this_map_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_5\ : std_logic;
signal \M_this_map_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_map_address_q_cry_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_7\ : std_logic;
signal \M_this_map_address_qZ0Z_8\ : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal \un1_M_this_map_address_q_cry_8\ : std_logic;
signal \M_this_map_address_qZ0Z_9\ : std_logic;
signal \this_vga_ramdac.i2_mux\ : std_logic;
signal \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\ : std_logic;
signal rgb_c_5 : std_logic;
signal \N_60_0\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal \M_this_map_ram_read_data_1\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_6_c_RNIP5LZ0Z8\ : std_logic;
signal \M_this_ppu_sprites_addr_7\ : std_logic;
signal \M_this_data_tmp_qZ0Z_15\ : std_logic;
signal \M_this_data_tmp_qZ0Z_8\ : std_logic;
signal \M_this_data_tmp_qZ0Z_11\ : std_logic;
signal \N_835_0\ : std_logic;
signal \N_897_0\ : std_logic;
signal \N_53_0\ : std_logic;
signal \M_this_oam_ram_write_data_2\ : std_logic;
signal \N_890_0\ : std_logic;
signal \M_this_oam_ram_write_data_12\ : std_logic;
signal \N_831_0\ : std_logic;
signal \M_this_oam_ram_write_data_24\ : std_logic;
signal \N_832_0\ : std_logic;
signal \N_893_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_19\ : std_logic;
signal \M_this_data_tmp_qZ0Z_20\ : std_logic;
signal \M_this_data_tmp_qZ0Z_21\ : std_logic;
signal \M_this_data_tmp_qZ0Z_22\ : std_logic;
signal \M_this_data_tmp_qZ0Z_23\ : std_logic;
signal \this_oam_ram.M_this_oam_ram_read_data_22\ : std_logic;
signal \M_this_oam_ram_read_data_i_22\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals.if_m2_0\ : std_logic;
signal \N_58_0\ : std_logic;
signal \N_3_0_cascade_\ : std_logic;
signal \G_480_cascade_\ : std_logic;
signal \this_vga_ramdac.N_2614_reto\ : std_logic;
signal \this_vga_ramdac.N_2611_reto\ : std_logic;
signal \this_vga_ramdac.N_2610_reto\ : std_logic;
signal \N_2_0\ : std_logic;
signal \N_2_0_cascade_\ : std_logic;
signal \M_this_vga_signals_pixel_clk_0_0\ : std_logic;
signal \this_vga_ramdac.i2_mux_0_cascade_\ : std_logic;
signal \this_vga_ramdac.N_2615_reto\ : std_logic;
signal \this_vga_ramdac.m16_cascade_\ : std_logic;
signal \G_480\ : std_logic;
signal \this_vga_ramdac.N_2613_reto\ : std_logic;
signal \N_73_0\ : std_logic;
signal \this_vga_ramdac.N_24_mux\ : std_logic;
signal \this_vga_ramdac.m19\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \this_vga_ramdac.m6\ : std_logic;
signal \M_this_data_tmp_qZ0Z_14\ : std_logic;
signal \M_this_data_tmp_qZ0Z_27\ : std_logic;
signal \M_this_data_tmp_qZ0Z_3\ : std_logic;
signal \M_this_data_tmp_qZ0Z_7\ : std_logic;
signal \M_this_data_tmp_qZ0Z_2\ : std_logic;
signal \M_this_data_tmp_qZ0Z_4\ : std_logic;
signal \M_this_data_tmp_qZ0Z_25\ : std_logic;
signal \M_this_data_tmp_qZ0Z_31\ : std_logic;
signal \M_this_data_tmp_qZ0Z_28\ : std_logic;
signal \N_833_0\ : std_logic;
signal \M_this_oam_ram_read_data_16\ : std_logic;
signal \M_this_ppu_vram_addr_i_6\ : std_logic;
signal \M_this_data_tmp_qZ0Z_18\ : std_logic;
signal \M_this_oam_ram_write_data_18\ : std_logic;
signal \M_this_ppu_map_addr_4\ : std_logic;
signal \M_this_data_tmp_qZ0Z_30\ : std_logic;
signal \N_830_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_16\ : std_logic;
signal \M_this_oam_ram_write_data_16\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1\ : std_logic;
signal \this_vga_signals.if_i4_mux_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.M_hcounter_q_RNIUULS4Z0Z_3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.if_m2_2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_3_1_cascade_\ : std_logic;
signal \this_vga_signals.d_N_3_0_i\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_axbxc3_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c3_0\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_1_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2\ : std_logic;
signal \this_vga_signals.SUM_3\ : std_logic;
signal \N_3_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_0\ : std_logic;
signal \this_vga_signals.N_17_0\ : std_logic;
signal \this_vga_signals.M_hcounter_q_RNI9JJM1Z0Z_0\ : std_logic;
signal \this_vga_signals.M_hcounter_q_RNIADGD1Z0Z_5_cascade_\ : std_logic;
signal this_vga_signals_hvisibility_i : std_logic;
signal \this_vga_signals.i5_mux\ : std_logic;
signal this_vga_signals_hsync_1_i : std_logic;
signal \M_this_ppu_map_addr_9\ : std_logic;
signal \N_63_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_3\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal \this_vga_signals.SUM_3_1\ : std_logic;
signal \M_this_vga_signals_address_6\ : std_logic;
signal \M_this_data_tmp_qZ0Z_29\ : std_logic;
signal \M_this_data_tmp_qZ0Z_5\ : std_logic;
signal \M_this_data_tmp_qZ0Z_12\ : std_logic;
signal \M_this_data_tmp_qZ0Z_13\ : std_logic;
signal \M_this_data_tmp_qZ0Z_9\ : std_logic;
signal \M_this_data_tmp_qZ0Z_0\ : std_logic;
signal \M_this_ppu_vram_data_0_cascade_\ : std_logic;
signal \this_ppu.N_134_cascade_\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c2_cascade_\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c5\ : std_logic;
signal \M_this_ppu_vram_addr_6\ : std_logic;
signal \M_this_ppu_map_addr_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c5_cascade_\ : std_logic;
signal \this_ppu.M_haddress_qZ0Z_7\ : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_12_22_0_\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_3_0\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_0\ : std_logic;
signal \N_815_0\ : std_logic;
signal \N_814_0\ : std_logic;
signal \this_ppu_M_vaddress_q_i_6\ : std_logic;
signal \M_this_data_tmp_qZ0Z_1\ : std_logic;
signal \M_this_data_tmp_qZ0Z_24\ : std_logic;
signal \M_this_data_tmp_qZ0Z_6\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_1_c_RNITOBZ0Z8\ : std_logic;
signal \M_this_ppu_sprites_addr_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c1_cascade_\ : std_logic;
signal \M_this_ppu_vram_en_0\ : std_logic;
signal \this_ppu.N_134\ : std_logic;
signal \M_this_ppu_map_addr_0\ : std_logic;
signal \M_this_ppu_vram_addr_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c2\ : std_logic;
signal \M_this_ppu_map_addr_1\ : std_logic;
signal \this_ppu.N_128\ : std_logic;
signal \this_ppu.M_state_qc_1_3\ : std_logic;
signal \M_this_ppu_vram_data_0\ : std_logic;
signal \this_ppu.M_state_qc_1_1_cascade_\ : std_logic;
signal \this_ppu.M_state_qZ0Z_4\ : std_logic;
signal \this_ppu.M_state_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.N_18_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.m23_1_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.N_1090_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \G_464\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \M_this_oam_ram_write_data_10\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_0_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_1_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_2_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_3_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_4_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_5_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_6_s1\ : std_logic;
signal \this_ppu.M_state_d_0_sqmuxa_1_cascade_\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\ : std_logic;
signal \this_ppu.N_1456_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_5\ : std_logic;
signal \this_ppu.M_count_qZ0Z_4\ : std_logic;
signal \this_ppu.M_count_qZ0Z_1\ : std_logic;
signal \this_ppu.M_state_q_RNIE20V4Z0Z_0\ : std_logic;
signal \M_this_vga_signals_line_clk_0_cascade_\ : std_logic;
signal \this_ppu.M_state_d_0_sqmuxa_cascade_\ : std_logic;
signal \this_vga_signals.N_1000_cascade_\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.i21_mux_cascade_\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_1\ : std_logic;
signal \N_817_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_10\ : std_logic;
signal \M_this_data_tmp_qZ0Z_17\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_3\ : std_logic;
signal \this_ppu.M_count_qZ0Z_0\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_2\ : std_logic;
signal \M_this_map_ram_read_data_2\ : std_logic;
signal \this_ppu.un10_sprites_addr_axb_0_cascade_\ : std_logic;
signal \M_this_ppu_sprites_addr_8\ : std_logic;
signal \this_ppu.un10_0\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\ : std_logic;
signal \this_ppu.N_1456_0\ : std_logic;
signal \this_ppu.M_count_qZ0Z_6\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_2_c_RNIVRCZ0Z8\ : std_logic;
signal \M_this_ppu_sprites_addr_3\ : std_logic;
signal \this_oam_ram.M_this_oam_ram_read_data_9\ : std_logic;
signal \M_this_map_ram_read_data_3\ : std_logic;
signal \M_this_ppu_sprites_addr_9\ : std_logic;
signal \this_ppu.M_state_d_0_sqmuxa_1\ : std_logic;
signal \this_ppu.M_count_q_RNO_0Z0Z_7\ : std_logic;
signal \this_ppu.M_count_qZ0Z_7\ : std_logic;
signal \this_vga_signals.N_129_mux\ : std_logic;
signal \this_vga_signals.N_1028\ : std_logic;
signal \this_vga_signals.N_1028_cascade_\ : std_logic;
signal \this_vga_signals.N_999\ : std_logic;
signal \this_vga_signals.N_1004_cascade_\ : std_logic;
signal \this_vga_signals.N_1013\ : std_logic;
signal \this_vga_signals.N_1013_cascade_\ : std_logic;
signal \this_vga_signals.N_105_mux_cascade_\ : std_logic;
signal \this_vga_signals.N_113_mux\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_4\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_5\ : std_logic;
signal this_vga_signals_vvisibility : std_logic;
signal \M_this_reset_cond_out_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_6\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_7\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_8\ : std_logic;
signal \this_vga_signals.vaddress_ac0_9_0_a0_2\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_6\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_c5\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_7\ : std_logic;
signal dma_0_i : std_logic;
signal \N_1430_0\ : std_logic;
signal \M_this_state_q_ns_17_cascade_\ : std_logic;
signal \M_this_state_q_ns_0_17\ : std_logic;
signal \M_this_map_ram_read_data_6\ : std_logic;
signal \M_this_oam_ram_read_data_8\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_iZ0Z_8\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \M_this_oam_ram_read_data_i_9\ : std_logic;
signal \this_ppu.un10_sprites_addr_cry_0_c_RNIMJ5BZ0\ : std_logic;
signal \this_ppu.un10_sprites_addr_cry_0\ : std_logic;
signal \M_this_oam_ram_read_data_i_10\ : std_logic;
signal \this_ppu.un10_sprites_addr_cry_1\ : std_logic;
signal \M_this_oam_ram_read_data_i_11\ : std_logic;
signal \this_ppu.un10_sprites_addr_cry_2\ : std_logic;
signal \M_this_oam_ram_read_data_i_12\ : std_logic;
signal \this_ppu.un10_sprites_addr_cry_3_c_RNISS8BZ0\ : std_logic;
signal \this_ppu.un10_sprites_addr_cry_3\ : std_logic;
signal \M_this_oam_ram_read_data_13\ : std_logic;
signal \this_ppu.un10_sprites_addr_cry_4\ : std_logic;
signal \this_ppu.M_last_q\ : std_logic;
signal \this_ppu.M_state_qZ0Z_0\ : std_logic;
signal \M_this_vga_signals_line_clk_0\ : std_logic;
signal \this_ppu.M_state_d_0_sqmuxa\ : std_logic;
signal \M_this_ppu_vram_addr_7\ : std_logic;
signal \M_this_ppu_map_addr_7\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_c3\ : std_logic;
signal \M_this_ppu_map_addr_5\ : std_logic;
signal \M_this_ppu_map_addr_6\ : std_logic;
signal \this_ppu.M_state_q_RNIELANCZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNI4KCU6Z0Z_9\ : std_logic;
signal \this_vga_signals.g1_2_0_0_cascade_\ : std_logic;
signal \M_this_vga_ramdac_en_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c3_0_0_0_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \this_vga_signals.un6_vvisibilitylt9_0\ : std_logic;
signal \this_vga_signals.g2_2\ : std_logic;
signal \this_vga_signals.SUM_2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_1_1_cascade_\ : std_logic;
signal \this_vga_signals.N_4_0_0_0\ : std_logic;
signal \this_vga_signals.g3_2_0\ : std_logic;
signal \this_vga_signals.N_6_cascade_\ : std_logic;
signal \this_vga_signals.g4\ : std_logic;
signal \N_1438_0\ : std_logic;
signal \this_start_data_delay.port_data_rw_0_a2Z0Z_1\ : std_logic;
signal port_data_rw_0_i : std_logic;
signal \this_sprites_ram.mem_out_bus5_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_2\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_2\ : std_logic;
signal \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\ : std_logic;
signal \M_this_ppu_vram_data_2\ : std_logic;
signal \this_ppu.un10_sprites_addr_cry_2_c_RNIQP7BZ0\ : std_logic;
signal \M_this_map_ram_read_data_5\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_2\ : std_logic;
signal \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_1\ : std_logic;
signal \this_ppu.M_state_q_srsts_i_a3_5_2\ : std_logic;
signal \this_ppu.M_state_q_srsts_i_a3_4_2\ : std_logic;
signal \N_2_cascade_\ : std_logic;
signal \this_vga_signals.N_6_1_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_N_4_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb1_i_1\ : std_logic;
signal \this_vga_signals.N_7_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0\ : std_logic;
signal \this_vga_signals.if_m2_3_1_cascade_\ : std_logic;
signal \this_vga_signals.g2_cascade_\ : std_logic;
signal \this_vga_signals.g0_4\ : std_logic;
signal \this_vga_signals.g1_0_0\ : std_logic;
signal \this_vga_signals.if_m1_0_cascade_\ : std_logic;
signal \this_vga_signals.N_129_i\ : std_logic;
signal \this_vga_signals.if_m1_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.g0_3_0_a3\ : std_logic;
signal \this_vga_signals.g1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_1_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x4_7_0_0\ : std_logic;
signal \this_vga_signals.g0_9_N_2L1_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x4_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_1_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_9_N_3L3\ : std_logic;
signal \this_vga_signals.g0_i_a4_4_0_0\ : std_logic;
signal \N_1422_0\ : std_logic;
signal \M_this_state_d_0_sqmuxa_2_cascade_\ : std_logic;
signal \M_this_state_d_0_sqmuxa_2\ : std_logic;
signal \this_start_data_delay.N_65_cascade_\ : std_logic;
signal \this_start_data_delay.N_42_0\ : std_logic;
signal \this_start_data_delay.N_43_0\ : std_logic;
signal dma_0 : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_0_2_cascade_\ : std_logic;
signal this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3 : std_logic;
signal \this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0\ : std_logic;
signal \this_vga_signals.if_m2\ : std_logic;
signal \this_vga_signals.if_m1_9_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m2_3_1\ : std_logic;
signal \this_vga_signals.if_i4_mux\ : std_logic;
signal \this_vga_signals.g0_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_a1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_0_2_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_0_2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb2_0_cascade_\ : std_logic;
signal this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d : std_logic;
signal \this_vga_signals.g2_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2\ : std_logic;
signal \this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb1_i_0\ : std_logic;
signal \this_vga_signals.N_4_2_cascade_\ : std_logic;
signal \this_vga_signals.if_m1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_d_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb2_0\ : std_logic;
signal this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1 : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb1_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_4_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.N_4_3_0_cascade_\ : std_logic;
signal \this_vga_signals.N_14_0\ : std_logic;
signal \this_vga_signals.g1\ : std_logic;
signal \this_vga_signals.g0_10_1\ : std_logic;
signal \this_vga_signals.N_24_mux\ : std_logic;
signal \this_vga_signals.g1_2\ : std_logic;
signal \this_vga_signals.g0_3_0_a3_3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals.if_N_9_i\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i\ : std_logic;
signal \this_vga_signals.SUM_2_0_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_1_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0\ : std_logic;
signal \this_vga_signals.g2_4\ : std_logic;
signal \this_vga_signals.m12_0_1\ : std_logic;
signal \this_start_data_delay.N_400\ : std_logic;
signal led23 : std_logic;
signal \this_start_data_delay.dmalto4_0_a2Z0Z_1\ : std_logic;
signal \this_start_data_delay.N_115\ : std_logic;
signal \this_start_data_delay.N_69\ : std_logic;
signal port_address_in_5 : std_logic;
signal port_address_in_6 : std_logic;
signal \this_start_data_delay.N_47_0_cascade_\ : std_logic;
signal \this_start_data_delay.N_48_0_cascade_\ : std_logic;
signal \N_28_0\ : std_logic;
signal \this_start_data_delay.N_82\ : std_logic;
signal \this_start_data_delay.N_82_cascade_\ : std_logic;
signal \M_this_substate_qZ0\ : std_logic;
signal \this_vga_signals.g0_0_x4_0_0\ : std_logic;
signal \this_vga_signals.vaddress_c2_cascade_\ : std_logic;
signal \this_vga_signals.N_5_2_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_5_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_1_1_cascade_\ : std_logic;
signal \this_vga_signals.N_3_2\ : std_logic;
signal \this_vga_signals.g0_1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.g0_5_2_0\ : std_logic;
signal \this_vga_signals.g2_1_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_2_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_0_a4\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_0_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_602_ns\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_4_x1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_2\ : std_logic;
signal \this_vga_signals.i1_mux\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc1_0\ : std_logic;
signal \this_vga_signals.vaddress_6\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_4_x0\ : std_logic;
signal \this_vga_signals.g1_7\ : std_logic;
signal \this_vga_signals.vaddress_3_6\ : std_logic;
signal \this_ppu.un3_sprites_addr_axb_0\ : std_logic;
signal \M_this_ppu_vram_addr_0\ : std_logic;
signal \M_this_ppu_sprites_addr_0\ : std_logic;
signal \M_this_state_qZ0Z_15\ : std_logic;
signal \M_this_state_qZ0Z_14\ : std_logic;
signal \M_this_state_qZ0Z_13\ : std_logic;
signal \this_start_data_delay.N_112_0\ : std_logic;
signal \this_start_data_delay.N_80_0\ : std_logic;
signal \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_aZ0Z2_cascade_\ : std_logic;
signal \this_start_data_delay.N_76_1\ : std_logic;
signal \this_start_data_delay.N_127_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_11\ : std_logic;
signal \this_start_data_delay.N_844_0_cascade_\ : std_logic;
signal \this_start_data_delay.N_151_cascade_\ : std_logic;
signal \this_start_data_delay.N_89_0\ : std_logic;
signal \M_this_state_qZ0Z_16\ : std_logic;
signal \this_start_data_delay.N_47_0\ : std_logic;
signal \this_start_data_delay.N_909_0_cascade_\ : std_logic;
signal led_c_1 : std_logic;
signal \this_start_data_delay.M_this_state_q_ns_0_i_0_0\ : std_logic;
signal \this_start_data_delay.M_this_state_q_ns_0_i_2_0_0\ : std_logic;
signal \N_822_0\ : std_logic;
signal \this_start_data_delay.N_910_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_10\ : std_logic;
signal \this_start_data_delay.N_90_0\ : std_logic;
signal port_address_in_1 : std_logic;
signal port_address_in_0 : std_logic;
signal port_address_in_2 : std_logic;
signal \this_start_data_delay.N_48_0\ : std_logic;
signal \this_start_data_delay.N_71\ : std_logic;
signal \this_start_data_delay.N_67\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_2_1_0\ : std_logic;
signal \this_vga_signals.N_4558_0\ : std_logic;
signal \this_vga_signals.g0_4_i_a3_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_4_i_1_cascade_\ : std_logic;
signal \this_vga_signals.N_6_2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_602_x0\ : std_logic;
signal \this_vga_signals.vaddress_c2\ : std_logic;
signal \this_vga_signals.r_N_4_mux\ : std_logic;
signal \this_vga_signals.r_N_4_mux_cascade_\ : std_logic;
signal \this_vga_signals.SUM_2\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a1_x1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a1_ns\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a1_x0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_602_x1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_3_x1\ : std_logic;
signal \this_vga_signals.N_4_0\ : std_logic;
signal \this_vga_signals.g0_6_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3\ : std_logic;
signal \this_vga_signals.N_4_0_0_1\ : std_logic;
signal \this_vga_signals.vaddress_0_5\ : std_logic;
signal \this_vga_signals.vaddress_0_6_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_5_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_repZ0Z1\ : std_logic;
signal \this_vga_signals.vaddress_5\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i\ : std_logic;
signal \this_vga_signals.g2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_2\ : std_logic;
signal \this_vga_signals.g0_i_x4_0_0\ : std_logic;
signal \this_vga_signals.g0_3_0_a3_1\ : std_logic;
signal \this_vga_signals.vaddress_1_6\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_0_c_RNIRLAZ0Z8\ : std_logic;
signal \M_this_ppu_vram_addr_1\ : std_logic;
signal \M_this_ppu_sprites_addr_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_1\ : std_logic;
signal \M_this_state_qZ0Z_12\ : std_logic;
signal \this_start_data_delay.N_125\ : std_logic;
signal \this_start_data_delay.un30_0_0_cascade_\ : std_logic;
signal \N_554_0_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_2\ : std_logic;
signal \this_start_data_delay.N_109_cascade_\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_4\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_3\ : std_logic;
signal \this_start_data_delay.M_last_qZ0\ : std_logic;
signal port_enb_c : std_logic;
signal \M_this_delay_clk_out_0\ : std_logic;
signal \this_start_data_delay.N_91_0_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_1\ : std_logic;
signal \this_start_data_delay.N_110_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_4\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_1\ : std_logic;
signal \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\ : std_logic;
signal \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\ : std_logic;
signal \M_this_ppu_vram_data_1\ : std_logic;
signal \this_start_data_delay.M_this_state_q_ns_0_i_2_0\ : std_logic;
signal \this_vga_signals_M_hcounter_d7_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \bfn_21_20_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_1\ : std_logic;
signal \G_442\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7\ : std_logic;
signal \bfn_21_21_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\ : std_logic;
signal \this_vga_signals.N_4557_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.M_vcounter_q_8_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_7_repZ0Z1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_601\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.N_1090_0\ : std_logic;
signal \this_vga_signals.N_1358_g\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.m58_1\ : std_logic;
signal \this_vga_signals.m58_0\ : std_logic;
signal \this_vga_signals.m58_4_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_6\ : std_logic;
signal this_vga_signals_vsync_1_i : std_logic;
signal \M_this_state_qZ0Z_3\ : std_logic;
signal \this_start_data_delay.N_123_cascade_\ : std_logic;
signal \N_812_0\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_7\ : std_logic;
signal \this_start_data_delay.N_129_cascade_\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_12_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_8\ : std_logic;
signal \this_start_data_delay.N_821_0_cascade_\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_11\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_10_cascade_\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_1\ : std_logic;
signal \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\ : std_logic;
signal \this_start_data_delay.N_55_0\ : std_logic;
signal \this_start_data_delay.N_84\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_2_cascade_\ : std_logic;
signal \this_start_data_delay.N_913_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_9\ : std_logic;
signal \M_this_state_qZ0Z_7\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_3_cascade_\ : std_logic;
signal \M_this_map_ram_read_data_7\ : std_logic;
signal \this_ppu.un10_sprites_addr_cry_4_c_RNIUV9BZ0\ : std_logic;
signal \this_start_data_delay.N_91_0\ : std_logic;
signal \this_start_data_delay.N_149_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_6\ : std_logic;
signal \this_start_data_delay.N_555_0\ : std_logic;
signal \this_start_data_delay.M_this_data_count_qlde_i_a3_0\ : std_logic;
signal \this_start_data_delay.M_this_data_count_qlde_i_2_tz_0\ : std_logic;
signal \this_start_data_delay.N_820_0_cascade_\ : std_logic;
signal \this_start_data_delay.N_151\ : std_logic;
signal \this_start_data_delay.N_820_0\ : std_logic;
signal \this_start_data_delay.M_this_data_count_qlde_i_1_cascade_\ : std_logic;
signal \this_start_data_delay.N_68\ : std_logic;
signal \M_this_state_qZ0Z_5\ : std_logic;
signal \N_554_0\ : std_logic;
signal \this_start_data_delay_M_this_data_count_q_3_0_a3_0_6_cascade_\ : std_logic;
signal \N_911\ : std_logic;
signal \M_this_data_count_q_3_0_13\ : std_logic;
signal \this_start_data_delay.N_93_0\ : std_logic;
signal \this_start_data_delay.N_122\ : std_logic;
signal \this_start_data_delay.N_149\ : std_logic;
signal \this_start_data_delay.N_121\ : std_logic;
signal \this_start_data_delay.N_938_0\ : std_logic;
signal \N_813_0\ : std_logic;
signal port_data_c_5 : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_6_cascade_\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_1_cascade_\ : std_logic;
signal \this_start_data_delay.N_993\ : std_logic;
signal \this_start_data_delay.N_109\ : std_logic;
signal \bfn_23_17_0_\ : std_logic;
signal \M_this_sprites_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_0_THRU_CO\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_1_THRU_CO\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_1\ : std_logic;
signal \M_this_sprites_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_2_THRU_CO\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_2\ : std_logic;
signal \M_this_sprites_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_3_THRU_CO\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_3\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_4\ : std_logic;
signal \M_this_sprites_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_5_THRU_CO\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_5\ : std_logic;
signal \M_this_sprites_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_6_THRU_CO\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_6\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_7\ : std_logic;
signal \bfn_23_18_0_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_8\ : std_logic;
signal \M_this_sprites_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_9_THRU_CO\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_9\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_10_THRU_CO\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_10\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_11_THRU_CO\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_11\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_13\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_12\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_0\ : std_logic;
signal un30_0 : std_logic;
signal \M_this_sprites_address_qZ0Z_0\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_9\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_8_THRU_CO\ : std_logic;
signal \M_this_sprites_address_qZ0Z_9\ : std_logic;
signal \this_start_data_delay.N_86_0\ : std_logic;
signal \M_this_reset_cond_out_g_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_3\ : std_logic;
signal \N_10_0\ : std_logic;
signal \this_start_data_delay.M_this_state_d62Z0Z_11\ : std_logic;
signal \this_start_data_delay.M_this_state_d62Z0Z_10\ : std_logic;
signal \this_start_data_delay.M_this_state_d62Z0Z_9_cascade_\ : std_logic;
signal \this_start_data_delay.M_this_state_d62Z0Z_8\ : std_logic;
signal \this_start_data_delay.M_this_state_dZ0Z62\ : std_logic;
signal \M_this_data_count_q_3_10\ : std_logic;
signal \this_start_data_delay_M_this_external_address_q_3_i_0_15\ : std_logic;
signal \N_116\ : std_logic;
signal \M_this_external_address_q_3_0_13\ : std_logic;
signal \M_this_map_ram_read_data_0\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_5_c_RNI55GZ0Z8\ : std_logic;
signal \M_this_ppu_sprites_addr_6\ : std_logic;
signal \this_sprites_ram.mem_WE_10\ : std_logic;
signal \this_sprites_ram.mem_WE_8\ : std_logic;
signal \this_sprites_ram.mem_WE_12\ : std_logic;
signal \this_sprites_ram.mem_WE_14\ : std_logic;
signal \N_811_0\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_5\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_4_THRU_CO\ : std_logic;
signal \M_this_sprites_address_qZ0Z_5\ : std_logic;
signal \this_sprites_ram.mem_WE_6\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_0\ : std_logic;
signal \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\ : std_logic;
signal port_data_c_0 : std_logic;
signal port_data_c_4 : std_logic;
signal port_data_c_6 : std_logic;
signal \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_3Z0Z_0_cascade_\ : std_logic;
signal \this_start_data_delay.N_902_0\ : std_logic;
signal \this_start_data_delay.N_821_0\ : std_logic;
signal port_data_c_7 : std_logic;
signal \this_start_data_delay.N_123\ : std_logic;
signal \N_41_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_3\ : std_logic;
signal \this_start_data_delay.N_992\ : std_logic;
signal \this_start_data_delay.N_110\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_7_THRU_CO\ : std_logic;
signal \this_start_data_delay.M_this_sprites_address_q_0_0_0_8_cascade_\ : std_logic;
signal \this_start_data_delay.N_990\ : std_logic;
signal \M_this_sprites_address_qZ0Z_8\ : std_logic;
signal \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\ : std_logic;
signal \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\ : std_logic;
signal \M_this_ppu_vram_data_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_0\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_12\ : std_logic;
signal \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0\ : std_logic;
signal \this_sprites_ram.mem_mem_2_0_RNINE6PZ0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_11\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_2\ : std_logic;
signal \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0\ : std_logic;
signal \this_sprites_ram.mem_WE_4\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_0\ : std_logic;
signal \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\ : std_logic;
signal \M_this_data_count_qZ0Z_0\ : std_logic;
signal \bfn_24_21_0_\ : std_logic;
signal \M_this_data_count_qZ0Z_1\ : std_logic;
signal \M_this_data_count_q_cry_0_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_0\ : std_logic;
signal \M_this_data_count_qZ0Z_2\ : std_logic;
signal \M_this_data_count_q_cry_1_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_1\ : std_logic;
signal \M_this_data_count_qZ0Z_3\ : std_logic;
signal \M_this_data_count_q_cry_2_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_2\ : std_logic;
signal \M_this_data_count_q_cry_3\ : std_logic;
signal \M_this_data_count_qZ0Z_5\ : std_logic;
signal \M_this_data_count_q_cry_4_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_4\ : std_logic;
signal \M_this_data_count_qZ0Z_6\ : std_logic;
signal \M_this_data_count_q_s_6\ : std_logic;
signal \M_this_data_count_q_cry_5\ : std_logic;
signal \M_this_data_count_qZ0Z_7\ : std_logic;
signal \M_this_data_count_q_cry_6_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_6\ : std_logic;
signal \M_this_data_count_q_cry_7\ : std_logic;
signal \M_this_data_count_qZ0Z_8\ : std_logic;
signal \M_this_data_count_q_s_8\ : std_logic;
signal \bfn_24_22_0_\ : std_logic;
signal \M_this_data_count_qZ0Z_9\ : std_logic;
signal \M_this_data_count_q_s_9\ : std_logic;
signal \M_this_data_count_q_cry_8\ : std_logic;
signal \M_this_data_count_qZ0Z_10\ : std_logic;
signal \M_this_data_count_q_cry_9_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_9\ : std_logic;
signal \M_this_data_count_qZ0Z_11\ : std_logic;
signal \M_this_data_count_q_s_11\ : std_logic;
signal \M_this_data_count_q_cry_10\ : std_logic;
signal \M_this_data_count_qZ0Z_12\ : std_logic;
signal \M_this_data_count_q_s_12\ : std_logic;
signal \M_this_data_count_q_cry_11\ : std_logic;
signal \M_this_data_count_qZ0Z_13\ : std_logic;
signal \M_this_data_count_q_cry_12_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_12\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \M_this_data_count_qZ0Z_14\ : std_logic;
signal \M_this_data_count_q_s_14\ : std_logic;
signal \M_this_data_count_q_cry_13\ : std_logic;
signal \M_this_data_count_qZ0Z_15\ : std_logic;
signal \M_this_data_count_q_cry_14\ : std_logic;
signal \M_this_data_count_q_s_15\ : std_logic;
signal \M_this_data_count_q_cry_3_THRU_CO\ : std_logic;
signal \N_33\ : std_logic;
signal \M_this_data_count_qZ0Z_4\ : std_logic;
signal \N_35\ : std_logic;
signal \M_this_external_address_q_3_0_12\ : std_logic;
signal \M_this_external_address_q_3_14\ : std_logic;
signal port_data_c_1 : std_logic;
signal \this_sprites_ram.mem_WE_2\ : std_logic;
signal \M_this_sprites_ram_write_en_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_12\ : std_logic;
signal \M_this_sprites_address_qZ0Z_11\ : std_logic;
signal \M_this_sprites_address_qZ0Z_13\ : std_logic;
signal \this_sprites_ram.mem_WE_0\ : std_logic;
signal \M_this_map_ram_read_data_4\ : std_logic;
signal \this_ppu.un10_sprites_addr_cry_1_c_RNIOM6BZ0\ : std_logic;
signal \M_this_ppu_sprites_addr_10\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_2\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_4_c_RNI32FZ0Z8\ : std_logic;
signal \M_this_ppu_sprites_addr_5\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_3\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_13\ : std_logic;
signal \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\ : std_logic;
signal \M_this_external_address_qZ0Z_0\ : std_logic;
signal \bfn_26_23_0_\ : std_logic;
signal \M_this_external_address_qZ0Z_1\ : std_logic;
signal \M_this_external_address_q_cry_0\ : std_logic;
signal \M_this_external_address_qZ0Z_2\ : std_logic;
signal \M_this_external_address_q_cry_1\ : std_logic;
signal \M_this_external_address_qZ0Z_3\ : std_logic;
signal \M_this_external_address_q_cry_2\ : std_logic;
signal \M_this_external_address_qZ0Z_4\ : std_logic;
signal \M_this_external_address_q_cry_3\ : std_logic;
signal \M_this_external_address_qZ0Z_5\ : std_logic;
signal \M_this_external_address_q_cry_4\ : std_logic;
signal \M_this_external_address_qZ0Z_6\ : std_logic;
signal \M_this_external_address_q_cry_5\ : std_logic;
signal \M_this_external_address_qZ0Z_7\ : std_logic;
signal \M_this_external_address_q_cry_6\ : std_logic;
signal \M_this_external_address_q_cry_7\ : std_logic;
signal \M_this_external_address_qZ0Z_8\ : std_logic;
signal \M_this_external_address_q_s_8\ : std_logic;
signal \bfn_26_24_0_\ : std_logic;
signal \M_this_external_address_qZ0Z_9\ : std_logic;
signal \M_this_external_address_q_s_9\ : std_logic;
signal \M_this_external_address_q_cry_8\ : std_logic;
signal \M_this_external_address_q_cry_9\ : std_logic;
signal \M_this_external_address_q_cry_10\ : std_logic;
signal \M_this_external_address_qZ0Z_12\ : std_logic;
signal \M_this_external_address_q_cry_11_THRU_CO\ : std_logic;
signal \M_this_external_address_q_cry_11\ : std_logic;
signal \M_this_external_address_qZ0Z_13\ : std_logic;
signal \M_this_external_address_q_cry_12_THRU_CO\ : std_logic;
signal \M_this_external_address_q_cry_12\ : std_logic;
signal \M_this_external_address_qZ0Z_14\ : std_logic;
signal \M_this_external_address_q_cry_13_THRU_CO\ : std_logic;
signal \M_this_external_address_q_cry_13\ : std_logic;
signal \M_this_external_address_qZ0Z_15\ : std_logic;
signal \M_this_external_address_q_cry_14\ : std_logic;
signal \M_this_external_address_q_s_15\ : std_logic;
signal \M_this_external_address_q_s_11\ : std_logic;
signal port_data_c_3 : std_logic;
signal \M_this_external_address_qZ0Z_11\ : std_logic;
signal \M_this_external_address_q_s_10\ : std_logic;
signal \M_this_external_address_d_1_sqmuxa\ : std_logic;
signal port_data_c_2 : std_logic;
signal \N_39\ : std_logic;
signal \M_this_external_address_qZ0Z_10\ : std_logic;
signal clk_0_c_g : std_logic;
signal \N_37\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_1\ : std_logic;
signal \this_ppu.M_state_qZ0Z_3\ : std_logic;
signal \this_ppu.M_state_qZ0Z_2\ : std_logic;
signal \this_ppu.un3_sprites_addr_cry_3_c_RNI1VDZ0Z8\ : std_logic;
signal \M_this_ppu_sprites_addr_4\ : std_logic;
signal port_address_in_7 : std_logic;
signal port_address_in_4 : std_logic;
signal port_rw_in : std_logic;
signal port_address_in_3 : std_logic;
signal \this_start_data_delay.un1_M_this_state_q_17_i_o2_1Z0Z_4\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic_vector(1 downto 0);
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal led_wire : std_logic_vector(7 downto 0);
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_map_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    led <= led_wire;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \M_this_map_ram_read_data_3\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_2\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_1\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_0\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&\N__13431\&\N__13662\&\N__16782\&\N__16638\&\N__16701\&\N__12840\&\N__12891\&\N__13584\&\N__13827\&\N__13962\;
    \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&\N__11931\&\N__11964\&\N__11994\&\N__11589\&\N__11619\&\N__11649\&\N__11679\&\N__11709\&\N__11739\&\N__11766\;
    \this_map_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&\N__13689\&'0'&'0'&'0'&\N__11796\&'0'&'0'&'0'&\N__15012\&'0'&'0'&'0'&\N__12633\&'0';
    \M_this_map_ram_read_data_7\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_6\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_5\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_4\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&\N__13425\&\N__13656\&\N__16776\&\N__16632\&\N__16695\&\N__12834\&\N__12885\&\N__13578\&\N__13821\&\N__13956\;
    \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&\N__11925\&\N__11958\&\N__11988\&\N__11583\&\N__11613\&\N__11643\&\N__11673\&\N__11703\&\N__11733\&\N__11760\;
    \this_map_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&\N__12405\&'0'&'0'&'0'&\N__11826\&'0'&'0'&'0'&\N__13410\&'0'&'0'&'0'&\N__13677\&'0';
    \M_this_oam_ram_read_data_13\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \this_oam_ram.M_this_oam_ram_read_data_12\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(12);
    \this_oam_ram.M_this_oam_ram_read_data_11\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_oam_ram.M_this_oam_ram_read_data_10\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(10);
    \this_oam_ram.M_this_oam_ram_read_data_9\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_oam_ram_read_data_8\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(8);
    \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__11211\&\N__11241\&\N__11010\&\N__11037\&\N__11067\&\N__11094\;
    \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ <= \N__11301\&\N__11289\&\N__11385\&\N__12258\&\N__11247\&\N__14709\&\N__12039\&\N__11259\&\N__11253\&\N__12018\&\N__11268\&\N__11394\&\N__12030\&\N__12006\&\N__11280\&\N__11559\;
    \M_this_oam_ram_read_data_23\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(7);
    \this_oam_ram.M_this_oam_ram_read_data_22\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(6);
    \this_oam_ram.M_this_oam_ram_read_data_21\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \this_oam_ram.M_this_oam_ram_read_data_20\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(4);
    \this_oam_ram.M_this_oam_ram_read_data_19\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_oam_ram.M_this_oam_ram_read_data_18\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(2);
    \this_oam_ram.M_this_oam_ram_read_data_17\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_16\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__11205\&\N__11235\&\N__11004\&\N__11031\&\N__11061\&\N__11088\;
    \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ <= \N__11340\&\N__12801\&\N__12270\&\N__11355\&\N__11376\&\N__11172\&\N__12249\&\N__12237\&\N__11160\&\N__12225\&\N__12213\&\N__11166\&\N__11349\&\N__12855\&\N__12921\&\N__12786\;
    \this_sprites_ram.mem_out_bus0_1\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_0\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ <= \N__30390\&\N__15570\&\N__15291\&\N__12162\&\N__26661\&\N__30234\&\N__31791\&\N__15714\&\N__14121\&\N__20877\&\N__19251\;
    \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ <= \N__25539\&\N__26409\&\N__27483\&\N__25689\&\N__25824\&\N__27174\&\N__24852\&\N__24996\&\N__25137\&\N__25272\&\N__26559\;
    \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22134\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24584\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus0_3\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_2\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ <= \N__30384\&\N__15564\&\N__15285\&\N__12156\&\N__26655\&\N__30228\&\N__31785\&\N__15708\&\N__14115\&\N__20871\&\N__19245\;
    \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ <= \N__25533\&\N__26403\&\N__27477\&\N__25683\&\N__25818\&\N__27168\&\N__24846\&\N__24990\&\N__25131\&\N__25266\&\N__26553\;
    \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27803\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__27246\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_1\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_0\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ <= \N__30378\&\N__15558\&\N__15279\&\N__12150\&\N__26649\&\N__30222\&\N__31779\&\N__15702\&\N__14109\&\N__20865\&\N__19239\;
    \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ <= \N__25527\&\N__26397\&\N__27471\&\N__25677\&\N__25812\&\N__27162\&\N__24840\&\N__24984\&\N__25125\&\N__25260\&\N__26547\;
    \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22129\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24576\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_3\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_2\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ <= \N__30372\&\N__15552\&\N__15273\&\N__12144\&\N__26643\&\N__30216\&\N__31773\&\N__15696\&\N__14103\&\N__20859\&\N__19233\;
    \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ <= \N__25521\&\N__26391\&\N__27465\&\N__25671\&\N__25806\&\N__27156\&\N__24834\&\N__24978\&\N__25119\&\N__25254\&\N__26541\;
    \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27795\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__27233\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_1\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_0\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ <= \N__30366\&\N__15546\&\N__15267\&\N__12138\&\N__26637\&\N__30210\&\N__31767\&\N__15690\&\N__14097\&\N__20853\&\N__19227\;
    \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ <= \N__25515\&\N__26385\&\N__27459\&\N__25665\&\N__25800\&\N__27150\&\N__24828\&\N__24972\&\N__25113\&\N__25248\&\N__26535\;
    \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22118\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24562\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_3\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_2\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ <= \N__30360\&\N__15540\&\N__15261\&\N__12132\&\N__26631\&\N__30204\&\N__31761\&\N__15684\&\N__14091\&\N__20847\&\N__19221\;
    \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ <= \N__25509\&\N__26379\&\N__27453\&\N__25659\&\N__25794\&\N__27144\&\N__24822\&\N__24966\&\N__25107\&\N__25242\&\N__26529\;
    \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27781\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__27218\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_1\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_0\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ <= \N__30354\&\N__15534\&\N__15255\&\N__12126\&\N__26625\&\N__30198\&\N__31755\&\N__15678\&\N__14085\&\N__20841\&\N__19215\;
    \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ <= \N__25503\&\N__26373\&\N__27447\&\N__25653\&\N__25788\&\N__27138\&\N__24816\&\N__24960\&\N__25101\&\N__25236\&\N__26523\;
    \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22092\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24544\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_3\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_2\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ <= \N__30348\&\N__15528\&\N__15249\&\N__12120\&\N__26619\&\N__30192\&\N__31749\&\N__15672\&\N__14079\&\N__20835\&\N__19209\;
    \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ <= \N__25497\&\N__26367\&\N__27441\&\N__25647\&\N__25782\&\N__27132\&\N__24810\&\N__24954\&\N__25095\&\N__25230\&\N__26517\;
    \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27763\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__27204\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_1\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_0\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ <= \N__30342\&\N__15522\&\N__15243\&\N__12114\&\N__26613\&\N__30186\&\N__31743\&\N__15666\&\N__14073\&\N__20829\&\N__19203\;
    \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ <= \N__25491\&\N__26361\&\N__27435\&\N__25641\&\N__25776\&\N__27126\&\N__24804\&\N__24948\&\N__25089\&\N__25224\&\N__26511\;
    \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22093\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24553\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_3\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_2\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ <= \N__30336\&\N__15516\&\N__15237\&\N__12108\&\N__26607\&\N__30180\&\N__31737\&\N__15660\&\N__14067\&\N__20823\&\N__19197\;
    \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ <= \N__25485\&\N__26355\&\N__27429\&\N__25635\&\N__25770\&\N__27120\&\N__24798\&\N__24942\&\N__25083\&\N__25218\&\N__26505\;
    \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27772\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__27237\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_1\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_0\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ <= \N__30330\&\N__15510\&\N__15231\&\N__12102\&\N__26601\&\N__30174\&\N__31731\&\N__15654\&\N__14061\&\N__20817\&\N__19191\;
    \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ <= \N__25479\&\N__26349\&\N__27423\&\N__25629\&\N__25764\&\N__27114\&\N__24792\&\N__24936\&\N__25077\&\N__25212\&\N__26499\;
    \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22111\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24569\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_3\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_2\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ <= \N__30324\&\N__15504\&\N__15225\&\N__12096\&\N__26595\&\N__30168\&\N__31725\&\N__15648\&\N__14055\&\N__20811\&\N__19185\;
    \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ <= \N__25473\&\N__26343\&\N__27417\&\N__25623\&\N__25758\&\N__27108\&\N__24786\&\N__24930\&\N__25071\&\N__25206\&\N__26493\;
    \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27788\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__27247\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_1\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_0\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ <= \N__30318\&\N__15498\&\N__15219\&\N__12090\&\N__26589\&\N__30162\&\N__31719\&\N__15642\&\N__14049\&\N__20805\&\N__19179\;
    \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ <= \N__25467\&\N__26337\&\N__27411\&\N__25617\&\N__25752\&\N__27102\&\N__24780\&\N__24924\&\N__25065\&\N__25200\&\N__26487\;
    \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22125\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24580\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_3\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_2\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ <= \N__30312\&\N__15492\&\N__15213\&\N__12084\&\N__26583\&\N__30156\&\N__31713\&\N__15636\&\N__14043\&\N__20799\&\N__19173\;
    \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ <= \N__25461\&\N__26331\&\N__27405\&\N__25611\&\N__25746\&\N__27096\&\N__24774\&\N__24918\&\N__25059\&\N__25194\&\N__26481\;
    \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27799\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__27254\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_1\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_0\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ <= \N__30306\&\N__15486\&\N__15207\&\N__12078\&\N__26577\&\N__30150\&\N__31707\&\N__15630\&\N__14037\&\N__20793\&\N__19167\;
    \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ <= \N__25455\&\N__26325\&\N__27399\&\N__25605\&\N__25740\&\N__27090\&\N__24768\&\N__24912\&\N__25053\&\N__25188\&\N__26475\;
    \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22133\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24585\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_3\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_2\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ <= \N__30300\&\N__15480\&\N__15201\&\N__12072\&\N__26571\&\N__30144\&\N__31701\&\N__15624\&\N__14031\&\N__20787\&\N__19161\;
    \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ <= \N__25449\&\N__26319\&\N__27393\&\N__25599\&\N__25734\&\N__27084\&\N__24762\&\N__24906\&\N__25047\&\N__25182\&\N__26469\;
    \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27804\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__27258\&'0'&'0'&'0';
    \M_this_vram_read_data_3\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_vram_read_data_2\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_vram_read_data_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_vram_read_data_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__17046\&\N__13323\&\N__11820\&\N__12195\&\N__13344\&\N__11805\&\N__11463\&\N__13197\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__16848\&\N__13623\&\N__13577\&\N__13820\&\N__13952\&\N__13890\&\N__20940\&\N__19335\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28790\&\N__17190\&\N__21162\&\N__14685\;

    \this_map_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32649\,
            RE => \N__29819\,
            WCLKE => \N__19898\,
            WCLK => \N__32650\,
            WE => \N__29837\
        );

    \this_map_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32655\,
            RE => \N__29841\,
            WCLKE => \N__19899\,
            WCLK => \N__32656\,
            WE => \N__29836\
        );

    \this_oam_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32605\,
            RE => \N__29755\,
            WCLKE => \N__18621\,
            WCLK => \N__32606\,
            WE => \N__29794\
        );

    \this_oam_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32621\,
            RE => \N__29790\,
            WCLKE => \N__18622\,
            WCLK => \N__32622\,
            WE => \N__29795\
        );

    \this_sprites_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32524\,
            RE => \N__29789\,
            WCLKE => \N__27282\,
            WCLK => \N__32525\,
            WE => \N__29787\
        );

    \this_sprites_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32526\,
            RE => \N__29788\,
            WCLKE => \N__27278\,
            WCLK => \N__32527\,
            WE => \N__29511\
        );

    \this_sprites_ram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32528\,
            RE => \N__29744\,
            WCLKE => \N__27303\,
            WCLK => \N__32529\,
            WE => \N__29739\
        );

    \this_sprites_ram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32532\,
            RE => \N__29743\,
            WCLKE => \N__27299\,
            WCLK => \N__32533\,
            WE => \N__29735\
        );

    \this_sprites_ram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32540\,
            RE => \N__29651\,
            WCLKE => \N__27348\,
            WCLK => \N__32539\,
            WE => \N__29664\
        );

    \this_sprites_ram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32558\,
            RE => \N__29650\,
            WCLKE => \N__27347\,
            WCLK => \N__32559\,
            WE => \N__29510\
        );

    \this_sprites_ram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32578\,
            RE => \N__29513\,
            WCLKE => \N__27326\,
            WCLK => \N__32579\,
            WE => \N__29539\
        );

    \this_sprites_ram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32595\,
            RE => \N__29512\,
            WCLKE => \N__27327\,
            WCLK => \N__32596\,
            WE => \N__29426\
        );

    \this_sprites_ram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32614\,
            RE => \N__29514\,
            WCLKE => \N__27035\,
            WCLK => \N__32615\,
            WE => \N__29519\
        );

    \this_sprites_ram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32628\,
            RE => \N__29515\,
            WCLKE => \N__27042\,
            WCLK => \N__32629\,
            WE => \N__29520\
        );

    \this_sprites_ram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32634\,
            RE => \N__29702\,
            WCLKE => \N__28571\,
            WCLK => \N__32635\,
            WE => \N__29629\
        );

    \this_sprites_ram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32645\,
            RE => \N__29628\,
            WCLKE => \N__28572\,
            WCLK => \N__32646\,
            WE => \N__29630\
        );

    \this_sprites_ram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32652\,
            RE => \N__29754\,
            WCLKE => \N__30785\,
            WCLK => \N__32653\,
            WE => \N__29720\
        );

    \this_sprites_ram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32657\,
            RE => \N__29725\,
            WCLKE => \N__30786\,
            WCLK => \N__32658\,
            WE => \N__29721\
        );

    \this_sprites_ram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32661\,
            RE => \N__29779\,
            WCLKE => \N__30446\,
            WCLK => \N__32662\,
            WE => \N__29778\
        );

    \this_sprites_ram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32663\,
            RE => \N__29780\,
            WCLKE => \N__30447\,
            WCLK => \N__32664\,
            WE => \N__29812\
        );

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__32659\,
            RE => \N__29842\,
            WCLKE => \N__14010\,
            WCLK => \N__32660\,
            WE => \N__29844\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__33433\,
            GLOBALBUFFEROUTPUT => clk_0_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33435\,
            DIN => \N__33434\,
            DOUT => \N__33433\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__33435\,
            PADOUT => \N__33434\,
            PADIN => \N__33433\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33424\,
            DIN => \N__33423\,
            DOUT => \N__33422\,
            PACKAGEPIN => debug_wire(0)
        );

    \debug_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33424\,
            PADOUT => \N__33423\,
            PADIN => \N__33422\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33415\,
            DIN => \N__33414\,
            DOUT => \N__33413\,
            PACKAGEPIN => debug_wire(1)
        );

    \debug_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33415\,
            PADOUT => \N__33414\,
            PADIN => \N__33413\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33406\,
            DIN => \N__33405\,
            DOUT => \N__33404\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33406\,
            PADOUT => \N__33405\,
            PADIN => \N__33404\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13224\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33397\,
            DIN => \N__33396\,
            DOUT => \N__33395\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33397\,
            PADOUT => \N__33396\,
            PADIN => \N__33395\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13443\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33388\,
            DIN => \N__33387\,
            DOUT => \N__33386\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33388\,
            PADOUT => \N__33387\,
            PADIN => \N__33386\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__29835\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33379\,
            DIN => \N__33378\,
            DOUT => \N__33377\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33379\,
            PADOUT => \N__33378\,
            PADIN => \N__33377\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__19953\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33370\,
            DIN => \N__33369\,
            DOUT => \N__33368\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33370\,
            PADOUT => \N__33369\,
            PADIN => \N__33368\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33361\,
            DIN => \N__33360\,
            DOUT => \N__33359\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33361\,
            PADOUT => \N__33360\,
            PADIN => \N__33359\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33352\,
            DIN => \N__33351\,
            DOUT => \N__33350\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33352\,
            PADOUT => \N__33351\,
            PADIN => \N__33350\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33343\,
            DIN => \N__33342\,
            DOUT => \N__33341\,
            PACKAGEPIN => led_wire(5)
        );

    \led_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33343\,
            PADOUT => \N__33342\,
            PADIN => \N__33341\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33334\,
            DIN => \N__33333\,
            DOUT => \N__33332\,
            PACKAGEPIN => led_wire(6)
        );

    \led_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33334\,
            PADOUT => \N__33333\,
            PADIN => \N__33332\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33325\,
            DIN => \N__33324\,
            DOUT => \N__33323\,
            PACKAGEPIN => led_wire(7)
        );

    \led_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33325\,
            PADOUT => \N__33324\,
            PADIN => \N__33323\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33316\,
            DIN => \N__33315\,
            DOUT => \N__33314\,
            PACKAGEPIN => port_address(0)
        );

    \port_address_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33316\,
            PADOUT => \N__33315\,
            PADIN => \N__33314\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__31191\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16079\
        );

    \port_address_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33307\,
            DIN => \N__33306\,
            DOUT => \N__33305\,
            PACKAGEPIN => port_address(1)
        );

    \port_address_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33307\,
            PADOUT => \N__33306\,
            PADIN => \N__33305\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__31164\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16048\
        );

    \port_address_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33298\,
            DIN => \N__33297\,
            DOUT => \N__33296\,
            PACKAGEPIN => port_address(2)
        );

    \port_address_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33298\,
            PADOUT => \N__33297\,
            PADIN => \N__33296\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__31143\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16113\
        );

    \port_address_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33289\,
            DIN => \N__33288\,
            DOUT => \N__33287\,
            PACKAGEPIN => port_address(3)
        );

    \port_address_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33289\,
            PADOUT => \N__33288\,
            PADIN => \N__33287\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__31116\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16049\
        );

    \port_address_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33280\,
            DIN => \N__33279\,
            DOUT => \N__33278\,
            PACKAGEPIN => port_address(4)
        );

    \port_address_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33280\,
            PADOUT => \N__33279\,
            PADIN => \N__33278\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__31089\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16122\
        );

    \port_address_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33271\,
            DIN => \N__33270\,
            DOUT => \N__33269\,
            PACKAGEPIN => port_address(5)
        );

    \port_address_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33271\,
            PADOUT => \N__33270\,
            PADIN => \N__33269\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__31071\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16120\
        );

    \port_address_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33262\,
            DIN => \N__33261\,
            DOUT => \N__33260\,
            PACKAGEPIN => port_address(6)
        );

    \port_address_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33262\,
            PADOUT => \N__33261\,
            PADIN => \N__33260\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__31047\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16091\
        );

    \port_address_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33253\,
            DIN => \N__33252\,
            DOUT => \N__33251\,
            PACKAGEPIN => port_address(7)
        );

    \port_address_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33253\,
            PADOUT => \N__33252\,
            PADIN => \N__33251\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__31026\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16136\
        );

    \port_address_obuft_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33244\,
            DIN => \N__33243\,
            DOUT => \N__33242\,
            PACKAGEPIN => port_address(10)
        );

    \port_address_obuft_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33244\,
            PADOUT => \N__33243\,
            PADIN => \N__33242\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__32682\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16112\
        );

    \port_address_obuft_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33235\,
            DIN => \N__33234\,
            DOUT => \N__33233\,
            PACKAGEPIN => port_address(11)
        );

    \port_address_obuft_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33235\,
            PADOUT => \N__33234\,
            PADIN => \N__33233\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__31212\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16137\
        );

    \port_address_obuft_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33226\,
            DIN => \N__33225\,
            DOUT => \N__33224\,
            PACKAGEPIN => port_address(12)
        );

    \port_address_obuft_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33226\,
            PADOUT => \N__33225\,
            PADIN => \N__33224\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__31542\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16123\
        );

    \port_address_obuft_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33217\,
            DIN => \N__33216\,
            DOUT => \N__33215\,
            PACKAGEPIN => port_address(13)
        );

    \port_address_obuft_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33217\,
            PADOUT => \N__33216\,
            PADIN => \N__33215\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__31500\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16121\
        );

    \port_address_obuft_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33208\,
            DIN => \N__33207\,
            DOUT => \N__33206\,
            PACKAGEPIN => port_address(14)
        );

    \port_address_obuft_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33208\,
            PADOUT => \N__33207\,
            PADIN => \N__33206\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__31452\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16015\
        );

    \port_address_obuft_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33199\,
            DIN => \N__33198\,
            DOUT => \N__33197\,
            PACKAGEPIN => port_address(15)
        );

    \port_address_obuft_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33199\,
            PADOUT => \N__33198\,
            PADIN => \N__33197\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__31404\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16135\
        );

    \port_address_obuft_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33190\,
            DIN => \N__33189\,
            DOUT => \N__33188\,
            PACKAGEPIN => port_address(8)
        );

    \port_address_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33190\,
            PADOUT => \N__33189\,
            PADIN => \N__33188\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__30996\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16011\
        );

    \port_address_obuft_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33181\,
            DIN => \N__33180\,
            DOUT => \N__33179\,
            PACKAGEPIN => port_address(9)
        );

    \port_address_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33181\,
            PADOUT => \N__33180\,
            PADIN => \N__33179\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__31584\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16131\
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33172\,
            DIN => \N__33171\,
            DOUT => \N__33170\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__33172\,
            PADOUT => \N__33171\,
            PADIN => \N__33170\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33163\,
            DIN => \N__33162\,
            DOUT => \N__33161\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__33163\,
            PADOUT => \N__33162\,
            PADIN => \N__33161\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33154\,
            DIN => \N__33153\,
            DOUT => \N__33152\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__33154\,
            PADOUT => \N__33153\,
            PADIN => \N__33152\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33145\,
            DIN => \N__33144\,
            DOUT => \N__33143\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__33145\,
            PADOUT => \N__33144\,
            PADIN => \N__33143\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33136\,
            DIN => \N__33135\,
            DOUT => \N__33134\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__33136\,
            PADOUT => \N__33135\,
            PADIN => \N__33134\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33127\,
            DIN => \N__33126\,
            DOUT => \N__33125\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__33127\,
            PADOUT => \N__33126\,
            PADIN => \N__33125\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33118\,
            DIN => \N__33117\,
            DOUT => \N__33116\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__33118\,
            PADOUT => \N__33117\,
            PADIN => \N__33116\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33109\,
            DIN => \N__33108\,
            DOUT => \N__33107\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__33109\,
            PADOUT => \N__33108\,
            PADIN => \N__33107\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33100\,
            DIN => \N__33099\,
            DOUT => \N__33098\,
            PACKAGEPIN => port_data_wire(7)
        );

    \port_data_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__33100\,
            PADOUT => \N__33099\,
            PADIN => \N__33098\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33091\,
            DIN => \N__33090\,
            DOUT => \N__33089\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33091\,
            PADOUT => \N__33090\,
            PADIN => \N__33089\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__17298\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33082\,
            DIN => \N__33081\,
            DOUT => \N__33080\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33082\,
            PADOUT => \N__33081\,
            PADIN => \N__33080\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__17745\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33073\,
            DIN => \N__33072\,
            DOUT => \N__33071\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__33073\,
            PADOUT => \N__33072\,
            PADIN => \N__33071\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33064\,
            DIN => \N__33063\,
            DOUT => \N__33062\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33064\,
            PADOUT => \N__33063\,
            PADIN => \N__33062\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__10980\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33055\,
            DIN => \N__33054\,
            DOUT => \N__33053\,
            PACKAGEPIN => port_rw
        );

    \port_rw_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__33055\,
            PADOUT => \N__33054\,
            PADIN => \N__33053\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_in,
            DIN1 => OPEN,
            DOUT0 => \N__29843\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__16130\
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33046\,
            DIN => \N__33045\,
            DOUT => \N__33044\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33046\,
            PADOUT => \N__33045\,
            PADIN => \N__33044\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11154\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33037\,
            DIN => \N__33036\,
            DOUT => \N__33035\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33037\,
            PADOUT => \N__33036\,
            PADIN => \N__33035\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11475\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33028\,
            DIN => \N__33027\,
            DOUT => \N__33026\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33028\,
            PADOUT => \N__33027\,
            PADIN => \N__33026\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11124\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33019\,
            DIN => \N__33018\,
            DOUT => \N__33017\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33019\,
            PADOUT => \N__33018\,
            PADIN => \N__33017\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11328\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33010\,
            DIN => \N__33009\,
            DOUT => \N__33008\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33010\,
            PADOUT => \N__33009\,
            PADIN => \N__33008\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11316\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__33001\,
            DIN => \N__33000\,
            DOUT => \N__32999\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__33001\,
            PADOUT => \N__33000\,
            PADIN => \N__32999\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11835\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__32992\,
            DIN => \N__32991\,
            DOUT => \N__32990\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__32992\,
            PADOUT => \N__32991\,
            PADIN => \N__32990\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__32983\,
            DIN => \N__32982\,
            DOUT => \N__32981\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__32983\,
            PADOUT => \N__32982\,
            PADIN => \N__32981\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11139\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__32974\,
            DIN => \N__32973\,
            DOUT => \N__32972\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__32974\,
            PADOUT => \N__32973\,
            PADIN => \N__32972\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__22200\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__8133\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32952\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__32952\,
            I => \M_this_external_address_q_s_10\
        );

    \I__8131\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32945\
        );

    \I__8130\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32942\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__32945\,
            I => \N__32936\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__32942\,
            I => \N__32936\
        );

    \I__8127\ : InMux
    port map (
            O => \N__32941\,
            I => \N__32933\
        );

    \I__8126\ : Span4Mux_v
    port map (
            O => \N__32936\,
            I => \N__32927\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__32933\,
            I => \N__32927\
        );

    \I__8124\ : InMux
    port map (
            O => \N__32932\,
            I => \N__32924\
        );

    \I__8123\ : Odrv4
    port map (
            O => \N__32927\,
            I => \M_this_external_address_d_1_sqmuxa\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__32924\,
            I => \M_this_external_address_d_1_sqmuxa\
        );

    \I__8121\ : InMux
    port map (
            O => \N__32919\,
            I => \N__32916\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__32916\,
            I => \N__32912\
        );

    \I__8119\ : InMux
    port map (
            O => \N__32915\,
            I => \N__32909\
        );

    \I__8118\ : Span4Mux_v
    port map (
            O => \N__32912\,
            I => \N__32905\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__32909\,
            I => \N__32900\
        );

    \I__8116\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32897\
        );

    \I__8115\ : Span4Mux_h
    port map (
            O => \N__32905\,
            I => \N__32893\
        );

    \I__8114\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32888\
        );

    \I__8113\ : CascadeMux
    port map (
            O => \N__32903\,
            I => \N__32885\
        );

    \I__8112\ : Span4Mux_h
    port map (
            O => \N__32900\,
            I => \N__32879\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__32897\,
            I => \N__32879\
        );

    \I__8110\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32876\
        );

    \I__8109\ : Span4Mux_h
    port map (
            O => \N__32893\,
            I => \N__32871\
        );

    \I__8108\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32868\
        );

    \I__8107\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32865\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__32888\,
            I => \N__32862\
        );

    \I__8105\ : InMux
    port map (
            O => \N__32885\,
            I => \N__32859\
        );

    \I__8104\ : CascadeMux
    port map (
            O => \N__32884\,
            I => \N__32855\
        );

    \I__8103\ : Span4Mux_v
    port map (
            O => \N__32879\,
            I => \N__32850\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__32876\,
            I => \N__32850\
        );

    \I__8101\ : InMux
    port map (
            O => \N__32875\,
            I => \N__32845\
        );

    \I__8100\ : InMux
    port map (
            O => \N__32874\,
            I => \N__32845\
        );

    \I__8099\ : Span4Mux_h
    port map (
            O => \N__32871\,
            I => \N__32840\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__32868\,
            I => \N__32840\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__32865\,
            I => \N__32833\
        );

    \I__8096\ : Span4Mux_h
    port map (
            O => \N__32862\,
            I => \N__32833\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__32859\,
            I => \N__32833\
        );

    \I__8094\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32830\
        );

    \I__8093\ : InMux
    port map (
            O => \N__32855\,
            I => \N__32827\
        );

    \I__8092\ : Span4Mux_v
    port map (
            O => \N__32850\,
            I => \N__32823\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__32845\,
            I => \N__32820\
        );

    \I__8090\ : Span4Mux_h
    port map (
            O => \N__32840\,
            I => \N__32810\
        );

    \I__8089\ : Span4Mux_v
    port map (
            O => \N__32833\,
            I => \N__32810\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__32830\,
            I => \N__32810\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__32827\,
            I => \N__32810\
        );

    \I__8086\ : InMux
    port map (
            O => \N__32826\,
            I => \N__32807\
        );

    \I__8085\ : Span4Mux_h
    port map (
            O => \N__32823\,
            I => \N__32804\
        );

    \I__8084\ : Span4Mux_v
    port map (
            O => \N__32820\,
            I => \N__32801\
        );

    \I__8083\ : CascadeMux
    port map (
            O => \N__32819\,
            I => \N__32797\
        );

    \I__8082\ : Span4Mux_v
    port map (
            O => \N__32810\,
            I => \N__32794\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__32807\,
            I => \N__32791\
        );

    \I__8080\ : Span4Mux_h
    port map (
            O => \N__32804\,
            I => \N__32786\
        );

    \I__8079\ : Span4Mux_v
    port map (
            O => \N__32801\,
            I => \N__32786\
        );

    \I__8078\ : InMux
    port map (
            O => \N__32800\,
            I => \N__32783\
        );

    \I__8077\ : InMux
    port map (
            O => \N__32797\,
            I => \N__32780\
        );

    \I__8076\ : Span4Mux_h
    port map (
            O => \N__32794\,
            I => \N__32777\
        );

    \I__8075\ : Span12Mux_v
    port map (
            O => \N__32791\,
            I => \N__32768\
        );

    \I__8074\ : Sp12to4
    port map (
            O => \N__32786\,
            I => \N__32768\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__32783\,
            I => \N__32768\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__32780\,
            I => \N__32768\
        );

    \I__8071\ : Sp12to4
    port map (
            O => \N__32777\,
            I => \N__32763\
        );

    \I__8070\ : Span12Mux_h
    port map (
            O => \N__32768\,
            I => \N__32763\
        );

    \I__8069\ : Odrv12
    port map (
            O => \N__32763\,
            I => port_data_c_2
        );

    \I__8068\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32741\
        );

    \I__8067\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32741\
        );

    \I__8066\ : InMux
    port map (
            O => \N__32758\,
            I => \N__32741\
        );

    \I__8065\ : InMux
    port map (
            O => \N__32757\,
            I => \N__32736\
        );

    \I__8064\ : InMux
    port map (
            O => \N__32756\,
            I => \N__32736\
        );

    \I__8063\ : InMux
    port map (
            O => \N__32755\,
            I => \N__32724\
        );

    \I__8062\ : InMux
    port map (
            O => \N__32754\,
            I => \N__32724\
        );

    \I__8061\ : InMux
    port map (
            O => \N__32753\,
            I => \N__32724\
        );

    \I__8060\ : InMux
    port map (
            O => \N__32752\,
            I => \N__32724\
        );

    \I__8059\ : InMux
    port map (
            O => \N__32751\,
            I => \N__32715\
        );

    \I__8058\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32715\
        );

    \I__8057\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32715\
        );

    \I__8056\ : InMux
    port map (
            O => \N__32748\,
            I => \N__32715\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__32741\,
            I => \N__32712\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__32736\,
            I => \N__32709\
        );

    \I__8053\ : InMux
    port map (
            O => \N__32735\,
            I => \N__32702\
        );

    \I__8052\ : InMux
    port map (
            O => \N__32734\,
            I => \N__32702\
        );

    \I__8051\ : InMux
    port map (
            O => \N__32733\,
            I => \N__32702\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__32724\,
            I => \N__32697\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__32715\,
            I => \N__32697\
        );

    \I__8048\ : Span4Mux_h
    port map (
            O => \N__32712\,
            I => \N__32694\
        );

    \I__8047\ : Span4Mux_h
    port map (
            O => \N__32709\,
            I => \N__32691\
        );

    \I__8046\ : LocalMux
    port map (
            O => \N__32702\,
            I => \N_39\
        );

    \I__8045\ : Odrv12
    port map (
            O => \N__32697\,
            I => \N_39\
        );

    \I__8044\ : Odrv4
    port map (
            O => \N__32694\,
            I => \N_39\
        );

    \I__8043\ : Odrv4
    port map (
            O => \N__32691\,
            I => \N_39\
        );

    \I__8042\ : IoInMux
    port map (
            O => \N__32682\,
            I => \N__32679\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__32679\,
            I => \N__32676\
        );

    \I__8040\ : Span12Mux_s7_v
    port map (
            O => \N__32676\,
            I => \N__32672\
        );

    \I__8039\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32669\
        );

    \I__8038\ : Odrv12
    port map (
            O => \N__32672\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__32669\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__8036\ : ClkMux
    port map (
            O => \N__32664\,
            I => \N__32241\
        );

    \I__8035\ : ClkMux
    port map (
            O => \N__32663\,
            I => \N__32241\
        );

    \I__8034\ : ClkMux
    port map (
            O => \N__32662\,
            I => \N__32241\
        );

    \I__8033\ : ClkMux
    port map (
            O => \N__32661\,
            I => \N__32241\
        );

    \I__8032\ : ClkMux
    port map (
            O => \N__32660\,
            I => \N__32241\
        );

    \I__8031\ : ClkMux
    port map (
            O => \N__32659\,
            I => \N__32241\
        );

    \I__8030\ : ClkMux
    port map (
            O => \N__32658\,
            I => \N__32241\
        );

    \I__8029\ : ClkMux
    port map (
            O => \N__32657\,
            I => \N__32241\
        );

    \I__8028\ : ClkMux
    port map (
            O => \N__32656\,
            I => \N__32241\
        );

    \I__8027\ : ClkMux
    port map (
            O => \N__32655\,
            I => \N__32241\
        );

    \I__8026\ : ClkMux
    port map (
            O => \N__32654\,
            I => \N__32241\
        );

    \I__8025\ : ClkMux
    port map (
            O => \N__32653\,
            I => \N__32241\
        );

    \I__8024\ : ClkMux
    port map (
            O => \N__32652\,
            I => \N__32241\
        );

    \I__8023\ : ClkMux
    port map (
            O => \N__32651\,
            I => \N__32241\
        );

    \I__8022\ : ClkMux
    port map (
            O => \N__32650\,
            I => \N__32241\
        );

    \I__8021\ : ClkMux
    port map (
            O => \N__32649\,
            I => \N__32241\
        );

    \I__8020\ : ClkMux
    port map (
            O => \N__32648\,
            I => \N__32241\
        );

    \I__8019\ : ClkMux
    port map (
            O => \N__32647\,
            I => \N__32241\
        );

    \I__8018\ : ClkMux
    port map (
            O => \N__32646\,
            I => \N__32241\
        );

    \I__8017\ : ClkMux
    port map (
            O => \N__32645\,
            I => \N__32241\
        );

    \I__8016\ : ClkMux
    port map (
            O => \N__32644\,
            I => \N__32241\
        );

    \I__8015\ : ClkMux
    port map (
            O => \N__32643\,
            I => \N__32241\
        );

    \I__8014\ : ClkMux
    port map (
            O => \N__32642\,
            I => \N__32241\
        );

    \I__8013\ : ClkMux
    port map (
            O => \N__32641\,
            I => \N__32241\
        );

    \I__8012\ : ClkMux
    port map (
            O => \N__32640\,
            I => \N__32241\
        );

    \I__8011\ : ClkMux
    port map (
            O => \N__32639\,
            I => \N__32241\
        );

    \I__8010\ : ClkMux
    port map (
            O => \N__32638\,
            I => \N__32241\
        );

    \I__8009\ : ClkMux
    port map (
            O => \N__32637\,
            I => \N__32241\
        );

    \I__8008\ : ClkMux
    port map (
            O => \N__32636\,
            I => \N__32241\
        );

    \I__8007\ : ClkMux
    port map (
            O => \N__32635\,
            I => \N__32241\
        );

    \I__8006\ : ClkMux
    port map (
            O => \N__32634\,
            I => \N__32241\
        );

    \I__8005\ : ClkMux
    port map (
            O => \N__32633\,
            I => \N__32241\
        );

    \I__8004\ : ClkMux
    port map (
            O => \N__32632\,
            I => \N__32241\
        );

    \I__8003\ : ClkMux
    port map (
            O => \N__32631\,
            I => \N__32241\
        );

    \I__8002\ : ClkMux
    port map (
            O => \N__32630\,
            I => \N__32241\
        );

    \I__8001\ : ClkMux
    port map (
            O => \N__32629\,
            I => \N__32241\
        );

    \I__8000\ : ClkMux
    port map (
            O => \N__32628\,
            I => \N__32241\
        );

    \I__7999\ : ClkMux
    port map (
            O => \N__32627\,
            I => \N__32241\
        );

    \I__7998\ : ClkMux
    port map (
            O => \N__32626\,
            I => \N__32241\
        );

    \I__7997\ : ClkMux
    port map (
            O => \N__32625\,
            I => \N__32241\
        );

    \I__7996\ : ClkMux
    port map (
            O => \N__32624\,
            I => \N__32241\
        );

    \I__7995\ : ClkMux
    port map (
            O => \N__32623\,
            I => \N__32241\
        );

    \I__7994\ : ClkMux
    port map (
            O => \N__32622\,
            I => \N__32241\
        );

    \I__7993\ : ClkMux
    port map (
            O => \N__32621\,
            I => \N__32241\
        );

    \I__7992\ : ClkMux
    port map (
            O => \N__32620\,
            I => \N__32241\
        );

    \I__7991\ : ClkMux
    port map (
            O => \N__32619\,
            I => \N__32241\
        );

    \I__7990\ : ClkMux
    port map (
            O => \N__32618\,
            I => \N__32241\
        );

    \I__7989\ : ClkMux
    port map (
            O => \N__32617\,
            I => \N__32241\
        );

    \I__7988\ : ClkMux
    port map (
            O => \N__32616\,
            I => \N__32241\
        );

    \I__7987\ : ClkMux
    port map (
            O => \N__32615\,
            I => \N__32241\
        );

    \I__7986\ : ClkMux
    port map (
            O => \N__32614\,
            I => \N__32241\
        );

    \I__7985\ : ClkMux
    port map (
            O => \N__32613\,
            I => \N__32241\
        );

    \I__7984\ : ClkMux
    port map (
            O => \N__32612\,
            I => \N__32241\
        );

    \I__7983\ : ClkMux
    port map (
            O => \N__32611\,
            I => \N__32241\
        );

    \I__7982\ : ClkMux
    port map (
            O => \N__32610\,
            I => \N__32241\
        );

    \I__7981\ : ClkMux
    port map (
            O => \N__32609\,
            I => \N__32241\
        );

    \I__7980\ : ClkMux
    port map (
            O => \N__32608\,
            I => \N__32241\
        );

    \I__7979\ : ClkMux
    port map (
            O => \N__32607\,
            I => \N__32241\
        );

    \I__7978\ : ClkMux
    port map (
            O => \N__32606\,
            I => \N__32241\
        );

    \I__7977\ : ClkMux
    port map (
            O => \N__32605\,
            I => \N__32241\
        );

    \I__7976\ : ClkMux
    port map (
            O => \N__32604\,
            I => \N__32241\
        );

    \I__7975\ : ClkMux
    port map (
            O => \N__32603\,
            I => \N__32241\
        );

    \I__7974\ : ClkMux
    port map (
            O => \N__32602\,
            I => \N__32241\
        );

    \I__7973\ : ClkMux
    port map (
            O => \N__32601\,
            I => \N__32241\
        );

    \I__7972\ : ClkMux
    port map (
            O => \N__32600\,
            I => \N__32241\
        );

    \I__7971\ : ClkMux
    port map (
            O => \N__32599\,
            I => \N__32241\
        );

    \I__7970\ : ClkMux
    port map (
            O => \N__32598\,
            I => \N__32241\
        );

    \I__7969\ : ClkMux
    port map (
            O => \N__32597\,
            I => \N__32241\
        );

    \I__7968\ : ClkMux
    port map (
            O => \N__32596\,
            I => \N__32241\
        );

    \I__7967\ : ClkMux
    port map (
            O => \N__32595\,
            I => \N__32241\
        );

    \I__7966\ : ClkMux
    port map (
            O => \N__32594\,
            I => \N__32241\
        );

    \I__7965\ : ClkMux
    port map (
            O => \N__32593\,
            I => \N__32241\
        );

    \I__7964\ : ClkMux
    port map (
            O => \N__32592\,
            I => \N__32241\
        );

    \I__7963\ : ClkMux
    port map (
            O => \N__32591\,
            I => \N__32241\
        );

    \I__7962\ : ClkMux
    port map (
            O => \N__32590\,
            I => \N__32241\
        );

    \I__7961\ : ClkMux
    port map (
            O => \N__32589\,
            I => \N__32241\
        );

    \I__7960\ : ClkMux
    port map (
            O => \N__32588\,
            I => \N__32241\
        );

    \I__7959\ : ClkMux
    port map (
            O => \N__32587\,
            I => \N__32241\
        );

    \I__7958\ : ClkMux
    port map (
            O => \N__32586\,
            I => \N__32241\
        );

    \I__7957\ : ClkMux
    port map (
            O => \N__32585\,
            I => \N__32241\
        );

    \I__7956\ : ClkMux
    port map (
            O => \N__32584\,
            I => \N__32241\
        );

    \I__7955\ : ClkMux
    port map (
            O => \N__32583\,
            I => \N__32241\
        );

    \I__7954\ : ClkMux
    port map (
            O => \N__32582\,
            I => \N__32241\
        );

    \I__7953\ : ClkMux
    port map (
            O => \N__32581\,
            I => \N__32241\
        );

    \I__7952\ : ClkMux
    port map (
            O => \N__32580\,
            I => \N__32241\
        );

    \I__7951\ : ClkMux
    port map (
            O => \N__32579\,
            I => \N__32241\
        );

    \I__7950\ : ClkMux
    port map (
            O => \N__32578\,
            I => \N__32241\
        );

    \I__7949\ : ClkMux
    port map (
            O => \N__32577\,
            I => \N__32241\
        );

    \I__7948\ : ClkMux
    port map (
            O => \N__32576\,
            I => \N__32241\
        );

    \I__7947\ : ClkMux
    port map (
            O => \N__32575\,
            I => \N__32241\
        );

    \I__7946\ : ClkMux
    port map (
            O => \N__32574\,
            I => \N__32241\
        );

    \I__7945\ : ClkMux
    port map (
            O => \N__32573\,
            I => \N__32241\
        );

    \I__7944\ : ClkMux
    port map (
            O => \N__32572\,
            I => \N__32241\
        );

    \I__7943\ : ClkMux
    port map (
            O => \N__32571\,
            I => \N__32241\
        );

    \I__7942\ : ClkMux
    port map (
            O => \N__32570\,
            I => \N__32241\
        );

    \I__7941\ : ClkMux
    port map (
            O => \N__32569\,
            I => \N__32241\
        );

    \I__7940\ : ClkMux
    port map (
            O => \N__32568\,
            I => \N__32241\
        );

    \I__7939\ : ClkMux
    port map (
            O => \N__32567\,
            I => \N__32241\
        );

    \I__7938\ : ClkMux
    port map (
            O => \N__32566\,
            I => \N__32241\
        );

    \I__7937\ : ClkMux
    port map (
            O => \N__32565\,
            I => \N__32241\
        );

    \I__7936\ : ClkMux
    port map (
            O => \N__32564\,
            I => \N__32241\
        );

    \I__7935\ : ClkMux
    port map (
            O => \N__32563\,
            I => \N__32241\
        );

    \I__7934\ : ClkMux
    port map (
            O => \N__32562\,
            I => \N__32241\
        );

    \I__7933\ : ClkMux
    port map (
            O => \N__32561\,
            I => \N__32241\
        );

    \I__7932\ : ClkMux
    port map (
            O => \N__32560\,
            I => \N__32241\
        );

    \I__7931\ : ClkMux
    port map (
            O => \N__32559\,
            I => \N__32241\
        );

    \I__7930\ : ClkMux
    port map (
            O => \N__32558\,
            I => \N__32241\
        );

    \I__7929\ : ClkMux
    port map (
            O => \N__32557\,
            I => \N__32241\
        );

    \I__7928\ : ClkMux
    port map (
            O => \N__32556\,
            I => \N__32241\
        );

    \I__7927\ : ClkMux
    port map (
            O => \N__32555\,
            I => \N__32241\
        );

    \I__7926\ : ClkMux
    port map (
            O => \N__32554\,
            I => \N__32241\
        );

    \I__7925\ : ClkMux
    port map (
            O => \N__32553\,
            I => \N__32241\
        );

    \I__7924\ : ClkMux
    port map (
            O => \N__32552\,
            I => \N__32241\
        );

    \I__7923\ : ClkMux
    port map (
            O => \N__32551\,
            I => \N__32241\
        );

    \I__7922\ : ClkMux
    port map (
            O => \N__32550\,
            I => \N__32241\
        );

    \I__7921\ : ClkMux
    port map (
            O => \N__32549\,
            I => \N__32241\
        );

    \I__7920\ : ClkMux
    port map (
            O => \N__32548\,
            I => \N__32241\
        );

    \I__7919\ : ClkMux
    port map (
            O => \N__32547\,
            I => \N__32241\
        );

    \I__7918\ : ClkMux
    port map (
            O => \N__32546\,
            I => \N__32241\
        );

    \I__7917\ : ClkMux
    port map (
            O => \N__32545\,
            I => \N__32241\
        );

    \I__7916\ : ClkMux
    port map (
            O => \N__32544\,
            I => \N__32241\
        );

    \I__7915\ : ClkMux
    port map (
            O => \N__32543\,
            I => \N__32241\
        );

    \I__7914\ : ClkMux
    port map (
            O => \N__32542\,
            I => \N__32241\
        );

    \I__7913\ : ClkMux
    port map (
            O => \N__32541\,
            I => \N__32241\
        );

    \I__7912\ : ClkMux
    port map (
            O => \N__32540\,
            I => \N__32241\
        );

    \I__7911\ : ClkMux
    port map (
            O => \N__32539\,
            I => \N__32241\
        );

    \I__7910\ : ClkMux
    port map (
            O => \N__32538\,
            I => \N__32241\
        );

    \I__7909\ : ClkMux
    port map (
            O => \N__32537\,
            I => \N__32241\
        );

    \I__7908\ : ClkMux
    port map (
            O => \N__32536\,
            I => \N__32241\
        );

    \I__7907\ : ClkMux
    port map (
            O => \N__32535\,
            I => \N__32241\
        );

    \I__7906\ : ClkMux
    port map (
            O => \N__32534\,
            I => \N__32241\
        );

    \I__7905\ : ClkMux
    port map (
            O => \N__32533\,
            I => \N__32241\
        );

    \I__7904\ : ClkMux
    port map (
            O => \N__32532\,
            I => \N__32241\
        );

    \I__7903\ : ClkMux
    port map (
            O => \N__32531\,
            I => \N__32241\
        );

    \I__7902\ : ClkMux
    port map (
            O => \N__32530\,
            I => \N__32241\
        );

    \I__7901\ : ClkMux
    port map (
            O => \N__32529\,
            I => \N__32241\
        );

    \I__7900\ : ClkMux
    port map (
            O => \N__32528\,
            I => \N__32241\
        );

    \I__7899\ : ClkMux
    port map (
            O => \N__32527\,
            I => \N__32241\
        );

    \I__7898\ : ClkMux
    port map (
            O => \N__32526\,
            I => \N__32241\
        );

    \I__7897\ : ClkMux
    port map (
            O => \N__32525\,
            I => \N__32241\
        );

    \I__7896\ : ClkMux
    port map (
            O => \N__32524\,
            I => \N__32241\
        );

    \I__7895\ : GlobalMux
    port map (
            O => \N__32241\,
            I => \N__32238\
        );

    \I__7894\ : gio2CtrlBuf
    port map (
            O => \N__32238\,
            I => clk_0_c_g
        );

    \I__7893\ : CEMux
    port map (
            O => \N__32235\,
            I => \N__32230\
        );

    \I__7892\ : CEMux
    port map (
            O => \N__32234\,
            I => \N__32227\
        );

    \I__7891\ : CEMux
    port map (
            O => \N__32233\,
            I => \N__32224\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__32230\,
            I => \N__32221\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__32227\,
            I => \N__32217\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__32224\,
            I => \N__32214\
        );

    \I__7887\ : Span4Mux_h
    port map (
            O => \N__32221\,
            I => \N__32211\
        );

    \I__7886\ : CEMux
    port map (
            O => \N__32220\,
            I => \N__32208\
        );

    \I__7885\ : Span4Mux_h
    port map (
            O => \N__32217\,
            I => \N__32205\
        );

    \I__7884\ : Span4Mux_h
    port map (
            O => \N__32214\,
            I => \N__32202\
        );

    \I__7883\ : Span4Mux_h
    port map (
            O => \N__32211\,
            I => \N__32199\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__32208\,
            I => \N__32196\
        );

    \I__7881\ : Odrv4
    port map (
            O => \N__32205\,
            I => \N_37\
        );

    \I__7880\ : Odrv4
    port map (
            O => \N__32202\,
            I => \N_37\
        );

    \I__7879\ : Odrv4
    port map (
            O => \N__32199\,
            I => \N_37\
        );

    \I__7878\ : Odrv4
    port map (
            O => \N__32196\,
            I => \N_37\
        );

    \I__7877\ : InMux
    port map (
            O => \N__32187\,
            I => \N__32184\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__32184\,
            I => \N__32181\
        );

    \I__7875\ : Span4Mux_h
    port map (
            O => \N__32181\,
            I => \N__32178\
        );

    \I__7874\ : Sp12to4
    port map (
            O => \N__32178\,
            I => \N__32171\
        );

    \I__7873\ : InMux
    port map (
            O => \N__32177\,
            I => \N__32168\
        );

    \I__7872\ : CascadeMux
    port map (
            O => \N__32176\,
            I => \N__32165\
        );

    \I__7871\ : InMux
    port map (
            O => \N__32175\,
            I => \N__32160\
        );

    \I__7870\ : InMux
    port map (
            O => \N__32174\,
            I => \N__32160\
        );

    \I__7869\ : Span12Mux_v
    port map (
            O => \N__32171\,
            I => \N__32157\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__32168\,
            I => \N__32154\
        );

    \I__7867\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32151\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__32160\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__7865\ : Odrv12
    port map (
            O => \N__32157\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__7864\ : Odrv4
    port map (
            O => \N__32154\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__32151\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__7862\ : InMux
    port map (
            O => \N__32142\,
            I => \N__32137\
        );

    \I__7861\ : InMux
    port map (
            O => \N__32141\,
            I => \N__32125\
        );

    \I__7860\ : InMux
    port map (
            O => \N__32140\,
            I => \N__32120\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__32137\,
            I => \N__32116\
        );

    \I__7858\ : InMux
    port map (
            O => \N__32136\,
            I => \N__32113\
        );

    \I__7857\ : InMux
    port map (
            O => \N__32135\,
            I => \N__32106\
        );

    \I__7856\ : InMux
    port map (
            O => \N__32134\,
            I => \N__32106\
        );

    \I__7855\ : InMux
    port map (
            O => \N__32133\,
            I => \N__32106\
        );

    \I__7854\ : InMux
    port map (
            O => \N__32132\,
            I => \N__32103\
        );

    \I__7853\ : InMux
    port map (
            O => \N__32131\,
            I => \N__32099\
        );

    \I__7852\ : InMux
    port map (
            O => \N__32130\,
            I => \N__32096\
        );

    \I__7851\ : InMux
    port map (
            O => \N__32129\,
            I => \N__32091\
        );

    \I__7850\ : InMux
    port map (
            O => \N__32128\,
            I => \N__32091\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__32125\,
            I => \N__32088\
        );

    \I__7848\ : InMux
    port map (
            O => \N__32124\,
            I => \N__32085\
        );

    \I__7847\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32082\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__32120\,
            I => \N__32079\
        );

    \I__7845\ : InMux
    port map (
            O => \N__32119\,
            I => \N__32072\
        );

    \I__7844\ : Span4Mux_h
    port map (
            O => \N__32116\,
            I => \N__32063\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__32113\,
            I => \N__32063\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__32106\,
            I => \N__32063\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__32103\,
            I => \N__32063\
        );

    \I__7840\ : InMux
    port map (
            O => \N__32102\,
            I => \N__32060\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__32099\,
            I => \N__32053\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__32096\,
            I => \N__32053\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__32091\,
            I => \N__32053\
        );

    \I__7836\ : Span4Mux_h
    port map (
            O => \N__32088\,
            I => \N__32048\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__32085\,
            I => \N__32048\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__32082\,
            I => \N__32045\
        );

    \I__7833\ : Span4Mux_h
    port map (
            O => \N__32079\,
            I => \N__32042\
        );

    \I__7832\ : InMux
    port map (
            O => \N__32078\,
            I => \N__32035\
        );

    \I__7831\ : InMux
    port map (
            O => \N__32077\,
            I => \N__32035\
        );

    \I__7830\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32035\
        );

    \I__7829\ : InMux
    port map (
            O => \N__32075\,
            I => \N__32032\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__32072\,
            I => \N__32029\
        );

    \I__7827\ : Span4Mux_v
    port map (
            O => \N__32063\,
            I => \N__32026\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__32060\,
            I => \N__32021\
        );

    \I__7825\ : Span4Mux_h
    port map (
            O => \N__32053\,
            I => \N__32021\
        );

    \I__7824\ : Span4Mux_h
    port map (
            O => \N__32048\,
            I => \N__32016\
        );

    \I__7823\ : Span4Mux_h
    port map (
            O => \N__32045\,
            I => \N__32016\
        );

    \I__7822\ : Sp12to4
    port map (
            O => \N__32042\,
            I => \N__32011\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__32035\,
            I => \N__32011\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__32032\,
            I => \N__32008\
        );

    \I__7819\ : Span4Mux_s2_v
    port map (
            O => \N__32029\,
            I => \N__32005\
        );

    \I__7818\ : Span4Mux_v
    port map (
            O => \N__32026\,
            I => \N__32002\
        );

    \I__7817\ : Span4Mux_h
    port map (
            O => \N__32021\,
            I => \N__31999\
        );

    \I__7816\ : Span4Mux_v
    port map (
            O => \N__32016\,
            I => \N__31996\
        );

    \I__7815\ : Span12Mux_v
    port map (
            O => \N__32011\,
            I => \N__31993\
        );

    \I__7814\ : Span4Mux_s2_v
    port map (
            O => \N__32008\,
            I => \N__31990\
        );

    \I__7813\ : Span4Mux_h
    port map (
            O => \N__32005\,
            I => \N__31985\
        );

    \I__7812\ : Span4Mux_v
    port map (
            O => \N__32002\,
            I => \N__31985\
        );

    \I__7811\ : Span4Mux_h
    port map (
            O => \N__31999\,
            I => \N__31980\
        );

    \I__7810\ : Span4Mux_v
    port map (
            O => \N__31996\,
            I => \N__31980\
        );

    \I__7809\ : Odrv12
    port map (
            O => \N__31993\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__7808\ : Odrv4
    port map (
            O => \N__31990\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__7807\ : Odrv4
    port map (
            O => \N__31985\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__7806\ : Odrv4
    port map (
            O => \N__31980\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__7805\ : CascadeMux
    port map (
            O => \N__31971\,
            I => \N__31966\
        );

    \I__7804\ : CascadeMux
    port map (
            O => \N__31970\,
            I => \N__31961\
        );

    \I__7803\ : CascadeMux
    port map (
            O => \N__31969\,
            I => \N__31957\
        );

    \I__7802\ : InMux
    port map (
            O => \N__31966\,
            I => \N__31954\
        );

    \I__7801\ : InMux
    port map (
            O => \N__31965\,
            I => \N__31951\
        );

    \I__7800\ : CascadeMux
    port map (
            O => \N__31964\,
            I => \N__31948\
        );

    \I__7799\ : InMux
    port map (
            O => \N__31961\,
            I => \N__31945\
        );

    \I__7798\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31940\
        );

    \I__7797\ : InMux
    port map (
            O => \N__31957\,
            I => \N__31940\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__31954\,
            I => \N__31936\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__31951\,
            I => \N__31931\
        );

    \I__7794\ : InMux
    port map (
            O => \N__31948\,
            I => \N__31928\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__31945\,
            I => \N__31923\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__31940\,
            I => \N__31923\
        );

    \I__7791\ : CascadeMux
    port map (
            O => \N__31939\,
            I => \N__31920\
        );

    \I__7790\ : Span4Mux_v
    port map (
            O => \N__31936\,
            I => \N__31916\
        );

    \I__7789\ : CascadeMux
    port map (
            O => \N__31935\,
            I => \N__31913\
        );

    \I__7788\ : CascadeMux
    port map (
            O => \N__31934\,
            I => \N__31909\
        );

    \I__7787\ : Span4Mux_v
    port map (
            O => \N__31931\,
            I => \N__31906\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__31928\,
            I => \N__31901\
        );

    \I__7785\ : Span4Mux_h
    port map (
            O => \N__31923\,
            I => \N__31901\
        );

    \I__7784\ : InMux
    port map (
            O => \N__31920\,
            I => \N__31898\
        );

    \I__7783\ : InMux
    port map (
            O => \N__31919\,
            I => \N__31895\
        );

    \I__7782\ : Span4Mux_v
    port map (
            O => \N__31916\,
            I => \N__31892\
        );

    \I__7781\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31889\
        );

    \I__7780\ : CascadeMux
    port map (
            O => \N__31912\,
            I => \N__31886\
        );

    \I__7779\ : InMux
    port map (
            O => \N__31909\,
            I => \N__31879\
        );

    \I__7778\ : Span4Mux_h
    port map (
            O => \N__31906\,
            I => \N__31872\
        );

    \I__7777\ : Span4Mux_h
    port map (
            O => \N__31901\,
            I => \N__31872\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__31898\,
            I => \N__31872\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__31895\,
            I => \N__31869\
        );

    \I__7774\ : Span4Mux_v
    port map (
            O => \N__31892\,
            I => \N__31864\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__31889\,
            I => \N__31864\
        );

    \I__7772\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31857\
        );

    \I__7771\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31857\
        );

    \I__7770\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31857\
        );

    \I__7769\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31853\
        );

    \I__7768\ : CascadeMux
    port map (
            O => \N__31882\,
            I => \N__31850\
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__31879\,
            I => \N__31845\
        );

    \I__7766\ : Sp12to4
    port map (
            O => \N__31872\,
            I => \N__31845\
        );

    \I__7765\ : Span4Mux_h
    port map (
            O => \N__31869\,
            I => \N__31842\
        );

    \I__7764\ : Span4Mux_h
    port map (
            O => \N__31864\,
            I => \N__31837\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__31857\,
            I => \N__31837\
        );

    \I__7762\ : InMux
    port map (
            O => \N__31856\,
            I => \N__31834\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__31853\,
            I => \N__31831\
        );

    \I__7760\ : InMux
    port map (
            O => \N__31850\,
            I => \N__31828\
        );

    \I__7759\ : Span12Mux_v
    port map (
            O => \N__31845\,
            I => \N__31825\
        );

    \I__7758\ : Span4Mux_h
    port map (
            O => \N__31842\,
            I => \N__31820\
        );

    \I__7757\ : Span4Mux_h
    port map (
            O => \N__31837\,
            I => \N__31820\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__31834\,
            I => \N__31815\
        );

    \I__7755\ : Span4Mux_h
    port map (
            O => \N__31831\,
            I => \N__31815\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__31828\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__7753\ : Odrv12
    port map (
            O => \N__31825\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__7752\ : Odrv4
    port map (
            O => \N__31820\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__7751\ : Odrv4
    port map (
            O => \N__31815\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__7750\ : InMux
    port map (
            O => \N__31806\,
            I => \N__31803\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__31803\,
            I => \N__31800\
        );

    \I__7748\ : Span12Mux_s11_h
    port map (
            O => \N__31800\,
            I => \N__31797\
        );

    \I__7747\ : Span12Mux_v
    port map (
            O => \N__31797\,
            I => \N__31794\
        );

    \I__7746\ : Odrv12
    port map (
            O => \N__31794\,
            I => \this_ppu.un3_sprites_addr_cry_3_c_RNI1VDZ0Z8\
        );

    \I__7745\ : CascadeMux
    port map (
            O => \N__31791\,
            I => \N__31788\
        );

    \I__7744\ : CascadeBuf
    port map (
            O => \N__31788\,
            I => \N__31785\
        );

    \I__7743\ : CascadeMux
    port map (
            O => \N__31785\,
            I => \N__31782\
        );

    \I__7742\ : CascadeBuf
    port map (
            O => \N__31782\,
            I => \N__31779\
        );

    \I__7741\ : CascadeMux
    port map (
            O => \N__31779\,
            I => \N__31776\
        );

    \I__7740\ : CascadeBuf
    port map (
            O => \N__31776\,
            I => \N__31773\
        );

    \I__7739\ : CascadeMux
    port map (
            O => \N__31773\,
            I => \N__31770\
        );

    \I__7738\ : CascadeBuf
    port map (
            O => \N__31770\,
            I => \N__31767\
        );

    \I__7737\ : CascadeMux
    port map (
            O => \N__31767\,
            I => \N__31764\
        );

    \I__7736\ : CascadeBuf
    port map (
            O => \N__31764\,
            I => \N__31761\
        );

    \I__7735\ : CascadeMux
    port map (
            O => \N__31761\,
            I => \N__31758\
        );

    \I__7734\ : CascadeBuf
    port map (
            O => \N__31758\,
            I => \N__31755\
        );

    \I__7733\ : CascadeMux
    port map (
            O => \N__31755\,
            I => \N__31752\
        );

    \I__7732\ : CascadeBuf
    port map (
            O => \N__31752\,
            I => \N__31749\
        );

    \I__7731\ : CascadeMux
    port map (
            O => \N__31749\,
            I => \N__31746\
        );

    \I__7730\ : CascadeBuf
    port map (
            O => \N__31746\,
            I => \N__31743\
        );

    \I__7729\ : CascadeMux
    port map (
            O => \N__31743\,
            I => \N__31740\
        );

    \I__7728\ : CascadeBuf
    port map (
            O => \N__31740\,
            I => \N__31737\
        );

    \I__7727\ : CascadeMux
    port map (
            O => \N__31737\,
            I => \N__31734\
        );

    \I__7726\ : CascadeBuf
    port map (
            O => \N__31734\,
            I => \N__31731\
        );

    \I__7725\ : CascadeMux
    port map (
            O => \N__31731\,
            I => \N__31728\
        );

    \I__7724\ : CascadeBuf
    port map (
            O => \N__31728\,
            I => \N__31725\
        );

    \I__7723\ : CascadeMux
    port map (
            O => \N__31725\,
            I => \N__31722\
        );

    \I__7722\ : CascadeBuf
    port map (
            O => \N__31722\,
            I => \N__31719\
        );

    \I__7721\ : CascadeMux
    port map (
            O => \N__31719\,
            I => \N__31716\
        );

    \I__7720\ : CascadeBuf
    port map (
            O => \N__31716\,
            I => \N__31713\
        );

    \I__7719\ : CascadeMux
    port map (
            O => \N__31713\,
            I => \N__31710\
        );

    \I__7718\ : CascadeBuf
    port map (
            O => \N__31710\,
            I => \N__31707\
        );

    \I__7717\ : CascadeMux
    port map (
            O => \N__31707\,
            I => \N__31704\
        );

    \I__7716\ : CascadeBuf
    port map (
            O => \N__31704\,
            I => \N__31701\
        );

    \I__7715\ : CascadeMux
    port map (
            O => \N__31701\,
            I => \N__31698\
        );

    \I__7714\ : InMux
    port map (
            O => \N__31698\,
            I => \N__31695\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__31695\,
            I => \N__31692\
        );

    \I__7712\ : Odrv4
    port map (
            O => \N__31692\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__7711\ : InMux
    port map (
            O => \N__31689\,
            I => \N__31686\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__31686\,
            I => \N__31683\
        );

    \I__7709\ : Span4Mux_v
    port map (
            O => \N__31683\,
            I => \N__31680\
        );

    \I__7708\ : Span4Mux_v
    port map (
            O => \N__31680\,
            I => \N__31677\
        );

    \I__7707\ : Span4Mux_v
    port map (
            O => \N__31677\,
            I => \N__31674\
        );

    \I__7706\ : Span4Mux_v
    port map (
            O => \N__31674\,
            I => \N__31671\
        );

    \I__7705\ : Odrv4
    port map (
            O => \N__31671\,
            I => port_address_in_7
        );

    \I__7704\ : InMux
    port map (
            O => \N__31668\,
            I => \N__31665\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__31665\,
            I => \N__31662\
        );

    \I__7702\ : IoSpan4Mux
    port map (
            O => \N__31662\,
            I => \N__31659\
        );

    \I__7701\ : Odrv4
    port map (
            O => \N__31659\,
            I => port_address_in_4
        );

    \I__7700\ : CascadeMux
    port map (
            O => \N__31656\,
            I => \N__31653\
        );

    \I__7699\ : InMux
    port map (
            O => \N__31653\,
            I => \N__31650\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__31650\,
            I => \N__31646\
        );

    \I__7697\ : InMux
    port map (
            O => \N__31649\,
            I => \N__31643\
        );

    \I__7696\ : Span4Mux_s2_h
    port map (
            O => \N__31646\,
            I => \N__31640\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__31643\,
            I => \N__31637\
        );

    \I__7694\ : Sp12to4
    port map (
            O => \N__31640\,
            I => \N__31634\
        );

    \I__7693\ : Span4Mux_h
    port map (
            O => \N__31637\,
            I => \N__31631\
        );

    \I__7692\ : Span12Mux_s11_v
    port map (
            O => \N__31634\,
            I => \N__31628\
        );

    \I__7691\ : Span4Mux_v
    port map (
            O => \N__31631\,
            I => \N__31625\
        );

    \I__7690\ : Span12Mux_h
    port map (
            O => \N__31628\,
            I => \N__31622\
        );

    \I__7689\ : Sp12to4
    port map (
            O => \N__31625\,
            I => \N__31619\
        );

    \I__7688\ : Span12Mux_h
    port map (
            O => \N__31622\,
            I => \N__31616\
        );

    \I__7687\ : Span12Mux_h
    port map (
            O => \N__31619\,
            I => \N__31613\
        );

    \I__7686\ : Odrv12
    port map (
            O => \N__31616\,
            I => port_rw_in
        );

    \I__7685\ : Odrv12
    port map (
            O => \N__31613\,
            I => port_rw_in
        );

    \I__7684\ : InMux
    port map (
            O => \N__31608\,
            I => \N__31605\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__31605\,
            I => \N__31602\
        );

    \I__7682\ : Span12Mux_v
    port map (
            O => \N__31602\,
            I => \N__31599\
        );

    \I__7681\ : Odrv12
    port map (
            O => \N__31599\,
            I => port_address_in_3
        );

    \I__7680\ : InMux
    port map (
            O => \N__31596\,
            I => \N__31593\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__31593\,
            I => \N__31590\
        );

    \I__7678\ : Span12Mux_h
    port map (
            O => \N__31590\,
            I => \N__31587\
        );

    \I__7677\ : Odrv12
    port map (
            O => \N__31587\,
            I => \this_start_data_delay.un1_M_this_state_q_17_i_o2_1Z0Z_4\
        );

    \I__7676\ : IoInMux
    port map (
            O => \N__31584\,
            I => \N__31581\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__31581\,
            I => \N__31578\
        );

    \I__7674\ : Span4Mux_s1_v
    port map (
            O => \N__31578\,
            I => \N__31574\
        );

    \I__7673\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31571\
        );

    \I__7672\ : Span4Mux_v
    port map (
            O => \N__31574\,
            I => \N__31568\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__31571\,
            I => \N__31565\
        );

    \I__7670\ : Odrv4
    port map (
            O => \N__31568\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__7669\ : Odrv4
    port map (
            O => \N__31565\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__7668\ : InMux
    port map (
            O => \N__31560\,
            I => \N__31557\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__31557\,
            I => \N__31554\
        );

    \I__7666\ : Odrv12
    port map (
            O => \N__31554\,
            I => \M_this_external_address_q_s_9\
        );

    \I__7665\ : InMux
    port map (
            O => \N__31551\,
            I => \M_this_external_address_q_cry_8\
        );

    \I__7664\ : InMux
    port map (
            O => \N__31548\,
            I => \M_this_external_address_q_cry_9\
        );

    \I__7663\ : InMux
    port map (
            O => \N__31545\,
            I => \M_this_external_address_q_cry_10\
        );

    \I__7662\ : IoInMux
    port map (
            O => \N__31542\,
            I => \N__31539\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__31539\,
            I => \N__31534\
        );

    \I__7660\ : CascadeMux
    port map (
            O => \N__31538\,
            I => \N__31531\
        );

    \I__7659\ : InMux
    port map (
            O => \N__31537\,
            I => \N__31528\
        );

    \I__7658\ : Sp12to4
    port map (
            O => \N__31534\,
            I => \N__31525\
        );

    \I__7657\ : InMux
    port map (
            O => \N__31531\,
            I => \N__31522\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__31528\,
            I => \N__31519\
        );

    \I__7655\ : Odrv12
    port map (
            O => \N__31525\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__31522\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__31519\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__7652\ : InMux
    port map (
            O => \N__31512\,
            I => \N__31509\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__31509\,
            I => \N__31506\
        );

    \I__7650\ : Odrv4
    port map (
            O => \N__31506\,
            I => \M_this_external_address_q_cry_11_THRU_CO\
        );

    \I__7649\ : InMux
    port map (
            O => \N__31503\,
            I => \M_this_external_address_q_cry_11\
        );

    \I__7648\ : IoInMux
    port map (
            O => \N__31500\,
            I => \N__31497\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__31497\,
            I => \N__31494\
        );

    \I__7646\ : IoSpan4Mux
    port map (
            O => \N__31494\,
            I => \N__31491\
        );

    \I__7645\ : Span4Mux_s2_h
    port map (
            O => \N__31491\,
            I => \N__31487\
        );

    \I__7644\ : InMux
    port map (
            O => \N__31490\,
            I => \N__31483\
        );

    \I__7643\ : Span4Mux_h
    port map (
            O => \N__31487\,
            I => \N__31480\
        );

    \I__7642\ : InMux
    port map (
            O => \N__31486\,
            I => \N__31477\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__31483\,
            I => \N__31474\
        );

    \I__7640\ : Odrv4
    port map (
            O => \N__31480\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__31477\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__7638\ : Odrv12
    port map (
            O => \N__31474\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__7637\ : CascadeMux
    port map (
            O => \N__31467\,
            I => \N__31464\
        );

    \I__7636\ : InMux
    port map (
            O => \N__31464\,
            I => \N__31461\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__31461\,
            I => \N__31458\
        );

    \I__7634\ : Odrv12
    port map (
            O => \N__31458\,
            I => \M_this_external_address_q_cry_12_THRU_CO\
        );

    \I__7633\ : InMux
    port map (
            O => \N__31455\,
            I => \M_this_external_address_q_cry_12\
        );

    \I__7632\ : IoInMux
    port map (
            O => \N__31452\,
            I => \N__31449\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__31449\,
            I => \N__31446\
        );

    \I__7630\ : Span4Mux_s3_h
    port map (
            O => \N__31446\,
            I => \N__31443\
        );

    \I__7629\ : Span4Mux_v
    port map (
            O => \N__31443\,
            I => \N__31438\
        );

    \I__7628\ : CascadeMux
    port map (
            O => \N__31442\,
            I => \N__31435\
        );

    \I__7627\ : InMux
    port map (
            O => \N__31441\,
            I => \N__31432\
        );

    \I__7626\ : Span4Mux_h
    port map (
            O => \N__31438\,
            I => \N__31429\
        );

    \I__7625\ : InMux
    port map (
            O => \N__31435\,
            I => \N__31426\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__31432\,
            I => \N__31423\
        );

    \I__7623\ : Odrv4
    port map (
            O => \N__31429\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__31426\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__7621\ : Odrv4
    port map (
            O => \N__31423\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__7620\ : InMux
    port map (
            O => \N__31416\,
            I => \N__31413\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__31413\,
            I => \N__31410\
        );

    \I__7618\ : Odrv4
    port map (
            O => \N__31410\,
            I => \M_this_external_address_q_cry_13_THRU_CO\
        );

    \I__7617\ : InMux
    port map (
            O => \N__31407\,
            I => \M_this_external_address_q_cry_13\
        );

    \I__7616\ : IoInMux
    port map (
            O => \N__31404\,
            I => \N__31401\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__31401\,
            I => \N__31398\
        );

    \I__7614\ : Span12Mux_s9_h
    port map (
            O => \N__31398\,
            I => \N__31394\
        );

    \I__7613\ : InMux
    port map (
            O => \N__31397\,
            I => \N__31391\
        );

    \I__7612\ : Span12Mux_v
    port map (
            O => \N__31394\,
            I => \N__31388\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__31391\,
            I => \N__31385\
        );

    \I__7610\ : Odrv12
    port map (
            O => \N__31388\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__7609\ : Odrv12
    port map (
            O => \N__31385\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__7608\ : InMux
    port map (
            O => \N__31380\,
            I => \M_this_external_address_q_cry_14\
        );

    \I__7607\ : CascadeMux
    port map (
            O => \N__31377\,
            I => \N__31374\
        );

    \I__7606\ : InMux
    port map (
            O => \N__31374\,
            I => \N__31371\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__31371\,
            I => \N__31368\
        );

    \I__7604\ : Odrv4
    port map (
            O => \N__31368\,
            I => \M_this_external_address_q_s_15\
        );

    \I__7603\ : InMux
    port map (
            O => \N__31365\,
            I => \N__31362\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__31362\,
            I => \M_this_external_address_q_s_11\
        );

    \I__7601\ : InMux
    port map (
            O => \N__31359\,
            I => \N__31352\
        );

    \I__7600\ : InMux
    port map (
            O => \N__31358\,
            I => \N__31349\
        );

    \I__7599\ : InMux
    port map (
            O => \N__31357\,
            I => \N__31346\
        );

    \I__7598\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31343\
        );

    \I__7597\ : CascadeMux
    port map (
            O => \N__31355\,
            I => \N__31339\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__31352\,
            I => \N__31334\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__31349\,
            I => \N__31334\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__31346\,
            I => \N__31331\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__31343\,
            I => \N__31327\
        );

    \I__7592\ : CascadeMux
    port map (
            O => \N__31342\,
            I => \N__31324\
        );

    \I__7591\ : InMux
    port map (
            O => \N__31339\,
            I => \N__31319\
        );

    \I__7590\ : Span4Mux_v
    port map (
            O => \N__31334\,
            I => \N__31314\
        );

    \I__7589\ : Span4Mux_h
    port map (
            O => \N__31331\,
            I => \N__31314\
        );

    \I__7588\ : InMux
    port map (
            O => \N__31330\,
            I => \N__31311\
        );

    \I__7587\ : Span4Mux_v
    port map (
            O => \N__31327\,
            I => \N__31308\
        );

    \I__7586\ : InMux
    port map (
            O => \N__31324\,
            I => \N__31305\
        );

    \I__7585\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31300\
        );

    \I__7584\ : InMux
    port map (
            O => \N__31322\,
            I => \N__31300\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__31319\,
            I => \N__31297\
        );

    \I__7582\ : Span4Mux_v
    port map (
            O => \N__31314\,
            I => \N__31290\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__31311\,
            I => \N__31290\
        );

    \I__7580\ : Span4Mux_h
    port map (
            O => \N__31308\,
            I => \N__31287\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__31305\,
            I => \N__31284\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__31300\,
            I => \N__31281\
        );

    \I__7577\ : Span4Mux_h
    port map (
            O => \N__31297\,
            I => \N__31278\
        );

    \I__7576\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31275\
        );

    \I__7575\ : CascadeMux
    port map (
            O => \N__31295\,
            I => \N__31272\
        );

    \I__7574\ : Span4Mux_v
    port map (
            O => \N__31290\,
            I => \N__31269\
        );

    \I__7573\ : Span4Mux_h
    port map (
            O => \N__31287\,
            I => \N__31264\
        );

    \I__7572\ : Span4Mux_v
    port map (
            O => \N__31284\,
            I => \N__31264\
        );

    \I__7571\ : Span4Mux_v
    port map (
            O => \N__31281\,
            I => \N__31257\
        );

    \I__7570\ : Span4Mux_h
    port map (
            O => \N__31278\,
            I => \N__31257\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__31275\,
            I => \N__31257\
        );

    \I__7568\ : InMux
    port map (
            O => \N__31272\,
            I => \N__31254\
        );

    \I__7567\ : Span4Mux_h
    port map (
            O => \N__31269\,
            I => \N__31251\
        );

    \I__7566\ : Sp12to4
    port map (
            O => \N__31264\,
            I => \N__31248\
        );

    \I__7565\ : Span4Mux_v
    port map (
            O => \N__31257\,
            I => \N__31245\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__31254\,
            I => \N__31242\
        );

    \I__7563\ : Sp12to4
    port map (
            O => \N__31251\,
            I => \N__31239\
        );

    \I__7562\ : Span12Mux_h
    port map (
            O => \N__31248\,
            I => \N__31236\
        );

    \I__7561\ : Sp12to4
    port map (
            O => \N__31245\,
            I => \N__31233\
        );

    \I__7560\ : Span4Mux_h
    port map (
            O => \N__31242\,
            I => \N__31230\
        );

    \I__7559\ : Span12Mux_h
    port map (
            O => \N__31239\,
            I => \N__31225\
        );

    \I__7558\ : Span12Mux_v
    port map (
            O => \N__31236\,
            I => \N__31225\
        );

    \I__7557\ : Span12Mux_h
    port map (
            O => \N__31233\,
            I => \N__31222\
        );

    \I__7556\ : Span4Mux_v
    port map (
            O => \N__31230\,
            I => \N__31219\
        );

    \I__7555\ : Odrv12
    port map (
            O => \N__31225\,
            I => port_data_c_3
        );

    \I__7554\ : Odrv12
    port map (
            O => \N__31222\,
            I => port_data_c_3
        );

    \I__7553\ : Odrv4
    port map (
            O => \N__31219\,
            I => port_data_c_3
        );

    \I__7552\ : IoInMux
    port map (
            O => \N__31212\,
            I => \N__31209\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__31209\,
            I => \N__31206\
        );

    \I__7550\ : Span4Mux_s3_v
    port map (
            O => \N__31206\,
            I => \N__31203\
        );

    \I__7549\ : Span4Mux_v
    port map (
            O => \N__31203\,
            I => \N__31199\
        );

    \I__7548\ : InMux
    port map (
            O => \N__31202\,
            I => \N__31196\
        );

    \I__7547\ : Odrv4
    port map (
            O => \N__31199\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__31196\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__7545\ : IoInMux
    port map (
            O => \N__31191\,
            I => \N__31188\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__31188\,
            I => \N__31185\
        );

    \I__7543\ : Span4Mux_s1_v
    port map (
            O => \N__31185\,
            I => \N__31182\
        );

    \I__7542\ : Sp12to4
    port map (
            O => \N__31182\,
            I => \N__31179\
        );

    \I__7541\ : Span12Mux_h
    port map (
            O => \N__31179\,
            I => \N__31175\
        );

    \I__7540\ : InMux
    port map (
            O => \N__31178\,
            I => \N__31172\
        );

    \I__7539\ : Odrv12
    port map (
            O => \N__31175\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__31172\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__7537\ : InMux
    port map (
            O => \N__31167\,
            I => \bfn_26_23_0_\
        );

    \I__7536\ : IoInMux
    port map (
            O => \N__31164\,
            I => \N__31161\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__31161\,
            I => \N__31158\
        );

    \I__7534\ : Sp12to4
    port map (
            O => \N__31158\,
            I => \N__31154\
        );

    \I__7533\ : InMux
    port map (
            O => \N__31157\,
            I => \N__31151\
        );

    \I__7532\ : Odrv12
    port map (
            O => \N__31154\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__31151\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__7530\ : InMux
    port map (
            O => \N__31146\,
            I => \M_this_external_address_q_cry_0\
        );

    \I__7529\ : IoInMux
    port map (
            O => \N__31143\,
            I => \N__31140\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__31140\,
            I => \N__31137\
        );

    \I__7527\ : IoSpan4Mux
    port map (
            O => \N__31137\,
            I => \N__31134\
        );

    \I__7526\ : Span4Mux_s2_v
    port map (
            O => \N__31134\,
            I => \N__31131\
        );

    \I__7525\ : Span4Mux_v
    port map (
            O => \N__31131\,
            I => \N__31127\
        );

    \I__7524\ : InMux
    port map (
            O => \N__31130\,
            I => \N__31124\
        );

    \I__7523\ : Odrv4
    port map (
            O => \N__31127\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__31124\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__7521\ : InMux
    port map (
            O => \N__31119\,
            I => \M_this_external_address_q_cry_1\
        );

    \I__7520\ : IoInMux
    port map (
            O => \N__31116\,
            I => \N__31113\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__31113\,
            I => \N__31110\
        );

    \I__7518\ : Span4Mux_s2_h
    port map (
            O => \N__31110\,
            I => \N__31107\
        );

    \I__7517\ : Span4Mux_h
    port map (
            O => \N__31107\,
            I => \N__31104\
        );

    \I__7516\ : Span4Mux_v
    port map (
            O => \N__31104\,
            I => \N__31100\
        );

    \I__7515\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31097\
        );

    \I__7514\ : Odrv4
    port map (
            O => \N__31100\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__31097\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__7512\ : InMux
    port map (
            O => \N__31092\,
            I => \M_this_external_address_q_cry_2\
        );

    \I__7511\ : IoInMux
    port map (
            O => \N__31089\,
            I => \N__31086\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__31086\,
            I => \N__31082\
        );

    \I__7509\ : InMux
    port map (
            O => \N__31085\,
            I => \N__31079\
        );

    \I__7508\ : Odrv12
    port map (
            O => \N__31082\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__31079\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__7506\ : InMux
    port map (
            O => \N__31074\,
            I => \M_this_external_address_q_cry_3\
        );

    \I__7505\ : IoInMux
    port map (
            O => \N__31071\,
            I => \N__31068\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__31068\,
            I => \N__31065\
        );

    \I__7503\ : IoSpan4Mux
    port map (
            O => \N__31065\,
            I => \N__31062\
        );

    \I__7502\ : Sp12to4
    port map (
            O => \N__31062\,
            I => \N__31058\
        );

    \I__7501\ : InMux
    port map (
            O => \N__31061\,
            I => \N__31055\
        );

    \I__7500\ : Odrv12
    port map (
            O => \N__31058\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__31055\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__7498\ : InMux
    port map (
            O => \N__31050\,
            I => \M_this_external_address_q_cry_4\
        );

    \I__7497\ : IoInMux
    port map (
            O => \N__31047\,
            I => \N__31044\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__31044\,
            I => \N__31041\
        );

    \I__7495\ : Span12Mux_s6_h
    port map (
            O => \N__31041\,
            I => \N__31037\
        );

    \I__7494\ : InMux
    port map (
            O => \N__31040\,
            I => \N__31034\
        );

    \I__7493\ : Odrv12
    port map (
            O => \N__31037\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__31034\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__7491\ : InMux
    port map (
            O => \N__31029\,
            I => \M_this_external_address_q_cry_5\
        );

    \I__7490\ : IoInMux
    port map (
            O => \N__31026\,
            I => \N__31023\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__31023\,
            I => \N__31020\
        );

    \I__7488\ : Span4Mux_s2_h
    port map (
            O => \N__31020\,
            I => \N__31017\
        );

    \I__7487\ : Span4Mux_h
    port map (
            O => \N__31017\,
            I => \N__31014\
        );

    \I__7486\ : Sp12to4
    port map (
            O => \N__31014\,
            I => \N__31011\
        );

    \I__7485\ : Span12Mux_v
    port map (
            O => \N__31011\,
            I => \N__31007\
        );

    \I__7484\ : InMux
    port map (
            O => \N__31010\,
            I => \N__31004\
        );

    \I__7483\ : Odrv12
    port map (
            O => \N__31007\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__31004\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__7481\ : InMux
    port map (
            O => \N__30999\,
            I => \M_this_external_address_q_cry_6\
        );

    \I__7480\ : IoInMux
    port map (
            O => \N__30996\,
            I => \N__30993\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__30993\,
            I => \N__30990\
        );

    \I__7478\ : Span4Mux_s0_v
    port map (
            O => \N__30990\,
            I => \N__30987\
        );

    \I__7477\ : Sp12to4
    port map (
            O => \N__30987\,
            I => \N__30983\
        );

    \I__7476\ : InMux
    port map (
            O => \N__30986\,
            I => \N__30980\
        );

    \I__7475\ : Span12Mux_h
    port map (
            O => \N__30983\,
            I => \N__30977\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__30980\,
            I => \N__30974\
        );

    \I__7473\ : Odrv12
    port map (
            O => \N__30977\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__7472\ : Odrv12
    port map (
            O => \N__30974\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__7471\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30966\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__30966\,
            I => \N__30963\
        );

    \I__7469\ : Span4Mux_h
    port map (
            O => \N__30963\,
            I => \N__30960\
        );

    \I__7468\ : Odrv4
    port map (
            O => \N__30960\,
            I => \M_this_external_address_q_s_8\
        );

    \I__7467\ : InMux
    port map (
            O => \N__30957\,
            I => \bfn_26_24_0_\
        );

    \I__7466\ : InMux
    port map (
            O => \N__30954\,
            I => \N__30951\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__30951\,
            I => \N__30948\
        );

    \I__7464\ : Odrv4
    port map (
            O => \N__30948\,
            I => \M_this_external_address_q_3_0_12\
        );

    \I__7463\ : InMux
    port map (
            O => \N__30945\,
            I => \N__30942\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__30942\,
            I => \N__30939\
        );

    \I__7461\ : Odrv4
    port map (
            O => \N__30939\,
            I => \M_this_external_address_q_3_14\
        );

    \I__7460\ : CascadeMux
    port map (
            O => \N__30936\,
            I => \N__30931\
        );

    \I__7459\ : InMux
    port map (
            O => \N__30935\,
            I => \N__30925\
        );

    \I__7458\ : CascadeMux
    port map (
            O => \N__30934\,
            I => \N__30922\
        );

    \I__7457\ : InMux
    port map (
            O => \N__30931\,
            I => \N__30919\
        );

    \I__7456\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30916\
        );

    \I__7455\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30910\
        );

    \I__7454\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30907\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__30925\,
            I => \N__30904\
        );

    \I__7452\ : InMux
    port map (
            O => \N__30922\,
            I => \N__30901\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__30919\,
            I => \N__30896\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__30916\,
            I => \N__30896\
        );

    \I__7449\ : CascadeMux
    port map (
            O => \N__30915\,
            I => \N__30893\
        );

    \I__7448\ : CascadeMux
    port map (
            O => \N__30914\,
            I => \N__30890\
        );

    \I__7447\ : InMux
    port map (
            O => \N__30913\,
            I => \N__30887\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__30910\,
            I => \N__30884\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__30907\,
            I => \N__30881\
        );

    \I__7444\ : Span4Mux_h
    port map (
            O => \N__30904\,
            I => \N__30876\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__30901\,
            I => \N__30876\
        );

    \I__7442\ : Span4Mux_v
    port map (
            O => \N__30896\,
            I => \N__30873\
        );

    \I__7441\ : InMux
    port map (
            O => \N__30893\,
            I => \N__30870\
        );

    \I__7440\ : InMux
    port map (
            O => \N__30890\,
            I => \N__30867\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__30887\,
            I => \N__30864\
        );

    \I__7438\ : Span4Mux_v
    port map (
            O => \N__30884\,
            I => \N__30858\
        );

    \I__7437\ : Span4Mux_h
    port map (
            O => \N__30881\,
            I => \N__30858\
        );

    \I__7436\ : Span4Mux_v
    port map (
            O => \N__30876\,
            I => \N__30855\
        );

    \I__7435\ : Span4Mux_v
    port map (
            O => \N__30873\,
            I => \N__30850\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__30870\,
            I => \N__30850\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__30867\,
            I => \N__30847\
        );

    \I__7432\ : Span4Mux_h
    port map (
            O => \N__30864\,
            I => \N__30843\
        );

    \I__7431\ : InMux
    port map (
            O => \N__30863\,
            I => \N__30840\
        );

    \I__7430\ : Span4Mux_v
    port map (
            O => \N__30858\,
            I => \N__30837\
        );

    \I__7429\ : Span4Mux_v
    port map (
            O => \N__30855\,
            I => \N__30832\
        );

    \I__7428\ : Span4Mux_v
    port map (
            O => \N__30850\,
            I => \N__30832\
        );

    \I__7427\ : Span4Mux_v
    port map (
            O => \N__30847\,
            I => \N__30829\
        );

    \I__7426\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30826\
        );

    \I__7425\ : Span4Mux_v
    port map (
            O => \N__30843\,
            I => \N__30823\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__30840\,
            I => \N__30820\
        );

    \I__7423\ : Span4Mux_v
    port map (
            O => \N__30837\,
            I => \N__30817\
        );

    \I__7422\ : Sp12to4
    port map (
            O => \N__30832\,
            I => \N__30812\
        );

    \I__7421\ : Sp12to4
    port map (
            O => \N__30829\,
            I => \N__30812\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__30826\,
            I => \N__30809\
        );

    \I__7419\ : Span4Mux_v
    port map (
            O => \N__30823\,
            I => \N__30804\
        );

    \I__7418\ : Span4Mux_h
    port map (
            O => \N__30820\,
            I => \N__30804\
        );

    \I__7417\ : Span4Mux_v
    port map (
            O => \N__30817\,
            I => \N__30801\
        );

    \I__7416\ : Span12Mux_h
    port map (
            O => \N__30812\,
            I => \N__30796\
        );

    \I__7415\ : Span12Mux_v
    port map (
            O => \N__30809\,
            I => \N__30796\
        );

    \I__7414\ : Span4Mux_v
    port map (
            O => \N__30804\,
            I => \N__30793\
        );

    \I__7413\ : Odrv4
    port map (
            O => \N__30801\,
            I => port_data_c_1
        );

    \I__7412\ : Odrv12
    port map (
            O => \N__30796\,
            I => port_data_c_1
        );

    \I__7411\ : Odrv4
    port map (
            O => \N__30793\,
            I => port_data_c_1
        );

    \I__7410\ : CEMux
    port map (
            O => \N__30786\,
            I => \N__30782\
        );

    \I__7409\ : CEMux
    port map (
            O => \N__30785\,
            I => \N__30779\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__30782\,
            I => \N__30776\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__30779\,
            I => \N__30773\
        );

    \I__7406\ : Span4Mux_v
    port map (
            O => \N__30776\,
            I => \N__30770\
        );

    \I__7405\ : Span4Mux_h
    port map (
            O => \N__30773\,
            I => \N__30767\
        );

    \I__7404\ : Odrv4
    port map (
            O => \N__30770\,
            I => \this_sprites_ram.mem_WE_2\
        );

    \I__7403\ : Odrv4
    port map (
            O => \N__30767\,
            I => \this_sprites_ram.mem_WE_2\
        );

    \I__7402\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30756\
        );

    \I__7401\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30756\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__30756\,
            I => \N__30748\
        );

    \I__7399\ : InMux
    port map (
            O => \N__30755\,
            I => \N__30745\
        );

    \I__7398\ : InMux
    port map (
            O => \N__30754\,
            I => \N__30740\
        );

    \I__7397\ : InMux
    port map (
            O => \N__30753\,
            I => \N__30740\
        );

    \I__7396\ : InMux
    port map (
            O => \N__30752\,
            I => \N__30734\
        );

    \I__7395\ : InMux
    port map (
            O => \N__30751\,
            I => \N__30734\
        );

    \I__7394\ : Span4Mux_v
    port map (
            O => \N__30748\,
            I => \N__30729\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__30745\,
            I => \N__30729\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__30740\,
            I => \N__30726\
        );

    \I__7391\ : InMux
    port map (
            O => \N__30739\,
            I => \N__30723\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__30734\,
            I => \N__30720\
        );

    \I__7389\ : Span4Mux_v
    port map (
            O => \N__30729\,
            I => \N__30713\
        );

    \I__7388\ : Span4Mux_v
    port map (
            O => \N__30726\,
            I => \N__30713\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__30723\,
            I => \N__30713\
        );

    \I__7386\ : Span4Mux_h
    port map (
            O => \N__30720\,
            I => \N__30708\
        );

    \I__7385\ : Span4Mux_h
    port map (
            O => \N__30713\,
            I => \N__30708\
        );

    \I__7384\ : Odrv4
    port map (
            O => \N__30708\,
            I => \M_this_sprites_ram_write_en_0\
        );

    \I__7383\ : CascadeMux
    port map (
            O => \N__30705\,
            I => \N__30701\
        );

    \I__7382\ : CascadeMux
    port map (
            O => \N__30704\,
            I => \N__30694\
        );

    \I__7381\ : InMux
    port map (
            O => \N__30701\,
            I => \N__30689\
        );

    \I__7380\ : InMux
    port map (
            O => \N__30700\,
            I => \N__30689\
        );

    \I__7379\ : CascadeMux
    port map (
            O => \N__30699\,
            I => \N__30686\
        );

    \I__7378\ : CascadeMux
    port map (
            O => \N__30698\,
            I => \N__30682\
        );

    \I__7377\ : CascadeMux
    port map (
            O => \N__30697\,
            I => \N__30678\
        );

    \I__7376\ : InMux
    port map (
            O => \N__30694\,
            I => \N__30674\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__30689\,
            I => \N__30671\
        );

    \I__7374\ : InMux
    port map (
            O => \N__30686\,
            I => \N__30668\
        );

    \I__7373\ : InMux
    port map (
            O => \N__30685\,
            I => \N__30663\
        );

    \I__7372\ : InMux
    port map (
            O => \N__30682\,
            I => \N__30663\
        );

    \I__7371\ : InMux
    port map (
            O => \N__30681\,
            I => \N__30658\
        );

    \I__7370\ : InMux
    port map (
            O => \N__30678\,
            I => \N__30658\
        );

    \I__7369\ : CascadeMux
    port map (
            O => \N__30677\,
            I => \N__30654\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__30674\,
            I => \N__30648\
        );

    \I__7367\ : Span4Mux_v
    port map (
            O => \N__30671\,
            I => \N__30648\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__30668\,
            I => \N__30643\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__30663\,
            I => \N__30643\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__30658\,
            I => \N__30640\
        );

    \I__7363\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30635\
        );

    \I__7362\ : InMux
    port map (
            O => \N__30654\,
            I => \N__30635\
        );

    \I__7361\ : InMux
    port map (
            O => \N__30653\,
            I => \N__30632\
        );

    \I__7360\ : Span4Mux_v
    port map (
            O => \N__30648\,
            I => \N__30627\
        );

    \I__7359\ : Span4Mux_v
    port map (
            O => \N__30643\,
            I => \N__30627\
        );

    \I__7358\ : Span4Mux_h
    port map (
            O => \N__30640\,
            I => \N__30624\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__30635\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__30632\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7355\ : Odrv4
    port map (
            O => \N__30627\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7354\ : Odrv4
    port map (
            O => \N__30624\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7353\ : CascadeMux
    port map (
            O => \N__30615\,
            I => \N__30611\
        );

    \I__7352\ : CascadeMux
    port map (
            O => \N__30614\,
            I => \N__30607\
        );

    \I__7351\ : InMux
    port map (
            O => \N__30611\,
            I => \N__30600\
        );

    \I__7350\ : InMux
    port map (
            O => \N__30610\,
            I => \N__30600\
        );

    \I__7349\ : InMux
    port map (
            O => \N__30607\,
            I => \N__30595\
        );

    \I__7348\ : InMux
    port map (
            O => \N__30606\,
            I => \N__30595\
        );

    \I__7347\ : InMux
    port map (
            O => \N__30605\,
            I => \N__30588\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__30600\,
            I => \N__30585\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__30595\,
            I => \N__30582\
        );

    \I__7344\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30577\
        );

    \I__7343\ : InMux
    port map (
            O => \N__30593\,
            I => \N__30577\
        );

    \I__7342\ : CascadeMux
    port map (
            O => \N__30592\,
            I => \N__30574\
        );

    \I__7341\ : InMux
    port map (
            O => \N__30591\,
            I => \N__30569\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__30588\,
            I => \N__30564\
        );

    \I__7339\ : Span4Mux_v
    port map (
            O => \N__30585\,
            I => \N__30564\
        );

    \I__7338\ : Span4Mux_h
    port map (
            O => \N__30582\,
            I => \N__30561\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__30577\,
            I => \N__30558\
        );

    \I__7336\ : InMux
    port map (
            O => \N__30574\,
            I => \N__30555\
        );

    \I__7335\ : InMux
    port map (
            O => \N__30573\,
            I => \N__30552\
        );

    \I__7334\ : InMux
    port map (
            O => \N__30572\,
            I => \N__30549\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__30569\,
            I => \N__30542\
        );

    \I__7332\ : Span4Mux_v
    port map (
            O => \N__30564\,
            I => \N__30542\
        );

    \I__7331\ : Span4Mux_v
    port map (
            O => \N__30561\,
            I => \N__30542\
        );

    \I__7330\ : Span4Mux_h
    port map (
            O => \N__30558\,
            I => \N__30539\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__30555\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__30552\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__30549\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7326\ : Odrv4
    port map (
            O => \N__30542\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7325\ : Odrv4
    port map (
            O => \N__30539\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7324\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30521\
        );

    \I__7323\ : InMux
    port map (
            O => \N__30527\,
            I => \N__30521\
        );

    \I__7322\ : CascadeMux
    port map (
            O => \N__30526\,
            I => \N__30516\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__30521\,
            I => \N__30510\
        );

    \I__7320\ : InMux
    port map (
            O => \N__30520\,
            I => \N__30505\
        );

    \I__7319\ : InMux
    port map (
            O => \N__30519\,
            I => \N__30505\
        );

    \I__7318\ : InMux
    port map (
            O => \N__30516\,
            I => \N__30500\
        );

    \I__7317\ : InMux
    port map (
            O => \N__30515\,
            I => \N__30500\
        );

    \I__7316\ : InMux
    port map (
            O => \N__30514\,
            I => \N__30497\
        );

    \I__7315\ : CascadeMux
    port map (
            O => \N__30513\,
            I => \N__30494\
        );

    \I__7314\ : Span4Mux_v
    port map (
            O => \N__30510\,
            I => \N__30491\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__30505\,
            I => \N__30488\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__30500\,
            I => \N__30485\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__30497\,
            I => \N__30482\
        );

    \I__7310\ : InMux
    port map (
            O => \N__30494\,
            I => \N__30477\
        );

    \I__7309\ : Span4Mux_v
    port map (
            O => \N__30491\,
            I => \N__30472\
        );

    \I__7308\ : Span4Mux_v
    port map (
            O => \N__30488\,
            I => \N__30472\
        );

    \I__7307\ : Span4Mux_h
    port map (
            O => \N__30485\,
            I => \N__30469\
        );

    \I__7306\ : Span4Mux_h
    port map (
            O => \N__30482\,
            I => \N__30466\
        );

    \I__7305\ : InMux
    port map (
            O => \N__30481\,
            I => \N__30463\
        );

    \I__7304\ : InMux
    port map (
            O => \N__30480\,
            I => \N__30460\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__30477\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7302\ : Odrv4
    port map (
            O => \N__30472\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7301\ : Odrv4
    port map (
            O => \N__30469\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7300\ : Odrv4
    port map (
            O => \N__30466\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__30463\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__30460\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7297\ : CEMux
    port map (
            O => \N__30447\,
            I => \N__30443\
        );

    \I__7296\ : CEMux
    port map (
            O => \N__30446\,
            I => \N__30440\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__30443\,
            I => \N__30435\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__30440\,
            I => \N__30435\
        );

    \I__7293\ : Span4Mux_v
    port map (
            O => \N__30435\,
            I => \N__30432\
        );

    \I__7292\ : Odrv4
    port map (
            O => \N__30432\,
            I => \this_sprites_ram.mem_WE_0\
        );

    \I__7291\ : CascadeMux
    port map (
            O => \N__30429\,
            I => \N__30426\
        );

    \I__7290\ : InMux
    port map (
            O => \N__30426\,
            I => \N__30423\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__30423\,
            I => \N__30420\
        );

    \I__7288\ : Span4Mux_v
    port map (
            O => \N__30420\,
            I => \N__30417\
        );

    \I__7287\ : Span4Mux_h
    port map (
            O => \N__30417\,
            I => \N__30414\
        );

    \I__7286\ : Span4Mux_h
    port map (
            O => \N__30414\,
            I => \N__30411\
        );

    \I__7285\ : Sp12to4
    port map (
            O => \N__30411\,
            I => \N__30408\
        );

    \I__7284\ : Odrv12
    port map (
            O => \N__30408\,
            I => \M_this_map_ram_read_data_4\
        );

    \I__7283\ : InMux
    port map (
            O => \N__30405\,
            I => \N__30402\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__30402\,
            I => \N__30399\
        );

    \I__7281\ : Span12Mux_s10_h
    port map (
            O => \N__30399\,
            I => \N__30396\
        );

    \I__7280\ : Span12Mux_v
    port map (
            O => \N__30396\,
            I => \N__30393\
        );

    \I__7279\ : Odrv12
    port map (
            O => \N__30393\,
            I => \this_ppu.un10_sprites_addr_cry_1_c_RNIOM6BZ0\
        );

    \I__7278\ : CascadeMux
    port map (
            O => \N__30390\,
            I => \N__30387\
        );

    \I__7277\ : CascadeBuf
    port map (
            O => \N__30387\,
            I => \N__30384\
        );

    \I__7276\ : CascadeMux
    port map (
            O => \N__30384\,
            I => \N__30381\
        );

    \I__7275\ : CascadeBuf
    port map (
            O => \N__30381\,
            I => \N__30378\
        );

    \I__7274\ : CascadeMux
    port map (
            O => \N__30378\,
            I => \N__30375\
        );

    \I__7273\ : CascadeBuf
    port map (
            O => \N__30375\,
            I => \N__30372\
        );

    \I__7272\ : CascadeMux
    port map (
            O => \N__30372\,
            I => \N__30369\
        );

    \I__7271\ : CascadeBuf
    port map (
            O => \N__30369\,
            I => \N__30366\
        );

    \I__7270\ : CascadeMux
    port map (
            O => \N__30366\,
            I => \N__30363\
        );

    \I__7269\ : CascadeBuf
    port map (
            O => \N__30363\,
            I => \N__30360\
        );

    \I__7268\ : CascadeMux
    port map (
            O => \N__30360\,
            I => \N__30357\
        );

    \I__7267\ : CascadeBuf
    port map (
            O => \N__30357\,
            I => \N__30354\
        );

    \I__7266\ : CascadeMux
    port map (
            O => \N__30354\,
            I => \N__30351\
        );

    \I__7265\ : CascadeBuf
    port map (
            O => \N__30351\,
            I => \N__30348\
        );

    \I__7264\ : CascadeMux
    port map (
            O => \N__30348\,
            I => \N__30345\
        );

    \I__7263\ : CascadeBuf
    port map (
            O => \N__30345\,
            I => \N__30342\
        );

    \I__7262\ : CascadeMux
    port map (
            O => \N__30342\,
            I => \N__30339\
        );

    \I__7261\ : CascadeBuf
    port map (
            O => \N__30339\,
            I => \N__30336\
        );

    \I__7260\ : CascadeMux
    port map (
            O => \N__30336\,
            I => \N__30333\
        );

    \I__7259\ : CascadeBuf
    port map (
            O => \N__30333\,
            I => \N__30330\
        );

    \I__7258\ : CascadeMux
    port map (
            O => \N__30330\,
            I => \N__30327\
        );

    \I__7257\ : CascadeBuf
    port map (
            O => \N__30327\,
            I => \N__30324\
        );

    \I__7256\ : CascadeMux
    port map (
            O => \N__30324\,
            I => \N__30321\
        );

    \I__7255\ : CascadeBuf
    port map (
            O => \N__30321\,
            I => \N__30318\
        );

    \I__7254\ : CascadeMux
    port map (
            O => \N__30318\,
            I => \N__30315\
        );

    \I__7253\ : CascadeBuf
    port map (
            O => \N__30315\,
            I => \N__30312\
        );

    \I__7252\ : CascadeMux
    port map (
            O => \N__30312\,
            I => \N__30309\
        );

    \I__7251\ : CascadeBuf
    port map (
            O => \N__30309\,
            I => \N__30306\
        );

    \I__7250\ : CascadeMux
    port map (
            O => \N__30306\,
            I => \N__30303\
        );

    \I__7249\ : CascadeBuf
    port map (
            O => \N__30303\,
            I => \N__30300\
        );

    \I__7248\ : CascadeMux
    port map (
            O => \N__30300\,
            I => \N__30297\
        );

    \I__7247\ : InMux
    port map (
            O => \N__30297\,
            I => \N__30294\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__30294\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__7245\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30288\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__30288\,
            I => \N__30285\
        );

    \I__7243\ : Span4Mux_s2_v
    port map (
            O => \N__30285\,
            I => \N__30282\
        );

    \I__7242\ : Sp12to4
    port map (
            O => \N__30282\,
            I => \N__30276\
        );

    \I__7241\ : InMux
    port map (
            O => \N__30281\,
            I => \N__30273\
        );

    \I__7240\ : CascadeMux
    port map (
            O => \N__30280\,
            I => \N__30270\
        );

    \I__7239\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30267\
        );

    \I__7238\ : Span12Mux_h
    port map (
            O => \N__30276\,
            I => \N__30264\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__30273\,
            I => \N__30261\
        );

    \I__7236\ : InMux
    port map (
            O => \N__30270\,
            I => \N__30258\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__30267\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7234\ : Odrv12
    port map (
            O => \N__30264\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7233\ : Odrv4
    port map (
            O => \N__30261\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__30258\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7231\ : InMux
    port map (
            O => \N__30249\,
            I => \N__30246\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__30246\,
            I => \N__30243\
        );

    \I__7229\ : Span12Mux_v
    port map (
            O => \N__30243\,
            I => \N__30240\
        );

    \I__7228\ : Span12Mux_h
    port map (
            O => \N__30240\,
            I => \N__30237\
        );

    \I__7227\ : Odrv12
    port map (
            O => \N__30237\,
            I => \this_ppu.un3_sprites_addr_cry_4_c_RNI32FZ0Z8\
        );

    \I__7226\ : CascadeMux
    port map (
            O => \N__30234\,
            I => \N__30231\
        );

    \I__7225\ : CascadeBuf
    port map (
            O => \N__30231\,
            I => \N__30228\
        );

    \I__7224\ : CascadeMux
    port map (
            O => \N__30228\,
            I => \N__30225\
        );

    \I__7223\ : CascadeBuf
    port map (
            O => \N__30225\,
            I => \N__30222\
        );

    \I__7222\ : CascadeMux
    port map (
            O => \N__30222\,
            I => \N__30219\
        );

    \I__7221\ : CascadeBuf
    port map (
            O => \N__30219\,
            I => \N__30216\
        );

    \I__7220\ : CascadeMux
    port map (
            O => \N__30216\,
            I => \N__30213\
        );

    \I__7219\ : CascadeBuf
    port map (
            O => \N__30213\,
            I => \N__30210\
        );

    \I__7218\ : CascadeMux
    port map (
            O => \N__30210\,
            I => \N__30207\
        );

    \I__7217\ : CascadeBuf
    port map (
            O => \N__30207\,
            I => \N__30204\
        );

    \I__7216\ : CascadeMux
    port map (
            O => \N__30204\,
            I => \N__30201\
        );

    \I__7215\ : CascadeBuf
    port map (
            O => \N__30201\,
            I => \N__30198\
        );

    \I__7214\ : CascadeMux
    port map (
            O => \N__30198\,
            I => \N__30195\
        );

    \I__7213\ : CascadeBuf
    port map (
            O => \N__30195\,
            I => \N__30192\
        );

    \I__7212\ : CascadeMux
    port map (
            O => \N__30192\,
            I => \N__30189\
        );

    \I__7211\ : CascadeBuf
    port map (
            O => \N__30189\,
            I => \N__30186\
        );

    \I__7210\ : CascadeMux
    port map (
            O => \N__30186\,
            I => \N__30183\
        );

    \I__7209\ : CascadeBuf
    port map (
            O => \N__30183\,
            I => \N__30180\
        );

    \I__7208\ : CascadeMux
    port map (
            O => \N__30180\,
            I => \N__30177\
        );

    \I__7207\ : CascadeBuf
    port map (
            O => \N__30177\,
            I => \N__30174\
        );

    \I__7206\ : CascadeMux
    port map (
            O => \N__30174\,
            I => \N__30171\
        );

    \I__7205\ : CascadeBuf
    port map (
            O => \N__30171\,
            I => \N__30168\
        );

    \I__7204\ : CascadeMux
    port map (
            O => \N__30168\,
            I => \N__30165\
        );

    \I__7203\ : CascadeBuf
    port map (
            O => \N__30165\,
            I => \N__30162\
        );

    \I__7202\ : CascadeMux
    port map (
            O => \N__30162\,
            I => \N__30159\
        );

    \I__7201\ : CascadeBuf
    port map (
            O => \N__30159\,
            I => \N__30156\
        );

    \I__7200\ : CascadeMux
    port map (
            O => \N__30156\,
            I => \N__30153\
        );

    \I__7199\ : CascadeBuf
    port map (
            O => \N__30153\,
            I => \N__30150\
        );

    \I__7198\ : CascadeMux
    port map (
            O => \N__30150\,
            I => \N__30147\
        );

    \I__7197\ : CascadeBuf
    port map (
            O => \N__30147\,
            I => \N__30144\
        );

    \I__7196\ : CascadeMux
    port map (
            O => \N__30144\,
            I => \N__30141\
        );

    \I__7195\ : InMux
    port map (
            O => \N__30141\,
            I => \N__30138\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__30138\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__7193\ : InMux
    port map (
            O => \N__30135\,
            I => \N__30132\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__30132\,
            I => \N__30129\
        );

    \I__7191\ : Span4Mux_v
    port map (
            O => \N__30129\,
            I => \N__30126\
        );

    \I__7190\ : Span4Mux_v
    port map (
            O => \N__30126\,
            I => \N__30123\
        );

    \I__7189\ : Span4Mux_v
    port map (
            O => \N__30123\,
            I => \N__30120\
        );

    \I__7188\ : Odrv4
    port map (
            O => \N__30120\,
            I => \this_sprites_ram.mem_out_bus7_3\
        );

    \I__7187\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30114\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__30114\,
            I => \N__30111\
        );

    \I__7185\ : Odrv4
    port map (
            O => \N__30111\,
            I => \this_sprites_ram.mem_out_bus3_3\
        );

    \I__7184\ : InMux
    port map (
            O => \N__30108\,
            I => \N__30102\
        );

    \I__7183\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30097\
        );

    \I__7182\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30092\
        );

    \I__7181\ : InMux
    port map (
            O => \N__30105\,
            I => \N__30085\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__30102\,
            I => \N__30082\
        );

    \I__7179\ : InMux
    port map (
            O => \N__30101\,
            I => \N__30077\
        );

    \I__7178\ : InMux
    port map (
            O => \N__30100\,
            I => \N__30077\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__30097\,
            I => \N__30073\
        );

    \I__7176\ : InMux
    port map (
            O => \N__30096\,
            I => \N__30068\
        );

    \I__7175\ : InMux
    port map (
            O => \N__30095\,
            I => \N__30068\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__30092\,
            I => \N__30065\
        );

    \I__7173\ : InMux
    port map (
            O => \N__30091\,
            I => \N__30060\
        );

    \I__7172\ : InMux
    port map (
            O => \N__30090\,
            I => \N__30060\
        );

    \I__7171\ : InMux
    port map (
            O => \N__30089\,
            I => \N__30057\
        );

    \I__7170\ : InMux
    port map (
            O => \N__30088\,
            I => \N__30053\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__30085\,
            I => \N__30050\
        );

    \I__7168\ : Span4Mux_v
    port map (
            O => \N__30082\,
            I => \N__30045\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__30077\,
            I => \N__30045\
        );

    \I__7166\ : InMux
    port map (
            O => \N__30076\,
            I => \N__30042\
        );

    \I__7165\ : Span4Mux_v
    port map (
            O => \N__30073\,
            I => \N__30037\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__30068\,
            I => \N__30037\
        );

    \I__7163\ : Span4Mux_v
    port map (
            O => \N__30065\,
            I => \N__30032\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__30060\,
            I => \N__30027\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__30057\,
            I => \N__30027\
        );

    \I__7160\ : InMux
    port map (
            O => \N__30056\,
            I => \N__30024\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__30053\,
            I => \N__30015\
        );

    \I__7158\ : Span4Mux_v
    port map (
            O => \N__30050\,
            I => \N__30015\
        );

    \I__7157\ : Span4Mux_h
    port map (
            O => \N__30045\,
            I => \N__30015\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__30042\,
            I => \N__30015\
        );

    \I__7155\ : Span4Mux_h
    port map (
            O => \N__30037\,
            I => \N__30012\
        );

    \I__7154\ : InMux
    port map (
            O => \N__30036\,
            I => \N__30007\
        );

    \I__7153\ : InMux
    port map (
            O => \N__30035\,
            I => \N__30007\
        );

    \I__7152\ : Span4Mux_v
    port map (
            O => \N__30032\,
            I => \N__30002\
        );

    \I__7151\ : Span4Mux_h
    port map (
            O => \N__30027\,
            I => \N__30002\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__30024\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7149\ : Odrv4
    port map (
            O => \N__30015\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7148\ : Odrv4
    port map (
            O => \N__30012\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__30007\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7146\ : Odrv4
    port map (
            O => \N__30002\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7145\ : InMux
    port map (
            O => \N__29991\,
            I => \N__29988\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__29988\,
            I => \N__29985\
        );

    \I__7143\ : Span4Mux_h
    port map (
            O => \N__29985\,
            I => \N__29982\
        );

    \I__7142\ : Odrv4
    port map (
            O => \N__29982\,
            I => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\
        );

    \I__7141\ : InMux
    port map (
            O => \N__29979\,
            I => \N__29976\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__29976\,
            I => \N__29973\
        );

    \I__7139\ : Odrv12
    port map (
            O => \N__29973\,
            I => \M_this_data_count_q_s_9\
        );

    \I__7138\ : InMux
    port map (
            O => \N__29970\,
            I => \M_this_data_count_q_cry_8\
        );

    \I__7137\ : CascadeMux
    port map (
            O => \N__29967\,
            I => \N__29964\
        );

    \I__7136\ : InMux
    port map (
            O => \N__29964\,
            I => \N__29961\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__29961\,
            I => \N__29956\
        );

    \I__7134\ : InMux
    port map (
            O => \N__29960\,
            I => \N__29951\
        );

    \I__7133\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29951\
        );

    \I__7132\ : Odrv4
    port map (
            O => \N__29956\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__29951\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__7130\ : InMux
    port map (
            O => \N__29946\,
            I => \N__29943\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__29943\,
            I => \M_this_data_count_q_cry_9_THRU_CO\
        );

    \I__7128\ : InMux
    port map (
            O => \N__29940\,
            I => \M_this_data_count_q_cry_9\
        );

    \I__7127\ : CascadeMux
    port map (
            O => \N__29937\,
            I => \N__29933\
        );

    \I__7126\ : InMux
    port map (
            O => \N__29936\,
            I => \N__29930\
        );

    \I__7125\ : InMux
    port map (
            O => \N__29933\,
            I => \N__29927\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__29930\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__29927\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__7122\ : InMux
    port map (
            O => \N__29922\,
            I => \N__29919\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__29919\,
            I => \M_this_data_count_q_s_11\
        );

    \I__7120\ : InMux
    port map (
            O => \N__29916\,
            I => \M_this_data_count_q_cry_10\
        );

    \I__7119\ : CascadeMux
    port map (
            O => \N__29913\,
            I => \N__29910\
        );

    \I__7118\ : InMux
    port map (
            O => \N__29910\,
            I => \N__29906\
        );

    \I__7117\ : InMux
    port map (
            O => \N__29909\,
            I => \N__29903\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__29906\,
            I => \N__29900\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__29903\,
            I => \N__29897\
        );

    \I__7114\ : Odrv4
    port map (
            O => \N__29900\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__7113\ : Odrv4
    port map (
            O => \N__29897\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__7112\ : InMux
    port map (
            O => \N__29892\,
            I => \N__29889\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__29889\,
            I => \N__29886\
        );

    \I__7110\ : Odrv4
    port map (
            O => \N__29886\,
            I => \M_this_data_count_q_s_12\
        );

    \I__7109\ : InMux
    port map (
            O => \N__29883\,
            I => \M_this_data_count_q_cry_11\
        );

    \I__7108\ : InMux
    port map (
            O => \N__29880\,
            I => \N__29876\
        );

    \I__7107\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29872\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__29876\,
            I => \N__29869\
        );

    \I__7105\ : InMux
    port map (
            O => \N__29875\,
            I => \N__29866\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__29872\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__7103\ : Odrv4
    port map (
            O => \N__29869\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__29866\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__7101\ : CascadeMux
    port map (
            O => \N__29859\,
            I => \N__29856\
        );

    \I__7100\ : InMux
    port map (
            O => \N__29856\,
            I => \N__29853\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__29853\,
            I => \N__29850\
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__29850\,
            I => \M_this_data_count_q_cry_12_THRU_CO\
        );

    \I__7097\ : InMux
    port map (
            O => \N__29847\,
            I => \M_this_data_count_q_cry_12\
        );

    \I__7096\ : SRMux
    port map (
            O => \N__29844\,
            I => \N__29838\
        );

    \I__7095\ : IoInMux
    port map (
            O => \N__29843\,
            I => \N__29832\
        );

    \I__7094\ : SRMux
    port map (
            O => \N__29842\,
            I => \N__29829\
        );

    \I__7093\ : SRMux
    port map (
            O => \N__29841\,
            I => \N__29826\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__29838\,
            I => \N__29823\
        );

    \I__7091\ : SRMux
    port map (
            O => \N__29837\,
            I => \N__29820\
        );

    \I__7090\ : SRMux
    port map (
            O => \N__29836\,
            I => \N__29816\
        );

    \I__7089\ : IoInMux
    port map (
            O => \N__29835\,
            I => \N__29813\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__29832\,
            I => \N__29809\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__29829\,
            I => \N__29804\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__29826\,
            I => \N__29804\
        );

    \I__7085\ : Span4Mux_s3_v
    port map (
            O => \N__29823\,
            I => \N__29799\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__29820\,
            I => \N__29799\
        );

    \I__7083\ : SRMux
    port map (
            O => \N__29819\,
            I => \N__29796\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__29816\,
            I => \N__29791\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__29813\,
            I => \N__29784\
        );

    \I__7080\ : SRMux
    port map (
            O => \N__29812\,
            I => \N__29781\
        );

    \I__7079\ : Span4Mux_s3_h
    port map (
            O => \N__29809\,
            I => \N__29775\
        );

    \I__7078\ : Span4Mux_v
    port map (
            O => \N__29804\,
            I => \N__29768\
        );

    \I__7077\ : Span4Mux_v
    port map (
            O => \N__29799\,
            I => \N__29768\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__29796\,
            I => \N__29768\
        );

    \I__7075\ : SRMux
    port map (
            O => \N__29795\,
            I => \N__29765\
        );

    \I__7074\ : SRMux
    port map (
            O => \N__29794\,
            I => \N__29762\
        );

    \I__7073\ : Span4Mux_v
    port map (
            O => \N__29791\,
            I => \N__29759\
        );

    \I__7072\ : SRMux
    port map (
            O => \N__29790\,
            I => \N__29756\
        );

    \I__7071\ : SRMux
    port map (
            O => \N__29789\,
            I => \N__29748\
        );

    \I__7070\ : SRMux
    port map (
            O => \N__29788\,
            I => \N__29745\
        );

    \I__7069\ : SRMux
    port map (
            O => \N__29787\,
            I => \N__29740\
        );

    \I__7068\ : IoSpan4Mux
    port map (
            O => \N__29784\,
            I => \N__29736\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__29781\,
            I => \N__29732\
        );

    \I__7066\ : SRMux
    port map (
            O => \N__29780\,
            I => \N__29729\
        );

    \I__7065\ : SRMux
    port map (
            O => \N__29779\,
            I => \N__29726\
        );

    \I__7064\ : SRMux
    port map (
            O => \N__29778\,
            I => \N__29722\
        );

    \I__7063\ : Span4Mux_h
    port map (
            O => \N__29775\,
            I => \N__29711\
        );

    \I__7062\ : Span4Mux_v
    port map (
            O => \N__29768\,
            I => \N__29711\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__29765\,
            I => \N__29711\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__29762\,
            I => \N__29711\
        );

    \I__7059\ : Span4Mux_v
    port map (
            O => \N__29759\,
            I => \N__29706\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__29756\,
            I => \N__29706\
        );

    \I__7057\ : SRMux
    port map (
            O => \N__29755\,
            I => \N__29703\
        );

    \I__7056\ : SRMux
    port map (
            O => \N__29754\,
            I => \N__29699\
        );

    \I__7055\ : CascadeMux
    port map (
            O => \N__29753\,
            I => \N__29695\
        );

    \I__7054\ : CascadeMux
    port map (
            O => \N__29752\,
            I => \N__29692\
        );

    \I__7053\ : CascadeMux
    port map (
            O => \N__29751\,
            I => \N__29686\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__29748\,
            I => \N__29671\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__29745\,
            I => \N__29671\
        );

    \I__7050\ : SRMux
    port map (
            O => \N__29744\,
            I => \N__29668\
        );

    \I__7049\ : SRMux
    port map (
            O => \N__29743\,
            I => \N__29665\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__29740\,
            I => \N__29661\
        );

    \I__7047\ : SRMux
    port map (
            O => \N__29739\,
            I => \N__29658\
        );

    \I__7046\ : Span4Mux_s2_h
    port map (
            O => \N__29736\,
            I => \N__29655\
        );

    \I__7045\ : SRMux
    port map (
            O => \N__29735\,
            I => \N__29652\
        );

    \I__7044\ : Span4Mux_h
    port map (
            O => \N__29732\,
            I => \N__29643\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__29729\,
            I => \N__29643\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__29726\,
            I => \N__29643\
        );

    \I__7041\ : SRMux
    port map (
            O => \N__29725\,
            I => \N__29640\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__29722\,
            I => \N__29637\
        );

    \I__7039\ : SRMux
    port map (
            O => \N__29721\,
            I => \N__29634\
        );

    \I__7038\ : SRMux
    port map (
            O => \N__29720\,
            I => \N__29631\
        );

    \I__7037\ : Span4Mux_v
    port map (
            O => \N__29711\,
            I => \N__29625\
        );

    \I__7036\ : Span4Mux_v
    port map (
            O => \N__29706\,
            I => \N__29620\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__29703\,
            I => \N__29620\
        );

    \I__7034\ : SRMux
    port map (
            O => \N__29702\,
            I => \N__29617\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__29699\,
            I => \N__29614\
        );

    \I__7032\ : InMux
    port map (
            O => \N__29698\,
            I => \N__29599\
        );

    \I__7031\ : InMux
    port map (
            O => \N__29695\,
            I => \N__29599\
        );

    \I__7030\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29599\
        );

    \I__7029\ : InMux
    port map (
            O => \N__29691\,
            I => \N__29599\
        );

    \I__7028\ : InMux
    port map (
            O => \N__29690\,
            I => \N__29599\
        );

    \I__7027\ : InMux
    port map (
            O => \N__29689\,
            I => \N__29599\
        );

    \I__7026\ : InMux
    port map (
            O => \N__29686\,
            I => \N__29599\
        );

    \I__7025\ : CascadeMux
    port map (
            O => \N__29685\,
            I => \N__29596\
        );

    \I__7024\ : CascadeMux
    port map (
            O => \N__29684\,
            I => \N__29593\
        );

    \I__7023\ : CascadeMux
    port map (
            O => \N__29683\,
            I => \N__29590\
        );

    \I__7022\ : CascadeMux
    port map (
            O => \N__29682\,
            I => \N__29587\
        );

    \I__7021\ : CascadeMux
    port map (
            O => \N__29681\,
            I => \N__29584\
        );

    \I__7020\ : CascadeMux
    port map (
            O => \N__29680\,
            I => \N__29581\
        );

    \I__7019\ : CascadeMux
    port map (
            O => \N__29679\,
            I => \N__29578\
        );

    \I__7018\ : CascadeMux
    port map (
            O => \N__29678\,
            I => \N__29574\
        );

    \I__7017\ : CascadeMux
    port map (
            O => \N__29677\,
            I => \N__29570\
        );

    \I__7016\ : CascadeMux
    port map (
            O => \N__29676\,
            I => \N__29566\
        );

    \I__7015\ : Span4Mux_s3_v
    port map (
            O => \N__29671\,
            I => \N__29559\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__29668\,
            I => \N__29559\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__29665\,
            I => \N__29559\
        );

    \I__7012\ : SRMux
    port map (
            O => \N__29664\,
            I => \N__29556\
        );

    \I__7011\ : Span4Mux_s3_v
    port map (
            O => \N__29661\,
            I => \N__29551\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__29658\,
            I => \N__29551\
        );

    \I__7009\ : Span4Mux_h
    port map (
            O => \N__29655\,
            I => \N__29546\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__29652\,
            I => \N__29546\
        );

    \I__7007\ : SRMux
    port map (
            O => \N__29651\,
            I => \N__29543\
        );

    \I__7006\ : SRMux
    port map (
            O => \N__29650\,
            I => \N__29540\
        );

    \I__7005\ : Span4Mux_v
    port map (
            O => \N__29643\,
            I => \N__29534\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__29640\,
            I => \N__29534\
        );

    \I__7003\ : Span4Mux_v
    port map (
            O => \N__29637\,
            I => \N__29527\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__29634\,
            I => \N__29527\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__29631\,
            I => \N__29527\
        );

    \I__7000\ : SRMux
    port map (
            O => \N__29630\,
            I => \N__29524\
        );

    \I__6999\ : SRMux
    port map (
            O => \N__29629\,
            I => \N__29521\
        );

    \I__6998\ : SRMux
    port map (
            O => \N__29628\,
            I => \N__29516\
        );

    \I__6997\ : Span4Mux_h
    port map (
            O => \N__29625\,
            I => \N__29505\
        );

    \I__6996\ : Span4Mux_h
    port map (
            O => \N__29620\,
            I => \N__29505\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__29617\,
            I => \N__29502\
        );

    \I__6994\ : Span4Mux_h
    port map (
            O => \N__29614\,
            I => \N__29497\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__29599\,
            I => \N__29497\
        );

    \I__6992\ : InMux
    port map (
            O => \N__29596\,
            I => \N__29488\
        );

    \I__6991\ : InMux
    port map (
            O => \N__29593\,
            I => \N__29488\
        );

    \I__6990\ : InMux
    port map (
            O => \N__29590\,
            I => \N__29488\
        );

    \I__6989\ : InMux
    port map (
            O => \N__29587\,
            I => \N__29488\
        );

    \I__6988\ : InMux
    port map (
            O => \N__29584\,
            I => \N__29481\
        );

    \I__6987\ : InMux
    port map (
            O => \N__29581\,
            I => \N__29481\
        );

    \I__6986\ : InMux
    port map (
            O => \N__29578\,
            I => \N__29481\
        );

    \I__6985\ : InMux
    port map (
            O => \N__29577\,
            I => \N__29468\
        );

    \I__6984\ : InMux
    port map (
            O => \N__29574\,
            I => \N__29468\
        );

    \I__6983\ : InMux
    port map (
            O => \N__29573\,
            I => \N__29468\
        );

    \I__6982\ : InMux
    port map (
            O => \N__29570\,
            I => \N__29468\
        );

    \I__6981\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29468\
        );

    \I__6980\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29468\
        );

    \I__6979\ : Span4Mux_v
    port map (
            O => \N__29559\,
            I => \N__29463\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__29556\,
            I => \N__29463\
        );

    \I__6977\ : Span4Mux_v
    port map (
            O => \N__29551\,
            I => \N__29454\
        );

    \I__6976\ : Span4Mux_h
    port map (
            O => \N__29546\,
            I => \N__29454\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__29543\,
            I => \N__29454\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__29540\,
            I => \N__29454\
        );

    \I__6973\ : SRMux
    port map (
            O => \N__29539\,
            I => \N__29451\
        );

    \I__6972\ : Span4Mux_v
    port map (
            O => \N__29534\,
            I => \N__29442\
        );

    \I__6971\ : Span4Mux_v
    port map (
            O => \N__29527\,
            I => \N__29442\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__29524\,
            I => \N__29442\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__29521\,
            I => \N__29442\
        );

    \I__6968\ : SRMux
    port map (
            O => \N__29520\,
            I => \N__29439\
        );

    \I__6967\ : SRMux
    port map (
            O => \N__29519\,
            I => \N__29436\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__29516\,
            I => \N__29433\
        );

    \I__6965\ : SRMux
    port map (
            O => \N__29515\,
            I => \N__29430\
        );

    \I__6964\ : SRMux
    port map (
            O => \N__29514\,
            I => \N__29427\
        );

    \I__6963\ : SRMux
    port map (
            O => \N__29513\,
            I => \N__29423\
        );

    \I__6962\ : SRMux
    port map (
            O => \N__29512\,
            I => \N__29420\
        );

    \I__6961\ : SRMux
    port map (
            O => \N__29511\,
            I => \N__29417\
        );

    \I__6960\ : SRMux
    port map (
            O => \N__29510\,
            I => \N__29414\
        );

    \I__6959\ : Span4Mux_h
    port map (
            O => \N__29505\,
            I => \N__29411\
        );

    \I__6958\ : Span4Mux_h
    port map (
            O => \N__29502\,
            I => \N__29402\
        );

    \I__6957\ : Span4Mux_v
    port map (
            O => \N__29497\,
            I => \N__29402\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__29488\,
            I => \N__29402\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__29481\,
            I => \N__29402\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__29468\,
            I => \N__29399\
        );

    \I__6953\ : Span4Mux_v
    port map (
            O => \N__29463\,
            I => \N__29392\
        );

    \I__6952\ : Span4Mux_v
    port map (
            O => \N__29454\,
            I => \N__29392\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__29451\,
            I => \N__29392\
        );

    \I__6950\ : Span4Mux_v
    port map (
            O => \N__29442\,
            I => \N__29385\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__29439\,
            I => \N__29385\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__29436\,
            I => \N__29385\
        );

    \I__6947\ : Span4Mux_v
    port map (
            O => \N__29433\,
            I => \N__29378\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__29430\,
            I => \N__29378\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__29427\,
            I => \N__29378\
        );

    \I__6944\ : SRMux
    port map (
            O => \N__29426\,
            I => \N__29375\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__29423\,
            I => \N__29370\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__29420\,
            I => \N__29370\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__29417\,
            I => \N__29367\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__29414\,
            I => \N__29364\
        );

    \I__6939\ : Span4Mux_h
    port map (
            O => \N__29411\,
            I => \N__29359\
        );

    \I__6938\ : Span4Mux_v
    port map (
            O => \N__29402\,
            I => \N__29359\
        );

    \I__6937\ : Span4Mux_v
    port map (
            O => \N__29399\,
            I => \N__29356\
        );

    \I__6936\ : Span4Mux_v
    port map (
            O => \N__29392\,
            I => \N__29351\
        );

    \I__6935\ : Span4Mux_v
    port map (
            O => \N__29385\,
            I => \N__29351\
        );

    \I__6934\ : Span4Mux_v
    port map (
            O => \N__29378\,
            I => \N__29344\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__29375\,
            I => \N__29344\
        );

    \I__6932\ : Span4Mux_v
    port map (
            O => \N__29370\,
            I => \N__29344\
        );

    \I__6931\ : Span12Mux_h
    port map (
            O => \N__29367\,
            I => \N__29341\
        );

    \I__6930\ : Span12Mux_h
    port map (
            O => \N__29364\,
            I => \N__29338\
        );

    \I__6929\ : Span4Mux_h
    port map (
            O => \N__29359\,
            I => \N__29335\
        );

    \I__6928\ : Span4Mux_h
    port map (
            O => \N__29356\,
            I => \N__29328\
        );

    \I__6927\ : Span4Mux_h
    port map (
            O => \N__29351\,
            I => \N__29328\
        );

    \I__6926\ : Span4Mux_h
    port map (
            O => \N__29344\,
            I => \N__29328\
        );

    \I__6925\ : Odrv12
    port map (
            O => \N__29341\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6924\ : Odrv12
    port map (
            O => \N__29338\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6923\ : Odrv4
    port map (
            O => \N__29335\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6922\ : Odrv4
    port map (
            O => \N__29328\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6921\ : CascadeMux
    port map (
            O => \N__29319\,
            I => \N__29316\
        );

    \I__6920\ : InMux
    port map (
            O => \N__29316\,
            I => \N__29312\
        );

    \I__6919\ : InMux
    port map (
            O => \N__29315\,
            I => \N__29309\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__29312\,
            I => \N__29304\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__29309\,
            I => \N__29304\
        );

    \I__6916\ : Span4Mux_h
    port map (
            O => \N__29304\,
            I => \N__29301\
        );

    \I__6915\ : Span4Mux_v
    port map (
            O => \N__29301\,
            I => \N__29298\
        );

    \I__6914\ : Odrv4
    port map (
            O => \N__29298\,
            I => \M_this_data_count_qZ0Z_14\
        );

    \I__6913\ : InMux
    port map (
            O => \N__29295\,
            I => \N__29292\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__29292\,
            I => \N__29289\
        );

    \I__6911\ : Span4Mux_h
    port map (
            O => \N__29289\,
            I => \N__29286\
        );

    \I__6910\ : Span4Mux_v
    port map (
            O => \N__29286\,
            I => \N__29283\
        );

    \I__6909\ : Span4Mux_h
    port map (
            O => \N__29283\,
            I => \N__29280\
        );

    \I__6908\ : Odrv4
    port map (
            O => \N__29280\,
            I => \M_this_data_count_q_s_14\
        );

    \I__6907\ : InMux
    port map (
            O => \N__29277\,
            I => \M_this_data_count_q_cry_13\
        );

    \I__6906\ : CascadeMux
    port map (
            O => \N__29274\,
            I => \N__29270\
        );

    \I__6905\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29267\
        );

    \I__6904\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29264\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__29267\,
            I => \M_this_data_count_qZ0Z_15\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__29264\,
            I => \M_this_data_count_qZ0Z_15\
        );

    \I__6901\ : InMux
    port map (
            O => \N__29259\,
            I => \M_this_data_count_q_cry_14\
        );

    \I__6900\ : InMux
    port map (
            O => \N__29256\,
            I => \N__29253\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__29253\,
            I => \N__29250\
        );

    \I__6898\ : Odrv4
    port map (
            O => \N__29250\,
            I => \M_this_data_count_q_s_15\
        );

    \I__6897\ : InMux
    port map (
            O => \N__29247\,
            I => \N__29244\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__29244\,
            I => \N__29241\
        );

    \I__6895\ : Odrv4
    port map (
            O => \N__29241\,
            I => \M_this_data_count_q_cry_3_THRU_CO\
        );

    \I__6894\ : CascadeMux
    port map (
            O => \N__29238\,
            I => \N__29228\
        );

    \I__6893\ : InMux
    port map (
            O => \N__29237\,
            I => \N__29220\
        );

    \I__6892\ : InMux
    port map (
            O => \N__29236\,
            I => \N__29220\
        );

    \I__6891\ : InMux
    port map (
            O => \N__29235\,
            I => \N__29213\
        );

    \I__6890\ : InMux
    port map (
            O => \N__29234\,
            I => \N__29213\
        );

    \I__6889\ : InMux
    port map (
            O => \N__29233\,
            I => \N__29213\
        );

    \I__6888\ : InMux
    port map (
            O => \N__29232\,
            I => \N__29209\
        );

    \I__6887\ : InMux
    port map (
            O => \N__29231\,
            I => \N__29202\
        );

    \I__6886\ : InMux
    port map (
            O => \N__29228\,
            I => \N__29202\
        );

    \I__6885\ : InMux
    port map (
            O => \N__29227\,
            I => \N__29202\
        );

    \I__6884\ : InMux
    port map (
            O => \N__29226\,
            I => \N__29197\
        );

    \I__6883\ : InMux
    port map (
            O => \N__29225\,
            I => \N__29197\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__29220\,
            I => \N__29189\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__29213\,
            I => \N__29189\
        );

    \I__6880\ : InMux
    port map (
            O => \N__29212\,
            I => \N__29185\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__29209\,
            I => \N__29182\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__29202\,
            I => \N__29177\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__29197\,
            I => \N__29177\
        );

    \I__6876\ : InMux
    port map (
            O => \N__29196\,
            I => \N__29170\
        );

    \I__6875\ : InMux
    port map (
            O => \N__29195\,
            I => \N__29170\
        );

    \I__6874\ : InMux
    port map (
            O => \N__29194\,
            I => \N__29170\
        );

    \I__6873\ : Span4Mux_h
    port map (
            O => \N__29189\,
            I => \N__29167\
        );

    \I__6872\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29164\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__29185\,
            I => \N__29161\
        );

    \I__6870\ : Span4Mux_v
    port map (
            O => \N__29182\,
            I => \N__29154\
        );

    \I__6869\ : Span4Mux_v
    port map (
            O => \N__29177\,
            I => \N__29154\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__29170\,
            I => \N__29154\
        );

    \I__6867\ : Span4Mux_v
    port map (
            O => \N__29167\,
            I => \N__29151\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__29164\,
            I => \N__29148\
        );

    \I__6865\ : Span4Mux_h
    port map (
            O => \N__29161\,
            I => \N__29143\
        );

    \I__6864\ : Span4Mux_h
    port map (
            O => \N__29154\,
            I => \N__29143\
        );

    \I__6863\ : Odrv4
    port map (
            O => \N__29151\,
            I => \N_33\
        );

    \I__6862\ : Odrv12
    port map (
            O => \N__29148\,
            I => \N_33\
        );

    \I__6861\ : Odrv4
    port map (
            O => \N__29143\,
            I => \N_33\
        );

    \I__6860\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29132\
        );

    \I__6859\ : InMux
    port map (
            O => \N__29135\,
            I => \N__29128\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__29132\,
            I => \N__29125\
        );

    \I__6857\ : InMux
    port map (
            O => \N__29131\,
            I => \N__29122\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__29128\,
            I => \N__29119\
        );

    \I__6855\ : Span4Mux_h
    port map (
            O => \N__29125\,
            I => \N__29116\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__29122\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__6853\ : Odrv4
    port map (
            O => \N__29119\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__6852\ : Odrv4
    port map (
            O => \N__29116\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__6851\ : CEMux
    port map (
            O => \N__29109\,
            I => \N__29105\
        );

    \I__6850\ : CEMux
    port map (
            O => \N__29108\,
            I => \N__29098\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__29105\,
            I => \N__29095\
        );

    \I__6848\ : CEMux
    port map (
            O => \N__29104\,
            I => \N__29092\
        );

    \I__6847\ : CEMux
    port map (
            O => \N__29103\,
            I => \N__29089\
        );

    \I__6846\ : CEMux
    port map (
            O => \N__29102\,
            I => \N__29086\
        );

    \I__6845\ : CEMux
    port map (
            O => \N__29101\,
            I => \N__29082\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__29098\,
            I => \N__29078\
        );

    \I__6843\ : Span4Mux_h
    port map (
            O => \N__29095\,
            I => \N__29073\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__29092\,
            I => \N__29073\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__29089\,
            I => \N__29070\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__29086\,
            I => \N__29067\
        );

    \I__6839\ : CEMux
    port map (
            O => \N__29085\,
            I => \N__29064\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__29082\,
            I => \N__29061\
        );

    \I__6837\ : CEMux
    port map (
            O => \N__29081\,
            I => \N__29058\
        );

    \I__6836\ : Span4Mux_v
    port map (
            O => \N__29078\,
            I => \N__29053\
        );

    \I__6835\ : Span4Mux_v
    port map (
            O => \N__29073\,
            I => \N__29053\
        );

    \I__6834\ : Span4Mux_h
    port map (
            O => \N__29070\,
            I => \N__29050\
        );

    \I__6833\ : Span4Mux_h
    port map (
            O => \N__29067\,
            I => \N__29045\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__29064\,
            I => \N__29045\
        );

    \I__6831\ : Span4Mux_v
    port map (
            O => \N__29061\,
            I => \N__29042\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__29058\,
            I => \N__29039\
        );

    \I__6829\ : Span4Mux_h
    port map (
            O => \N__29053\,
            I => \N__29036\
        );

    \I__6828\ : Odrv4
    port map (
            O => \N__29050\,
            I => \N_35\
        );

    \I__6827\ : Odrv4
    port map (
            O => \N__29045\,
            I => \N_35\
        );

    \I__6826\ : Odrv4
    port map (
            O => \N__29042\,
            I => \N_35\
        );

    \I__6825\ : Odrv4
    port map (
            O => \N__29039\,
            I => \N_35\
        );

    \I__6824\ : Odrv4
    port map (
            O => \N__29036\,
            I => \N_35\
        );

    \I__6823\ : InMux
    port map (
            O => \N__29025\,
            I => \M_this_data_count_q_cry_0\
        );

    \I__6822\ : InMux
    port map (
            O => \N__29022\,
            I => \N__29017\
        );

    \I__6821\ : InMux
    port map (
            O => \N__29021\,
            I => \N__29012\
        );

    \I__6820\ : InMux
    port map (
            O => \N__29020\,
            I => \N__29012\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__29017\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__29012\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__6817\ : InMux
    port map (
            O => \N__29007\,
            I => \N__29004\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__29004\,
            I => \N__29001\
        );

    \I__6815\ : Odrv4
    port map (
            O => \N__29001\,
            I => \M_this_data_count_q_cry_1_THRU_CO\
        );

    \I__6814\ : InMux
    port map (
            O => \N__28998\,
            I => \M_this_data_count_q_cry_1\
        );

    \I__6813\ : CascadeMux
    port map (
            O => \N__28995\,
            I => \N__28991\
        );

    \I__6812\ : InMux
    port map (
            O => \N__28994\,
            I => \N__28988\
        );

    \I__6811\ : InMux
    port map (
            O => \N__28991\,
            I => \N__28985\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__28988\,
            I => \N__28980\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__28985\,
            I => \N__28980\
        );

    \I__6808\ : Span4Mux_h
    port map (
            O => \N__28980\,
            I => \N__28976\
        );

    \I__6807\ : InMux
    port map (
            O => \N__28979\,
            I => \N__28973\
        );

    \I__6806\ : Span4Mux_v
    port map (
            O => \N__28976\,
            I => \N__28970\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__28973\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__6804\ : Odrv4
    port map (
            O => \N__28970\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__6803\ : InMux
    port map (
            O => \N__28965\,
            I => \N__28962\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__28962\,
            I => \N__28959\
        );

    \I__6801\ : Span4Mux_h
    port map (
            O => \N__28959\,
            I => \N__28956\
        );

    \I__6800\ : Span4Mux_h
    port map (
            O => \N__28956\,
            I => \N__28953\
        );

    \I__6799\ : Odrv4
    port map (
            O => \N__28953\,
            I => \M_this_data_count_q_cry_2_THRU_CO\
        );

    \I__6798\ : InMux
    port map (
            O => \N__28950\,
            I => \M_this_data_count_q_cry_2\
        );

    \I__6797\ : InMux
    port map (
            O => \N__28947\,
            I => \M_this_data_count_q_cry_3\
        );

    \I__6796\ : InMux
    port map (
            O => \N__28944\,
            I => \N__28941\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__28941\,
            I => \N__28936\
        );

    \I__6794\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28931\
        );

    \I__6793\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28931\
        );

    \I__6792\ : Odrv4
    port map (
            O => \N__28936\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__28931\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__6790\ : InMux
    port map (
            O => \N__28926\,
            I => \N__28923\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__28923\,
            I => \N__28920\
        );

    \I__6788\ : Odrv4
    port map (
            O => \N__28920\,
            I => \M_this_data_count_q_cry_4_THRU_CO\
        );

    \I__6787\ : InMux
    port map (
            O => \N__28917\,
            I => \M_this_data_count_q_cry_4\
        );

    \I__6786\ : InMux
    port map (
            O => \N__28914\,
            I => \N__28911\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__28911\,
            I => \N__28907\
        );

    \I__6784\ : InMux
    port map (
            O => \N__28910\,
            I => \N__28904\
        );

    \I__6783\ : Odrv4
    port map (
            O => \N__28907\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__28904\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__6781\ : InMux
    port map (
            O => \N__28899\,
            I => \N__28896\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__28896\,
            I => \N__28893\
        );

    \I__6779\ : Odrv12
    port map (
            O => \N__28893\,
            I => \M_this_data_count_q_s_6\
        );

    \I__6778\ : InMux
    port map (
            O => \N__28890\,
            I => \M_this_data_count_q_cry_5\
        );

    \I__6777\ : InMux
    port map (
            O => \N__28887\,
            I => \N__28883\
        );

    \I__6776\ : CascadeMux
    port map (
            O => \N__28886\,
            I => \N__28879\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__28883\,
            I => \N__28876\
        );

    \I__6774\ : InMux
    port map (
            O => \N__28882\,
            I => \N__28871\
        );

    \I__6773\ : InMux
    port map (
            O => \N__28879\,
            I => \N__28871\
        );

    \I__6772\ : Odrv4
    port map (
            O => \N__28876\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__28871\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__6770\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28863\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__28863\,
            I => \N__28860\
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__28860\,
            I => \M_this_data_count_q_cry_6_THRU_CO\
        );

    \I__6767\ : InMux
    port map (
            O => \N__28857\,
            I => \M_this_data_count_q_cry_6\
        );

    \I__6766\ : CascadeMux
    port map (
            O => \N__28854\,
            I => \N__28851\
        );

    \I__6765\ : InMux
    port map (
            O => \N__28851\,
            I => \N__28848\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__28848\,
            I => \N__28845\
        );

    \I__6763\ : Span4Mux_v
    port map (
            O => \N__28845\,
            I => \N__28841\
        );

    \I__6762\ : InMux
    port map (
            O => \N__28844\,
            I => \N__28838\
        );

    \I__6761\ : Odrv4
    port map (
            O => \N__28841\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__28838\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__6759\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28830\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__28830\,
            I => \N__28827\
        );

    \I__6757\ : Odrv4
    port map (
            O => \N__28827\,
            I => \M_this_data_count_q_s_8\
        );

    \I__6756\ : InMux
    port map (
            O => \N__28824\,
            I => \bfn_24_22_0_\
        );

    \I__6755\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28818\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__28818\,
            I => \N__28814\
        );

    \I__6753\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28811\
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__28814\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__28811\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__6750\ : InMux
    port map (
            O => \N__28806\,
            I => \N__28803\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__28803\,
            I => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\
        );

    \I__6748\ : CascadeMux
    port map (
            O => \N__28800\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\
        );

    \I__6747\ : InMux
    port map (
            O => \N__28797\,
            I => \N__28794\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__28794\,
            I => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\
        );

    \I__6745\ : InMux
    port map (
            O => \N__28791\,
            I => \N__28787\
        );

    \I__6744\ : InMux
    port map (
            O => \N__28790\,
            I => \N__28784\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__28787\,
            I => \N__28780\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__28784\,
            I => \N__28777\
        );

    \I__6741\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28774\
        );

    \I__6740\ : Span4Mux_v
    port map (
            O => \N__28780\,
            I => \N__28771\
        );

    \I__6739\ : Span12Mux_s11_h
    port map (
            O => \N__28777\,
            I => \N__28766\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__28774\,
            I => \N__28766\
        );

    \I__6737\ : Sp12to4
    port map (
            O => \N__28771\,
            I => \N__28761\
        );

    \I__6736\ : Span12Mux_v
    port map (
            O => \N__28766\,
            I => \N__28761\
        );

    \I__6735\ : Span12Mux_h
    port map (
            O => \N__28761\,
            I => \N__28758\
        );

    \I__6734\ : Odrv12
    port map (
            O => \N__28758\,
            I => \M_this_ppu_vram_data_3\
        );

    \I__6733\ : InMux
    port map (
            O => \N__28755\,
            I => \N__28752\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__28752\,
            I => \N__28749\
        );

    \I__6731\ : Span4Mux_v
    port map (
            O => \N__28749\,
            I => \N__28746\
        );

    \I__6730\ : Odrv4
    port map (
            O => \N__28746\,
            I => \this_sprites_ram.mem_out_bus6_0\
        );

    \I__6729\ : InMux
    port map (
            O => \N__28743\,
            I => \N__28740\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__28740\,
            I => \N__28737\
        );

    \I__6727\ : Span4Mux_v
    port map (
            O => \N__28737\,
            I => \N__28734\
        );

    \I__6726\ : Span4Mux_v
    port map (
            O => \N__28734\,
            I => \N__28731\
        );

    \I__6725\ : Odrv4
    port map (
            O => \N__28731\,
            I => \this_sprites_ram.mem_out_bus2_0\
        );

    \I__6724\ : CascadeMux
    port map (
            O => \N__28728\,
            I => \N__28724\
        );

    \I__6723\ : InMux
    port map (
            O => \N__28727\,
            I => \N__28721\
        );

    \I__6722\ : InMux
    port map (
            O => \N__28724\,
            I => \N__28716\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__28721\,
            I => \N__28713\
        );

    \I__6720\ : InMux
    port map (
            O => \N__28720\,
            I => \N__28710\
        );

    \I__6719\ : InMux
    port map (
            O => \N__28719\,
            I => \N__28707\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__28716\,
            I => \N__28702\
        );

    \I__6717\ : Span4Mux_v
    port map (
            O => \N__28713\,
            I => \N__28702\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__28710\,
            I => \N__28699\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__28707\,
            I => \N__28692\
        );

    \I__6714\ : Span4Mux_h
    port map (
            O => \N__28702\,
            I => \N__28692\
        );

    \I__6713\ : Span4Mux_h
    port map (
            O => \N__28699\,
            I => \N__28692\
        );

    \I__6712\ : Span4Mux_h
    port map (
            O => \N__28692\,
            I => \N__28689\
        );

    \I__6711\ : Odrv4
    port map (
            O => \N__28689\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__6710\ : InMux
    port map (
            O => \N__28686\,
            I => \N__28683\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__28683\,
            I => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0\
        );

    \I__6708\ : CascadeMux
    port map (
            O => \N__28680\,
            I => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0_cascade_\
        );

    \I__6707\ : CascadeMux
    port map (
            O => \N__28677\,
            I => \N__28673\
        );

    \I__6706\ : InMux
    port map (
            O => \N__28676\,
            I => \N__28670\
        );

    \I__6705\ : InMux
    port map (
            O => \N__28673\,
            I => \N__28663\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__28670\,
            I => \N__28658\
        );

    \I__6703\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28653\
        );

    \I__6702\ : InMux
    port map (
            O => \N__28668\,
            I => \N__28653\
        );

    \I__6701\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28648\
        );

    \I__6700\ : InMux
    port map (
            O => \N__28666\,
            I => \N__28648\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__28663\,
            I => \N__28645\
        );

    \I__6698\ : InMux
    port map (
            O => \N__28662\,
            I => \N__28640\
        );

    \I__6697\ : InMux
    port map (
            O => \N__28661\,
            I => \N__28640\
        );

    \I__6696\ : Sp12to4
    port map (
            O => \N__28658\,
            I => \N__28633\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__28653\,
            I => \N__28633\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__28648\,
            I => \N__28633\
        );

    \I__6693\ : Odrv12
    port map (
            O => \N__28645\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__28640\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__6691\ : Odrv12
    port map (
            O => \N__28633\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__6690\ : InMux
    port map (
            O => \N__28626\,
            I => \N__28623\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__28623\,
            I => \N__28620\
        );

    \I__6688\ : Span12Mux_h
    port map (
            O => \N__28620\,
            I => \N__28617\
        );

    \I__6687\ : Odrv12
    port map (
            O => \N__28617\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0\
        );

    \I__6686\ : InMux
    port map (
            O => \N__28614\,
            I => \N__28611\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__28611\,
            I => \N__28608\
        );

    \I__6684\ : Sp12to4
    port map (
            O => \N__28608\,
            I => \N__28605\
        );

    \I__6683\ : Odrv12
    port map (
            O => \N__28605\,
            I => \this_sprites_ram.mem_out_bus6_2\
        );

    \I__6682\ : InMux
    port map (
            O => \N__28602\,
            I => \N__28599\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__28599\,
            I => \N__28596\
        );

    \I__6680\ : Span4Mux_v
    port map (
            O => \N__28596\,
            I => \N__28593\
        );

    \I__6679\ : Span4Mux_v
    port map (
            O => \N__28593\,
            I => \N__28590\
        );

    \I__6678\ : Odrv4
    port map (
            O => \N__28590\,
            I => \this_sprites_ram.mem_out_bus2_2\
        );

    \I__6677\ : InMux
    port map (
            O => \N__28587\,
            I => \N__28584\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__28584\,
            I => \N__28581\
        );

    \I__6675\ : Span4Mux_v
    port map (
            O => \N__28581\,
            I => \N__28578\
        );

    \I__6674\ : Span4Mux_h
    port map (
            O => \N__28578\,
            I => \N__28575\
        );

    \I__6673\ : Odrv4
    port map (
            O => \N__28575\,
            I => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0\
        );

    \I__6672\ : CEMux
    port map (
            O => \N__28572\,
            I => \N__28568\
        );

    \I__6671\ : CEMux
    port map (
            O => \N__28571\,
            I => \N__28565\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__28568\,
            I => \N__28560\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__28565\,
            I => \N__28560\
        );

    \I__6668\ : Span4Mux_v
    port map (
            O => \N__28560\,
            I => \N__28557\
        );

    \I__6667\ : Odrv4
    port map (
            O => \N__28557\,
            I => \this_sprites_ram.mem_WE_4\
        );

    \I__6666\ : InMux
    port map (
            O => \N__28554\,
            I => \N__28551\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__28551\,
            I => \N__28548\
        );

    \I__6664\ : Span4Mux_v
    port map (
            O => \N__28548\,
            I => \N__28545\
        );

    \I__6663\ : Span4Mux_v
    port map (
            O => \N__28545\,
            I => \N__28542\
        );

    \I__6662\ : Odrv4
    port map (
            O => \N__28542\,
            I => \this_sprites_ram.mem_out_bus7_0\
        );

    \I__6661\ : InMux
    port map (
            O => \N__28539\,
            I => \N__28536\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__28536\,
            I => \N__28533\
        );

    \I__6659\ : Span4Mux_v
    port map (
            O => \N__28533\,
            I => \N__28530\
        );

    \I__6658\ : Odrv4
    port map (
            O => \N__28530\,
            I => \this_sprites_ram.mem_out_bus3_0\
        );

    \I__6657\ : InMux
    port map (
            O => \N__28527\,
            I => \N__28524\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28521\
        );

    \I__6655\ : Span12Mux_v
    port map (
            O => \N__28521\,
            I => \N__28518\
        );

    \I__6654\ : Span12Mux_h
    port map (
            O => \N__28518\,
            I => \N__28515\
        );

    \I__6653\ : Odrv12
    port map (
            O => \N__28515\,
            I => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\
        );

    \I__6652\ : InMux
    port map (
            O => \N__28512\,
            I => \N__28507\
        );

    \I__6651\ : InMux
    port map (
            O => \N__28511\,
            I => \N__28504\
        );

    \I__6650\ : InMux
    port map (
            O => \N__28510\,
            I => \N__28501\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__28507\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__28504\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__28501\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__6646\ : InMux
    port map (
            O => \N__28494\,
            I => \N__28489\
        );

    \I__6645\ : InMux
    port map (
            O => \N__28493\,
            I => \N__28484\
        );

    \I__6644\ : InMux
    port map (
            O => \N__28492\,
            I => \N__28484\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__28489\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__28484\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__6641\ : InMux
    port map (
            O => \N__28479\,
            I => \N__28476\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__28476\,
            I => \M_this_data_count_q_cry_0_THRU_CO\
        );

    \I__6639\ : InMux
    port map (
            O => \N__28473\,
            I => \N__28465\
        );

    \I__6638\ : InMux
    port map (
            O => \N__28472\,
            I => \N__28462\
        );

    \I__6637\ : InMux
    port map (
            O => \N__28471\,
            I => \N__28459\
        );

    \I__6636\ : CascadeMux
    port map (
            O => \N__28470\,
            I => \N__28456\
        );

    \I__6635\ : InMux
    port map (
            O => \N__28469\,
            I => \N__28451\
        );

    \I__6634\ : InMux
    port map (
            O => \N__28468\,
            I => \N__28448\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__28465\,
            I => \N__28444\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__28462\,
            I => \N__28441\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__28459\,
            I => \N__28438\
        );

    \I__6630\ : InMux
    port map (
            O => \N__28456\,
            I => \N__28435\
        );

    \I__6629\ : CascadeMux
    port map (
            O => \N__28455\,
            I => \N__28432\
        );

    \I__6628\ : InMux
    port map (
            O => \N__28454\,
            I => \N__28429\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__28451\,
            I => \N__28426\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__28448\,
            I => \N__28423\
        );

    \I__6625\ : InMux
    port map (
            O => \N__28447\,
            I => \N__28420\
        );

    \I__6624\ : Span4Mux_v
    port map (
            O => \N__28444\,
            I => \N__28416\
        );

    \I__6623\ : Span4Mux_v
    port map (
            O => \N__28441\,
            I => \N__28409\
        );

    \I__6622\ : Span4Mux_v
    port map (
            O => \N__28438\,
            I => \N__28409\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__28435\,
            I => \N__28409\
        );

    \I__6620\ : InMux
    port map (
            O => \N__28432\,
            I => \N__28406\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__28429\,
            I => \N__28403\
        );

    \I__6618\ : Span4Mux_v
    port map (
            O => \N__28426\,
            I => \N__28396\
        );

    \I__6617\ : Span4Mux_v
    port map (
            O => \N__28423\,
            I => \N__28396\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__28420\,
            I => \N__28396\
        );

    \I__6615\ : InMux
    port map (
            O => \N__28419\,
            I => \N__28392\
        );

    \I__6614\ : Span4Mux_v
    port map (
            O => \N__28416\,
            I => \N__28389\
        );

    \I__6613\ : Span4Mux_v
    port map (
            O => \N__28409\,
            I => \N__28386\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__28406\,
            I => \N__28383\
        );

    \I__6611\ : Span4Mux_v
    port map (
            O => \N__28403\,
            I => \N__28378\
        );

    \I__6610\ : Span4Mux_h
    port map (
            O => \N__28396\,
            I => \N__28378\
        );

    \I__6609\ : InMux
    port map (
            O => \N__28395\,
            I => \N__28375\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__28392\,
            I => \N__28372\
        );

    \I__6607\ : Span4Mux_v
    port map (
            O => \N__28389\,
            I => \N__28369\
        );

    \I__6606\ : Span4Mux_v
    port map (
            O => \N__28386\,
            I => \N__28364\
        );

    \I__6605\ : Span4Mux_v
    port map (
            O => \N__28383\,
            I => \N__28364\
        );

    \I__6604\ : Span4Mux_v
    port map (
            O => \N__28378\,
            I => \N__28361\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__28375\,
            I => \N__28358\
        );

    \I__6602\ : Span12Mux_h
    port map (
            O => \N__28372\,
            I => \N__28355\
        );

    \I__6601\ : Sp12to4
    port map (
            O => \N__28369\,
            I => \N__28350\
        );

    \I__6600\ : Sp12to4
    port map (
            O => \N__28364\,
            I => \N__28350\
        );

    \I__6599\ : Span4Mux_v
    port map (
            O => \N__28361\,
            I => \N__28347\
        );

    \I__6598\ : Span4Mux_h
    port map (
            O => \N__28358\,
            I => \N__28344\
        );

    \I__6597\ : Span12Mux_v
    port map (
            O => \N__28355\,
            I => \N__28339\
        );

    \I__6596\ : Span12Mux_h
    port map (
            O => \N__28350\,
            I => \N__28339\
        );

    \I__6595\ : Span4Mux_v
    port map (
            O => \N__28347\,
            I => \N__28336\
        );

    \I__6594\ : Span4Mux_v
    port map (
            O => \N__28344\,
            I => \N__28333\
        );

    \I__6593\ : Odrv12
    port map (
            O => \N__28339\,
            I => port_data_c_0
        );

    \I__6592\ : Odrv4
    port map (
            O => \N__28336\,
            I => port_data_c_0
        );

    \I__6591\ : Odrv4
    port map (
            O => \N__28333\,
            I => port_data_c_0
        );

    \I__6590\ : InMux
    port map (
            O => \N__28326\,
            I => \N__28321\
        );

    \I__6589\ : InMux
    port map (
            O => \N__28325\,
            I => \N__28317\
        );

    \I__6588\ : InMux
    port map (
            O => \N__28324\,
            I => \N__28314\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__28321\,
            I => \N__28311\
        );

    \I__6586\ : CascadeMux
    port map (
            O => \N__28320\,
            I => \N__28308\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__28317\,
            I => \N__28303\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__28314\,
            I => \N__28303\
        );

    \I__6583\ : Span4Mux_v
    port map (
            O => \N__28311\,
            I => \N__28298\
        );

    \I__6582\ : InMux
    port map (
            O => \N__28308\,
            I => \N__28295\
        );

    \I__6581\ : Span4Mux_h
    port map (
            O => \N__28303\,
            I => \N__28291\
        );

    \I__6580\ : InMux
    port map (
            O => \N__28302\,
            I => \N__28286\
        );

    \I__6579\ : InMux
    port map (
            O => \N__28301\,
            I => \N__28286\
        );

    \I__6578\ : Span4Mux_h
    port map (
            O => \N__28298\,
            I => \N__28282\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__28295\,
            I => \N__28279\
        );

    \I__6576\ : CascadeMux
    port map (
            O => \N__28294\,
            I => \N__28276\
        );

    \I__6575\ : Span4Mux_h
    port map (
            O => \N__28291\,
            I => \N__28270\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__28286\,
            I => \N__28270\
        );

    \I__6573\ : InMux
    port map (
            O => \N__28285\,
            I => \N__28267\
        );

    \I__6572\ : Span4Mux_h
    port map (
            O => \N__28282\,
            I => \N__28263\
        );

    \I__6571\ : Span4Mux_h
    port map (
            O => \N__28279\,
            I => \N__28260\
        );

    \I__6570\ : InMux
    port map (
            O => \N__28276\,
            I => \N__28257\
        );

    \I__6569\ : CascadeMux
    port map (
            O => \N__28275\,
            I => \N__28254\
        );

    \I__6568\ : Span4Mux_h
    port map (
            O => \N__28270\,
            I => \N__28249\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__28267\,
            I => \N__28249\
        );

    \I__6566\ : InMux
    port map (
            O => \N__28266\,
            I => \N__28246\
        );

    \I__6565\ : Span4Mux_h
    port map (
            O => \N__28263\,
            I => \N__28238\
        );

    \I__6564\ : Span4Mux_v
    port map (
            O => \N__28260\,
            I => \N__28238\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__28257\,
            I => \N__28238\
        );

    \I__6562\ : InMux
    port map (
            O => \N__28254\,
            I => \N__28235\
        );

    \I__6561\ : Span4Mux_h
    port map (
            O => \N__28249\,
            I => \N__28232\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__28246\,
            I => \N__28229\
        );

    \I__6559\ : InMux
    port map (
            O => \N__28245\,
            I => \N__28226\
        );

    \I__6558\ : Span4Mux_v
    port map (
            O => \N__28238\,
            I => \N__28223\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__28235\,
            I => \N__28220\
        );

    \I__6556\ : Sp12to4
    port map (
            O => \N__28232\,
            I => \N__28217\
        );

    \I__6555\ : Span12Mux_v
    port map (
            O => \N__28229\,
            I => \N__28212\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__28226\,
            I => \N__28212\
        );

    \I__6553\ : Span4Mux_v
    port map (
            O => \N__28223\,
            I => \N__28209\
        );

    \I__6552\ : Span4Mux_v
    port map (
            O => \N__28220\,
            I => \N__28206\
        );

    \I__6551\ : Span12Mux_v
    port map (
            O => \N__28217\,
            I => \N__28203\
        );

    \I__6550\ : Span12Mux_h
    port map (
            O => \N__28212\,
            I => \N__28196\
        );

    \I__6549\ : Sp12to4
    port map (
            O => \N__28209\,
            I => \N__28196\
        );

    \I__6548\ : Sp12to4
    port map (
            O => \N__28206\,
            I => \N__28196\
        );

    \I__6547\ : Odrv12
    port map (
            O => \N__28203\,
            I => port_data_c_4
        );

    \I__6546\ : Odrv12
    port map (
            O => \N__28196\,
            I => port_data_c_4
        );

    \I__6545\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28186\
        );

    \I__6544\ : InMux
    port map (
            O => \N__28190\,
            I => \N__28183\
        );

    \I__6543\ : InMux
    port map (
            O => \N__28189\,
            I => \N__28180\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__28186\,
            I => \N__28176\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__28183\,
            I => \N__28171\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__28180\,
            I => \N__28171\
        );

    \I__6539\ : InMux
    port map (
            O => \N__28179\,
            I => \N__28168\
        );

    \I__6538\ : Span4Mux_v
    port map (
            O => \N__28176\,
            I => \N__28163\
        );

    \I__6537\ : Span4Mux_v
    port map (
            O => \N__28171\,
            I => \N__28158\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__28168\,
            I => \N__28158\
        );

    \I__6535\ : CascadeMux
    port map (
            O => \N__28167\,
            I => \N__28155\
        );

    \I__6534\ : CascadeMux
    port map (
            O => \N__28166\,
            I => \N__28152\
        );

    \I__6533\ : Span4Mux_h
    port map (
            O => \N__28163\,
            I => \N__28149\
        );

    \I__6532\ : Span4Mux_h
    port map (
            O => \N__28158\,
            I => \N__28145\
        );

    \I__6531\ : InMux
    port map (
            O => \N__28155\,
            I => \N__28142\
        );

    \I__6530\ : InMux
    port map (
            O => \N__28152\,
            I => \N__28139\
        );

    \I__6529\ : Span4Mux_v
    port map (
            O => \N__28149\,
            I => \N__28136\
        );

    \I__6528\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28133\
        );

    \I__6527\ : Span4Mux_h
    port map (
            O => \N__28145\,
            I => \N__28128\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__28142\,
            I => \N__28128\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__28139\,
            I => \N__28124\
        );

    \I__6524\ : Span4Mux_v
    port map (
            O => \N__28136\,
            I => \N__28119\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__28133\,
            I => \N__28119\
        );

    \I__6522\ : Span4Mux_v
    port map (
            O => \N__28128\,
            I => \N__28116\
        );

    \I__6521\ : InMux
    port map (
            O => \N__28127\,
            I => \N__28113\
        );

    \I__6520\ : Span4Mux_v
    port map (
            O => \N__28124\,
            I => \N__28110\
        );

    \I__6519\ : Span4Mux_v
    port map (
            O => \N__28119\,
            I => \N__28105\
        );

    \I__6518\ : Span4Mux_h
    port map (
            O => \N__28116\,
            I => \N__28100\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__28113\,
            I => \N__28100\
        );

    \I__6516\ : Span4Mux_h
    port map (
            O => \N__28110\,
            I => \N__28097\
        );

    \I__6515\ : InMux
    port map (
            O => \N__28109\,
            I => \N__28093\
        );

    \I__6514\ : CascadeMux
    port map (
            O => \N__28108\,
            I => \N__28090\
        );

    \I__6513\ : Span4Mux_v
    port map (
            O => \N__28105\,
            I => \N__28087\
        );

    \I__6512\ : Span4Mux_v
    port map (
            O => \N__28100\,
            I => \N__28084\
        );

    \I__6511\ : Sp12to4
    port map (
            O => \N__28097\,
            I => \N__28081\
        );

    \I__6510\ : InMux
    port map (
            O => \N__28096\,
            I => \N__28078\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__28093\,
            I => \N__28075\
        );

    \I__6508\ : InMux
    port map (
            O => \N__28090\,
            I => \N__28072\
        );

    \I__6507\ : Sp12to4
    port map (
            O => \N__28087\,
            I => \N__28069\
        );

    \I__6506\ : Span4Mux_v
    port map (
            O => \N__28084\,
            I => \N__28066\
        );

    \I__6505\ : Span12Mux_s8_h
    port map (
            O => \N__28081\,
            I => \N__28057\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__28078\,
            I => \N__28057\
        );

    \I__6503\ : Sp12to4
    port map (
            O => \N__28075\,
            I => \N__28057\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__28072\,
            I => \N__28057\
        );

    \I__6501\ : Span12Mux_h
    port map (
            O => \N__28069\,
            I => \N__28050\
        );

    \I__6500\ : Sp12to4
    port map (
            O => \N__28066\,
            I => \N__28050\
        );

    \I__6499\ : Span12Mux_v
    port map (
            O => \N__28057\,
            I => \N__28050\
        );

    \I__6498\ : Odrv12
    port map (
            O => \N__28050\,
            I => port_data_c_6
        );

    \I__6497\ : CascadeMux
    port map (
            O => \N__28047\,
            I => \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_3Z0Z_0_cascade_\
        );

    \I__6496\ : CascadeMux
    port map (
            O => \N__28044\,
            I => \N__28041\
        );

    \I__6495\ : InMux
    port map (
            O => \N__28041\,
            I => \N__28037\
        );

    \I__6494\ : CascadeMux
    port map (
            O => \N__28040\,
            I => \N__28033\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__28037\,
            I => \N__28029\
        );

    \I__6492\ : InMux
    port map (
            O => \N__28036\,
            I => \N__28026\
        );

    \I__6491\ : InMux
    port map (
            O => \N__28033\,
            I => \N__28023\
        );

    \I__6490\ : InMux
    port map (
            O => \N__28032\,
            I => \N__28020\
        );

    \I__6489\ : Span4Mux_v
    port map (
            O => \N__28029\,
            I => \N__28015\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__28026\,
            I => \N__28015\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__28023\,
            I => \N__28011\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__28020\,
            I => \N__28008\
        );

    \I__6485\ : Span4Mux_v
    port map (
            O => \N__28015\,
            I => \N__28005\
        );

    \I__6484\ : InMux
    port map (
            O => \N__28014\,
            I => \N__28002\
        );

    \I__6483\ : Span4Mux_v
    port map (
            O => \N__28011\,
            I => \N__27999\
        );

    \I__6482\ : Span4Mux_h
    port map (
            O => \N__28008\,
            I => \N__27996\
        );

    \I__6481\ : Sp12to4
    port map (
            O => \N__28005\,
            I => \N__27991\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__28002\,
            I => \N__27991\
        );

    \I__6479\ : Odrv4
    port map (
            O => \N__27999\,
            I => \this_start_data_delay.N_902_0\
        );

    \I__6478\ : Odrv4
    port map (
            O => \N__27996\,
            I => \this_start_data_delay.N_902_0\
        );

    \I__6477\ : Odrv12
    port map (
            O => \N__27991\,
            I => \this_start_data_delay.N_902_0\
        );

    \I__6476\ : InMux
    port map (
            O => \N__27984\,
            I => \N__27981\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__27981\,
            I => \N__27975\
        );

    \I__6474\ : InMux
    port map (
            O => \N__27980\,
            I => \N__27972\
        );

    \I__6473\ : InMux
    port map (
            O => \N__27979\,
            I => \N__27969\
        );

    \I__6472\ : InMux
    port map (
            O => \N__27978\,
            I => \N__27966\
        );

    \I__6471\ : Span4Mux_h
    port map (
            O => \N__27975\,
            I => \N__27963\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__27972\,
            I => \N__27960\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__27969\,
            I => \N__27957\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__27966\,
            I => \N__27954\
        );

    \I__6467\ : Odrv4
    port map (
            O => \N__27963\,
            I => \this_start_data_delay.N_821_0\
        );

    \I__6466\ : Odrv4
    port map (
            O => \N__27960\,
            I => \this_start_data_delay.N_821_0\
        );

    \I__6465\ : Odrv4
    port map (
            O => \N__27957\,
            I => \this_start_data_delay.N_821_0\
        );

    \I__6464\ : Odrv4
    port map (
            O => \N__27954\,
            I => \this_start_data_delay.N_821_0\
        );

    \I__6463\ : InMux
    port map (
            O => \N__27945\,
            I => \N__27942\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__27942\,
            I => \N__27938\
        );

    \I__6461\ : CascadeMux
    port map (
            O => \N__27941\,
            I => \N__27934\
        );

    \I__6460\ : Span4Mux_h
    port map (
            O => \N__27938\,
            I => \N__27930\
        );

    \I__6459\ : InMux
    port map (
            O => \N__27937\,
            I => \N__27926\
        );

    \I__6458\ : InMux
    port map (
            O => \N__27934\,
            I => \N__27923\
        );

    \I__6457\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27920\
        );

    \I__6456\ : Span4Mux_h
    port map (
            O => \N__27930\,
            I => \N__27917\
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__27929\,
            I => \N__27913\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27908\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__27923\,
            I => \N__27902\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__27920\,
            I => \N__27902\
        );

    \I__6451\ : Span4Mux_h
    port map (
            O => \N__27917\,
            I => \N__27899\
        );

    \I__6450\ : InMux
    port map (
            O => \N__27916\,
            I => \N__27894\
        );

    \I__6449\ : InMux
    port map (
            O => \N__27913\,
            I => \N__27894\
        );

    \I__6448\ : InMux
    port map (
            O => \N__27912\,
            I => \N__27891\
        );

    \I__6447\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27888\
        );

    \I__6446\ : Span4Mux_h
    port map (
            O => \N__27908\,
            I => \N__27885\
        );

    \I__6445\ : InMux
    port map (
            O => \N__27907\,
            I => \N__27882\
        );

    \I__6444\ : Span4Mux_v
    port map (
            O => \N__27902\,
            I => \N__27879\
        );

    \I__6443\ : Span4Mux_h
    port map (
            O => \N__27899\,
            I => \N__27874\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__27894\,
            I => \N__27874\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__27891\,
            I => \N__27865\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__27888\,
            I => \N__27865\
        );

    \I__6439\ : Sp12to4
    port map (
            O => \N__27885\,
            I => \N__27865\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__27882\,
            I => \N__27865\
        );

    \I__6437\ : Sp12to4
    port map (
            O => \N__27879\,
            I => \N__27862\
        );

    \I__6436\ : Span4Mux_v
    port map (
            O => \N__27874\,
            I => \N__27859\
        );

    \I__6435\ : Span12Mux_v
    port map (
            O => \N__27865\,
            I => \N__27856\
        );

    \I__6434\ : Span12Mux_h
    port map (
            O => \N__27862\,
            I => \N__27853\
        );

    \I__6433\ : Span4Mux_h
    port map (
            O => \N__27859\,
            I => \N__27850\
        );

    \I__6432\ : Span12Mux_h
    port map (
            O => \N__27856\,
            I => \N__27847\
        );

    \I__6431\ : Span12Mux_v
    port map (
            O => \N__27853\,
            I => \N__27844\
        );

    \I__6430\ : IoSpan4Mux
    port map (
            O => \N__27850\,
            I => \N__27841\
        );

    \I__6429\ : Odrv12
    port map (
            O => \N__27847\,
            I => port_data_c_7
        );

    \I__6428\ : Odrv12
    port map (
            O => \N__27844\,
            I => port_data_c_7
        );

    \I__6427\ : Odrv4
    port map (
            O => \N__27841\,
            I => port_data_c_7
        );

    \I__6426\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27831\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__27831\,
            I => \N__27827\
        );

    \I__6424\ : InMux
    port map (
            O => \N__27830\,
            I => \N__27824\
        );

    \I__6423\ : Span4Mux_v
    port map (
            O => \N__27827\,
            I => \N__27817\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__27824\,
            I => \N__27817\
        );

    \I__6421\ : InMux
    port map (
            O => \N__27823\,
            I => \N__27814\
        );

    \I__6420\ : InMux
    port map (
            O => \N__27822\,
            I => \N__27811\
        );

    \I__6419\ : Odrv4
    port map (
            O => \N__27817\,
            I => \this_start_data_delay.N_123\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__27814\,
            I => \this_start_data_delay.N_123\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__27811\,
            I => \this_start_data_delay.N_123\
        );

    \I__6416\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27800\
        );

    \I__6415\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27796\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__27800\,
            I => \N__27792\
        );

    \I__6413\ : InMux
    port map (
            O => \N__27799\,
            I => \N__27789\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__27796\,
            I => \N__27785\
        );

    \I__6411\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27782\
        );

    \I__6410\ : Span4Mux_v
    port map (
            O => \N__27792\,
            I => \N__27776\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__27789\,
            I => \N__27776\
        );

    \I__6408\ : InMux
    port map (
            O => \N__27788\,
            I => \N__27773\
        );

    \I__6407\ : Span4Mux_v
    port map (
            O => \N__27785\,
            I => \N__27767\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__27782\,
            I => \N__27767\
        );

    \I__6405\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27764\
        );

    \I__6404\ : Span4Mux_v
    port map (
            O => \N__27776\,
            I => \N__27758\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__27773\,
            I => \N__27758\
        );

    \I__6402\ : InMux
    port map (
            O => \N__27772\,
            I => \N__27755\
        );

    \I__6401\ : Span4Mux_v
    port map (
            O => \N__27767\,
            I => \N__27750\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__27764\,
            I => \N__27750\
        );

    \I__6399\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27747\
        );

    \I__6398\ : Span4Mux_v
    port map (
            O => \N__27758\,
            I => \N__27742\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__27755\,
            I => \N__27742\
        );

    \I__6396\ : Span4Mux_v
    port map (
            O => \N__27750\,
            I => \N__27737\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__27747\,
            I => \N__27737\
        );

    \I__6394\ : Odrv4
    port map (
            O => \N__27742\,
            I => \N_41_0\
        );

    \I__6393\ : Odrv4
    port map (
            O => \N__27737\,
            I => \N_41_0\
        );

    \I__6392\ : InMux
    port map (
            O => \N__27732\,
            I => \N__27729\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__27729\,
            I => \this_sprites_ram.mem_out_bus4_0\
        );

    \I__6390\ : InMux
    port map (
            O => \N__27726\,
            I => \N__27723\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__27723\,
            I => \N__27720\
        );

    \I__6388\ : Sp12to4
    port map (
            O => \N__27720\,
            I => \N__27717\
        );

    \I__6387\ : Span12Mux_v
    port map (
            O => \N__27717\,
            I => \N__27714\
        );

    \I__6386\ : Odrv12
    port map (
            O => \N__27714\,
            I => \this_sprites_ram.mem_out_bus0_0\
        );

    \I__6385\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27708\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__27708\,
            I => \this_sprites_ram.mem_out_bus4_3\
        );

    \I__6383\ : InMux
    port map (
            O => \N__27705\,
            I => \N__27702\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__27702\,
            I => \N__27699\
        );

    \I__6381\ : Span4Mux_v
    port map (
            O => \N__27699\,
            I => \N__27696\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__27696\,
            I => \N__27693\
        );

    \I__6379\ : Span4Mux_v
    port map (
            O => \N__27693\,
            I => \N__27690\
        );

    \I__6378\ : Odrv4
    port map (
            O => \N__27690\,
            I => \this_sprites_ram.mem_out_bus0_3\
        );

    \I__6377\ : InMux
    port map (
            O => \N__27687\,
            I => \N__27684\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__27684\,
            I => \N__27681\
        );

    \I__6375\ : Sp12to4
    port map (
            O => \N__27681\,
            I => \N__27678\
        );

    \I__6374\ : Odrv12
    port map (
            O => \N__27678\,
            I => \this_sprites_ram.mem_out_bus6_3\
        );

    \I__6373\ : InMux
    port map (
            O => \N__27675\,
            I => \N__27672\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__27672\,
            I => \N__27669\
        );

    \I__6371\ : Span4Mux_v
    port map (
            O => \N__27669\,
            I => \N__27666\
        );

    \I__6370\ : Odrv4
    port map (
            O => \N__27666\,
            I => \this_sprites_ram.mem_out_bus2_3\
        );

    \I__6369\ : InMux
    port map (
            O => \N__27663\,
            I => \N__27660\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__27660\,
            I => \N__27654\
        );

    \I__6367\ : CascadeMux
    port map (
            O => \N__27659\,
            I => \N__27650\
        );

    \I__6366\ : CascadeMux
    port map (
            O => \N__27658\,
            I => \N__27647\
        );

    \I__6365\ : InMux
    port map (
            O => \N__27657\,
            I => \N__27642\
        );

    \I__6364\ : Span4Mux_h
    port map (
            O => \N__27654\,
            I => \N__27639\
        );

    \I__6363\ : InMux
    port map (
            O => \N__27653\,
            I => \N__27634\
        );

    \I__6362\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27634\
        );

    \I__6361\ : InMux
    port map (
            O => \N__27647\,
            I => \N__27631\
        );

    \I__6360\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27628\
        );

    \I__6359\ : InMux
    port map (
            O => \N__27645\,
            I => \N__27625\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__27642\,
            I => \this_start_data_delay.N_992\
        );

    \I__6357\ : Odrv4
    port map (
            O => \N__27639\,
            I => \this_start_data_delay.N_992\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__27634\,
            I => \this_start_data_delay.N_992\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__27631\,
            I => \this_start_data_delay.N_992\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__27628\,
            I => \this_start_data_delay.N_992\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__27625\,
            I => \this_start_data_delay.N_992\
        );

    \I__6352\ : InMux
    port map (
            O => \N__27612\,
            I => \N__27608\
        );

    \I__6351\ : InMux
    port map (
            O => \N__27611\,
            I => \N__27604\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__27608\,
            I => \N__27598\
        );

    \I__6349\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27595\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__27604\,
            I => \N__27592\
        );

    \I__6347\ : InMux
    port map (
            O => \N__27603\,
            I => \N__27589\
        );

    \I__6346\ : InMux
    port map (
            O => \N__27602\,
            I => \N__27584\
        );

    \I__6345\ : InMux
    port map (
            O => \N__27601\,
            I => \N__27584\
        );

    \I__6344\ : Odrv4
    port map (
            O => \N__27598\,
            I => \this_start_data_delay.N_110\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__27595\,
            I => \this_start_data_delay.N_110\
        );

    \I__6342\ : Odrv4
    port map (
            O => \N__27592\,
            I => \this_start_data_delay.N_110\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__27589\,
            I => \this_start_data_delay.N_110\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__27584\,
            I => \this_start_data_delay.N_110\
        );

    \I__6339\ : InMux
    port map (
            O => \N__27573\,
            I => \N__27570\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__27570\,
            I => \un1_M_this_sprites_address_q_cry_7_THRU_CO\
        );

    \I__6337\ : CascadeMux
    port map (
            O => \N__27567\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_8_cascade_\
        );

    \I__6336\ : InMux
    port map (
            O => \N__27564\,
            I => \N__27554\
        );

    \I__6335\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27547\
        );

    \I__6334\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27547\
        );

    \I__6333\ : InMux
    port map (
            O => \N__27561\,
            I => \N__27547\
        );

    \I__6332\ : InMux
    port map (
            O => \N__27560\,
            I => \N__27544\
        );

    \I__6331\ : InMux
    port map (
            O => \N__27559\,
            I => \N__27537\
        );

    \I__6330\ : InMux
    port map (
            O => \N__27558\,
            I => \N__27537\
        );

    \I__6329\ : InMux
    port map (
            O => \N__27557\,
            I => \N__27534\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__27554\,
            I => \N__27527\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__27547\,
            I => \N__27527\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__27544\,
            I => \N__27524\
        );

    \I__6325\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27519\
        );

    \I__6324\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27519\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__27537\,
            I => \N__27512\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__27534\,
            I => \N__27512\
        );

    \I__6321\ : InMux
    port map (
            O => \N__27533\,
            I => \N__27507\
        );

    \I__6320\ : InMux
    port map (
            O => \N__27532\,
            I => \N__27507\
        );

    \I__6319\ : Span4Mux_v
    port map (
            O => \N__27527\,
            I => \N__27500\
        );

    \I__6318\ : Span4Mux_h
    port map (
            O => \N__27524\,
            I => \N__27500\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__27519\,
            I => \N__27500\
        );

    \I__6316\ : InMux
    port map (
            O => \N__27518\,
            I => \N__27497\
        );

    \I__6315\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27494\
        );

    \I__6314\ : Odrv4
    port map (
            O => \N__27512\,
            I => \this_start_data_delay.N_990\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__27507\,
            I => \this_start_data_delay.N_990\
        );

    \I__6312\ : Odrv4
    port map (
            O => \N__27500\,
            I => \this_start_data_delay.N_990\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__27497\,
            I => \this_start_data_delay.N_990\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__27494\,
            I => \this_start_data_delay.N_990\
        );

    \I__6309\ : CascadeMux
    port map (
            O => \N__27483\,
            I => \N__27480\
        );

    \I__6308\ : CascadeBuf
    port map (
            O => \N__27480\,
            I => \N__27477\
        );

    \I__6307\ : CascadeMux
    port map (
            O => \N__27477\,
            I => \N__27474\
        );

    \I__6306\ : CascadeBuf
    port map (
            O => \N__27474\,
            I => \N__27471\
        );

    \I__6305\ : CascadeMux
    port map (
            O => \N__27471\,
            I => \N__27468\
        );

    \I__6304\ : CascadeBuf
    port map (
            O => \N__27468\,
            I => \N__27465\
        );

    \I__6303\ : CascadeMux
    port map (
            O => \N__27465\,
            I => \N__27462\
        );

    \I__6302\ : CascadeBuf
    port map (
            O => \N__27462\,
            I => \N__27459\
        );

    \I__6301\ : CascadeMux
    port map (
            O => \N__27459\,
            I => \N__27456\
        );

    \I__6300\ : CascadeBuf
    port map (
            O => \N__27456\,
            I => \N__27453\
        );

    \I__6299\ : CascadeMux
    port map (
            O => \N__27453\,
            I => \N__27450\
        );

    \I__6298\ : CascadeBuf
    port map (
            O => \N__27450\,
            I => \N__27447\
        );

    \I__6297\ : CascadeMux
    port map (
            O => \N__27447\,
            I => \N__27444\
        );

    \I__6296\ : CascadeBuf
    port map (
            O => \N__27444\,
            I => \N__27441\
        );

    \I__6295\ : CascadeMux
    port map (
            O => \N__27441\,
            I => \N__27438\
        );

    \I__6294\ : CascadeBuf
    port map (
            O => \N__27438\,
            I => \N__27435\
        );

    \I__6293\ : CascadeMux
    port map (
            O => \N__27435\,
            I => \N__27432\
        );

    \I__6292\ : CascadeBuf
    port map (
            O => \N__27432\,
            I => \N__27429\
        );

    \I__6291\ : CascadeMux
    port map (
            O => \N__27429\,
            I => \N__27426\
        );

    \I__6290\ : CascadeBuf
    port map (
            O => \N__27426\,
            I => \N__27423\
        );

    \I__6289\ : CascadeMux
    port map (
            O => \N__27423\,
            I => \N__27420\
        );

    \I__6288\ : CascadeBuf
    port map (
            O => \N__27420\,
            I => \N__27417\
        );

    \I__6287\ : CascadeMux
    port map (
            O => \N__27417\,
            I => \N__27414\
        );

    \I__6286\ : CascadeBuf
    port map (
            O => \N__27414\,
            I => \N__27411\
        );

    \I__6285\ : CascadeMux
    port map (
            O => \N__27411\,
            I => \N__27408\
        );

    \I__6284\ : CascadeBuf
    port map (
            O => \N__27408\,
            I => \N__27405\
        );

    \I__6283\ : CascadeMux
    port map (
            O => \N__27405\,
            I => \N__27402\
        );

    \I__6282\ : CascadeBuf
    port map (
            O => \N__27402\,
            I => \N__27399\
        );

    \I__6281\ : CascadeMux
    port map (
            O => \N__27399\,
            I => \N__27396\
        );

    \I__6280\ : CascadeBuf
    port map (
            O => \N__27396\,
            I => \N__27393\
        );

    \I__6279\ : CascadeMux
    port map (
            O => \N__27393\,
            I => \N__27390\
        );

    \I__6278\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27387\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__27387\,
            I => \N__27384\
        );

    \I__6276\ : Span4Mux_s3_v
    port map (
            O => \N__27384\,
            I => \N__27381\
        );

    \I__6275\ : Span4Mux_v
    port map (
            O => \N__27381\,
            I => \N__27375\
        );

    \I__6274\ : InMux
    port map (
            O => \N__27380\,
            I => \N__27372\
        );

    \I__6273\ : InMux
    port map (
            O => \N__27379\,
            I => \N__27369\
        );

    \I__6272\ : InMux
    port map (
            O => \N__27378\,
            I => \N__27366\
        );

    \I__6271\ : Span4Mux_v
    port map (
            O => \N__27375\,
            I => \N__27363\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__27372\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__27369\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__27366\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__6267\ : Odrv4
    port map (
            O => \N__27363\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__6266\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27351\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__27351\,
            I => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\
        );

    \I__6264\ : CEMux
    port map (
            O => \N__27348\,
            I => \N__27344\
        );

    \I__6263\ : CEMux
    port map (
            O => \N__27347\,
            I => \N__27341\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__27344\,
            I => \N__27336\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__27341\,
            I => \N__27336\
        );

    \I__6260\ : Span4Mux_v
    port map (
            O => \N__27336\,
            I => \N__27333\
        );

    \I__6259\ : Span4Mux_h
    port map (
            O => \N__27333\,
            I => \N__27330\
        );

    \I__6258\ : Odrv4
    port map (
            O => \N__27330\,
            I => \this_sprites_ram.mem_WE_10\
        );

    \I__6257\ : CEMux
    port map (
            O => \N__27327\,
            I => \N__27323\
        );

    \I__6256\ : CEMux
    port map (
            O => \N__27326\,
            I => \N__27320\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__27323\,
            I => \N__27317\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__27320\,
            I => \N__27314\
        );

    \I__6253\ : Span4Mux_h
    port map (
            O => \N__27317\,
            I => \N__27311\
        );

    \I__6252\ : Span4Mux_h
    port map (
            O => \N__27314\,
            I => \N__27308\
        );

    \I__6251\ : Odrv4
    port map (
            O => \N__27311\,
            I => \this_sprites_ram.mem_WE_8\
        );

    \I__6250\ : Odrv4
    port map (
            O => \N__27308\,
            I => \this_sprites_ram.mem_WE_8\
        );

    \I__6249\ : CEMux
    port map (
            O => \N__27303\,
            I => \N__27300\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__27300\,
            I => \N__27296\
        );

    \I__6247\ : CEMux
    port map (
            O => \N__27299\,
            I => \N__27293\
        );

    \I__6246\ : Span4Mux_v
    port map (
            O => \N__27296\,
            I => \N__27288\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__27293\,
            I => \N__27288\
        );

    \I__6244\ : Span4Mux_v
    port map (
            O => \N__27288\,
            I => \N__27285\
        );

    \I__6243\ : Odrv4
    port map (
            O => \N__27285\,
            I => \this_sprites_ram.mem_WE_12\
        );

    \I__6242\ : CEMux
    port map (
            O => \N__27282\,
            I => \N__27279\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__27279\,
            I => \N__27275\
        );

    \I__6240\ : CEMux
    port map (
            O => \N__27278\,
            I => \N__27272\
        );

    \I__6239\ : Span4Mux_s1_v
    port map (
            O => \N__27275\,
            I => \N__27267\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__27272\,
            I => \N__27267\
        );

    \I__6237\ : Span4Mux_v
    port map (
            O => \N__27267\,
            I => \N__27264\
        );

    \I__6236\ : Span4Mux_v
    port map (
            O => \N__27264\,
            I => \N__27261\
        );

    \I__6235\ : Odrv4
    port map (
            O => \N__27261\,
            I => \this_sprites_ram.mem_WE_14\
        );

    \I__6234\ : InMux
    port map (
            O => \N__27258\,
            I => \N__27255\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__27255\,
            I => \N__27251\
        );

    \I__6232\ : InMux
    port map (
            O => \N__27254\,
            I => \N__27248\
        );

    \I__6231\ : Span4Mux_v
    port map (
            O => \N__27251\,
            I => \N__27241\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__27248\,
            I => \N__27241\
        );

    \I__6229\ : InMux
    port map (
            O => \N__27247\,
            I => \N__27238\
        );

    \I__6228\ : InMux
    port map (
            O => \N__27246\,
            I => \N__27234\
        );

    \I__6227\ : Span4Mux_v
    port map (
            O => \N__27241\,
            I => \N__27228\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__27238\,
            I => \N__27228\
        );

    \I__6225\ : InMux
    port map (
            O => \N__27237\,
            I => \N__27225\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__27234\,
            I => \N__27222\
        );

    \I__6223\ : InMux
    port map (
            O => \N__27233\,
            I => \N__27219\
        );

    \I__6222\ : Span4Mux_v
    port map (
            O => \N__27228\,
            I => \N__27213\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__27225\,
            I => \N__27213\
        );

    \I__6220\ : Span4Mux_v
    port map (
            O => \N__27222\,
            I => \N__27208\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__27219\,
            I => \N__27208\
        );

    \I__6218\ : InMux
    port map (
            O => \N__27218\,
            I => \N__27205\
        );

    \I__6217\ : Span4Mux_v
    port map (
            O => \N__27213\,
            I => \N__27201\
        );

    \I__6216\ : Span4Mux_v
    port map (
            O => \N__27208\,
            I => \N__27196\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__27205\,
            I => \N__27196\
        );

    \I__6214\ : InMux
    port map (
            O => \N__27204\,
            I => \N__27193\
        );

    \I__6213\ : Odrv4
    port map (
            O => \N__27201\,
            I => \N_811_0\
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__27196\,
            I => \N_811_0\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__27193\,
            I => \N_811_0\
        );

    \I__6210\ : InMux
    port map (
            O => \N__27186\,
            I => \N__27183\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__27183\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_5\
        );

    \I__6208\ : InMux
    port map (
            O => \N__27180\,
            I => \N__27177\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__27177\,
            I => \un1_M_this_sprites_address_q_cry_4_THRU_CO\
        );

    \I__6206\ : CascadeMux
    port map (
            O => \N__27174\,
            I => \N__27171\
        );

    \I__6205\ : CascadeBuf
    port map (
            O => \N__27171\,
            I => \N__27168\
        );

    \I__6204\ : CascadeMux
    port map (
            O => \N__27168\,
            I => \N__27165\
        );

    \I__6203\ : CascadeBuf
    port map (
            O => \N__27165\,
            I => \N__27162\
        );

    \I__6202\ : CascadeMux
    port map (
            O => \N__27162\,
            I => \N__27159\
        );

    \I__6201\ : CascadeBuf
    port map (
            O => \N__27159\,
            I => \N__27156\
        );

    \I__6200\ : CascadeMux
    port map (
            O => \N__27156\,
            I => \N__27153\
        );

    \I__6199\ : CascadeBuf
    port map (
            O => \N__27153\,
            I => \N__27150\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__27150\,
            I => \N__27147\
        );

    \I__6197\ : CascadeBuf
    port map (
            O => \N__27147\,
            I => \N__27144\
        );

    \I__6196\ : CascadeMux
    port map (
            O => \N__27144\,
            I => \N__27141\
        );

    \I__6195\ : CascadeBuf
    port map (
            O => \N__27141\,
            I => \N__27138\
        );

    \I__6194\ : CascadeMux
    port map (
            O => \N__27138\,
            I => \N__27135\
        );

    \I__6193\ : CascadeBuf
    port map (
            O => \N__27135\,
            I => \N__27132\
        );

    \I__6192\ : CascadeMux
    port map (
            O => \N__27132\,
            I => \N__27129\
        );

    \I__6191\ : CascadeBuf
    port map (
            O => \N__27129\,
            I => \N__27126\
        );

    \I__6190\ : CascadeMux
    port map (
            O => \N__27126\,
            I => \N__27123\
        );

    \I__6189\ : CascadeBuf
    port map (
            O => \N__27123\,
            I => \N__27120\
        );

    \I__6188\ : CascadeMux
    port map (
            O => \N__27120\,
            I => \N__27117\
        );

    \I__6187\ : CascadeBuf
    port map (
            O => \N__27117\,
            I => \N__27114\
        );

    \I__6186\ : CascadeMux
    port map (
            O => \N__27114\,
            I => \N__27111\
        );

    \I__6185\ : CascadeBuf
    port map (
            O => \N__27111\,
            I => \N__27108\
        );

    \I__6184\ : CascadeMux
    port map (
            O => \N__27108\,
            I => \N__27105\
        );

    \I__6183\ : CascadeBuf
    port map (
            O => \N__27105\,
            I => \N__27102\
        );

    \I__6182\ : CascadeMux
    port map (
            O => \N__27102\,
            I => \N__27099\
        );

    \I__6181\ : CascadeBuf
    port map (
            O => \N__27099\,
            I => \N__27096\
        );

    \I__6180\ : CascadeMux
    port map (
            O => \N__27096\,
            I => \N__27093\
        );

    \I__6179\ : CascadeBuf
    port map (
            O => \N__27093\,
            I => \N__27090\
        );

    \I__6178\ : CascadeMux
    port map (
            O => \N__27090\,
            I => \N__27087\
        );

    \I__6177\ : CascadeBuf
    port map (
            O => \N__27087\,
            I => \N__27084\
        );

    \I__6176\ : CascadeMux
    port map (
            O => \N__27084\,
            I => \N__27081\
        );

    \I__6175\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27078\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__27078\,
            I => \N__27075\
        );

    \I__6173\ : Span4Mux_h
    port map (
            O => \N__27075\,
            I => \N__27071\
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__27074\,
            I => \N__27066\
        );

    \I__6171\ : Sp12to4
    port map (
            O => \N__27071\,
            I => \N__27063\
        );

    \I__6170\ : InMux
    port map (
            O => \N__27070\,
            I => \N__27060\
        );

    \I__6169\ : InMux
    port map (
            O => \N__27069\,
            I => \N__27057\
        );

    \I__6168\ : InMux
    port map (
            O => \N__27066\,
            I => \N__27054\
        );

    \I__6167\ : Span12Mux_s6_v
    port map (
            O => \N__27063\,
            I => \N__27051\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__27060\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__27057\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__27054\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__6163\ : Odrv12
    port map (
            O => \N__27051\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__6162\ : CEMux
    port map (
            O => \N__27042\,
            I => \N__27039\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__27039\,
            I => \N__27036\
        );

    \I__6160\ : Span4Mux_v
    port map (
            O => \N__27036\,
            I => \N__27032\
        );

    \I__6159\ : CEMux
    port map (
            O => \N__27035\,
            I => \N__27029\
        );

    \I__6158\ : Span4Mux_v
    port map (
            O => \N__27032\,
            I => \N__27024\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__27029\,
            I => \N__27024\
        );

    \I__6156\ : Span4Mux_h
    port map (
            O => \N__27024\,
            I => \N__27021\
        );

    \I__6155\ : Odrv4
    port map (
            O => \N__27021\,
            I => \this_sprites_ram.mem_WE_6\
        );

    \I__6154\ : InMux
    port map (
            O => \N__27018\,
            I => \N__27015\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__27015\,
            I => \N__27012\
        );

    \I__6152\ : Span4Mux_v
    port map (
            O => \N__27012\,
            I => \N__27009\
        );

    \I__6151\ : Odrv4
    port map (
            O => \N__27009\,
            I => \this_sprites_ram.mem_out_bus5_0\
        );

    \I__6150\ : InMux
    port map (
            O => \N__27006\,
            I => \N__27003\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__27003\,
            I => \N__27000\
        );

    \I__6148\ : Span4Mux_v
    port map (
            O => \N__27000\,
            I => \N__26997\
        );

    \I__6147\ : Span4Mux_v
    port map (
            O => \N__26997\,
            I => \N__26994\
        );

    \I__6146\ : Odrv4
    port map (
            O => \N__26994\,
            I => \this_sprites_ram.mem_out_bus1_0\
        );

    \I__6145\ : InMux
    port map (
            O => \N__26991\,
            I => \N__26988\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__26988\,
            I => \N__26985\
        );

    \I__6143\ : Span12Mux_h
    port map (
            O => \N__26985\,
            I => \N__26982\
        );

    \I__6142\ : Odrv12
    port map (
            O => \N__26982\,
            I => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\
        );

    \I__6141\ : CascadeMux
    port map (
            O => \N__26979\,
            I => \N__26976\
        );

    \I__6140\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26968\
        );

    \I__6139\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26964\
        );

    \I__6138\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26958\
        );

    \I__6137\ : InMux
    port map (
            O => \N__26973\,
            I => \N__26958\
        );

    \I__6136\ : InMux
    port map (
            O => \N__26972\,
            I => \N__26955\
        );

    \I__6135\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26952\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__26968\,
            I => \N__26949\
        );

    \I__6133\ : InMux
    port map (
            O => \N__26967\,
            I => \N__26946\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__26964\,
            I => \N__26943\
        );

    \I__6131\ : InMux
    port map (
            O => \N__26963\,
            I => \N__26940\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__26958\,
            I => \N__26937\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__26955\,
            I => \N__26934\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__26952\,
            I => \N__26931\
        );

    \I__6127\ : Span4Mux_v
    port map (
            O => \N__26949\,
            I => \N__26928\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__26946\,
            I => \N__26925\
        );

    \I__6125\ : Span4Mux_h
    port map (
            O => \N__26943\,
            I => \N__26922\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__26940\,
            I => \N__26917\
        );

    \I__6123\ : Span4Mux_v
    port map (
            O => \N__26937\,
            I => \N__26917\
        );

    \I__6122\ : Span4Mux_h
    port map (
            O => \N__26934\,
            I => \N__26912\
        );

    \I__6121\ : Span4Mux_h
    port map (
            O => \N__26931\,
            I => \N__26912\
        );

    \I__6120\ : Span4Mux_h
    port map (
            O => \N__26928\,
            I => \N__26907\
        );

    \I__6119\ : Span4Mux_h
    port map (
            O => \N__26925\,
            I => \N__26907\
        );

    \I__6118\ : Odrv4
    port map (
            O => \N__26922\,
            I => \N_10_0\
        );

    \I__6117\ : Odrv4
    port map (
            O => \N__26917\,
            I => \N_10_0\
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__26912\,
            I => \N_10_0\
        );

    \I__6115\ : Odrv4
    port map (
            O => \N__26907\,
            I => \N_10_0\
        );

    \I__6114\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26895\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__26895\,
            I => \this_start_data_delay.M_this_state_d62Z0Z_11\
        );

    \I__6112\ : InMux
    port map (
            O => \N__26892\,
            I => \N__26889\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__26889\,
            I => \this_start_data_delay.M_this_state_d62Z0Z_10\
        );

    \I__6110\ : CascadeMux
    port map (
            O => \N__26886\,
            I => \this_start_data_delay.M_this_state_d62Z0Z_9_cascade_\
        );

    \I__6109\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26880\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__26880\,
            I => \this_start_data_delay.M_this_state_d62Z0Z_8\
        );

    \I__6107\ : InMux
    port map (
            O => \N__26877\,
            I => \N__26872\
        );

    \I__6106\ : InMux
    port map (
            O => \N__26876\,
            I => \N__26868\
        );

    \I__6105\ : InMux
    port map (
            O => \N__26875\,
            I => \N__26864\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__26872\,
            I => \N__26861\
        );

    \I__6103\ : InMux
    port map (
            O => \N__26871\,
            I => \N__26858\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__26868\,
            I => \N__26855\
        );

    \I__6101\ : InMux
    port map (
            O => \N__26867\,
            I => \N__26852\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__26864\,
            I => \N__26848\
        );

    \I__6099\ : Span4Mux_h
    port map (
            O => \N__26861\,
            I => \N__26845\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__26858\,
            I => \N__26840\
        );

    \I__6097\ : Span4Mux_h
    port map (
            O => \N__26855\,
            I => \N__26840\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__26852\,
            I => \N__26837\
        );

    \I__6095\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26834\
        );

    \I__6094\ : Span4Mux_v
    port map (
            O => \N__26848\,
            I => \N__26831\
        );

    \I__6093\ : Span4Mux_v
    port map (
            O => \N__26845\,
            I => \N__26828\
        );

    \I__6092\ : Span4Mux_v
    port map (
            O => \N__26840\,
            I => \N__26825\
        );

    \I__6091\ : Span4Mux_h
    port map (
            O => \N__26837\,
            I => \N__26820\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__26834\,
            I => \N__26820\
        );

    \I__6089\ : Odrv4
    port map (
            O => \N__26831\,
            I => \this_start_data_delay.M_this_state_dZ0Z62\
        );

    \I__6088\ : Odrv4
    port map (
            O => \N__26828\,
            I => \this_start_data_delay.M_this_state_dZ0Z62\
        );

    \I__6087\ : Odrv4
    port map (
            O => \N__26825\,
            I => \this_start_data_delay.M_this_state_dZ0Z62\
        );

    \I__6086\ : Odrv4
    port map (
            O => \N__26820\,
            I => \this_start_data_delay.M_this_state_dZ0Z62\
        );

    \I__6085\ : CascadeMux
    port map (
            O => \N__26811\,
            I => \N__26808\
        );

    \I__6084\ : InMux
    port map (
            O => \N__26808\,
            I => \N__26805\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__26805\,
            I => \M_this_data_count_q_3_10\
        );

    \I__6082\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26799\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__26799\,
            I => \N__26796\
        );

    \I__6080\ : Odrv12
    port map (
            O => \N__26796\,
            I => \this_start_data_delay_M_this_external_address_q_3_i_0_15\
        );

    \I__6079\ : InMux
    port map (
            O => \N__26793\,
            I => \N__26781\
        );

    \I__6078\ : InMux
    port map (
            O => \N__26792\,
            I => \N__26781\
        );

    \I__6077\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26772\
        );

    \I__6076\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26772\
        );

    \I__6075\ : InMux
    port map (
            O => \N__26789\,
            I => \N__26772\
        );

    \I__6074\ : InMux
    port map (
            O => \N__26788\,
            I => \N__26772\
        );

    \I__6073\ : InMux
    port map (
            O => \N__26787\,
            I => \N__26769\
        );

    \I__6072\ : CascadeMux
    port map (
            O => \N__26786\,
            I => \N__26766\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__26781\,
            I => \N__26762\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__26772\,
            I => \N__26759\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__26769\,
            I => \N__26756\
        );

    \I__6068\ : InMux
    port map (
            O => \N__26766\,
            I => \N__26752\
        );

    \I__6067\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26749\
        );

    \I__6066\ : Span4Mux_v
    port map (
            O => \N__26762\,
            I => \N__26746\
        );

    \I__6065\ : Span4Mux_v
    port map (
            O => \N__26759\,
            I => \N__26743\
        );

    \I__6064\ : Span4Mux_h
    port map (
            O => \N__26756\,
            I => \N__26740\
        );

    \I__6063\ : InMux
    port map (
            O => \N__26755\,
            I => \N__26737\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__26752\,
            I => \N__26734\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__26749\,
            I => \N__26731\
        );

    \I__6060\ : Span4Mux_h
    port map (
            O => \N__26746\,
            I => \N__26726\
        );

    \I__6059\ : Span4Mux_h
    port map (
            O => \N__26743\,
            I => \N__26726\
        );

    \I__6058\ : Sp12to4
    port map (
            O => \N__26740\,
            I => \N__26721\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__26737\,
            I => \N__26721\
        );

    \I__6056\ : Span4Mux_v
    port map (
            O => \N__26734\,
            I => \N__26716\
        );

    \I__6055\ : Span4Mux_v
    port map (
            O => \N__26731\,
            I => \N__26716\
        );

    \I__6054\ : Sp12to4
    port map (
            O => \N__26726\,
            I => \N__26713\
        );

    \I__6053\ : Span12Mux_s10_v
    port map (
            O => \N__26721\,
            I => \N__26710\
        );

    \I__6052\ : Odrv4
    port map (
            O => \N__26716\,
            I => \N_116\
        );

    \I__6051\ : Odrv12
    port map (
            O => \N__26713\,
            I => \N_116\
        );

    \I__6050\ : Odrv12
    port map (
            O => \N__26710\,
            I => \N_116\
        );

    \I__6049\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26700\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__26700\,
            I => \M_this_external_address_q_3_0_13\
        );

    \I__6047\ : InMux
    port map (
            O => \N__26697\,
            I => \N__26694\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__26694\,
            I => \N__26691\
        );

    \I__6045\ : Span4Mux_s2_v
    port map (
            O => \N__26691\,
            I => \N__26688\
        );

    \I__6044\ : Span4Mux_h
    port map (
            O => \N__26688\,
            I => \N__26685\
        );

    \I__6043\ : Span4Mux_v
    port map (
            O => \N__26685\,
            I => \N__26682\
        );

    \I__6042\ : Sp12to4
    port map (
            O => \N__26682\,
            I => \N__26679\
        );

    \I__6041\ : Odrv12
    port map (
            O => \N__26679\,
            I => \M_this_map_ram_read_data_0\
        );

    \I__6040\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26673\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__26673\,
            I => \N__26670\
        );

    \I__6038\ : Span12Mux_h
    port map (
            O => \N__26670\,
            I => \N__26667\
        );

    \I__6037\ : Span12Mux_v
    port map (
            O => \N__26667\,
            I => \N__26664\
        );

    \I__6036\ : Odrv12
    port map (
            O => \N__26664\,
            I => \this_ppu.un3_sprites_addr_cry_5_c_RNI55GZ0Z8\
        );

    \I__6035\ : CascadeMux
    port map (
            O => \N__26661\,
            I => \N__26658\
        );

    \I__6034\ : CascadeBuf
    port map (
            O => \N__26658\,
            I => \N__26655\
        );

    \I__6033\ : CascadeMux
    port map (
            O => \N__26655\,
            I => \N__26652\
        );

    \I__6032\ : CascadeBuf
    port map (
            O => \N__26652\,
            I => \N__26649\
        );

    \I__6031\ : CascadeMux
    port map (
            O => \N__26649\,
            I => \N__26646\
        );

    \I__6030\ : CascadeBuf
    port map (
            O => \N__26646\,
            I => \N__26643\
        );

    \I__6029\ : CascadeMux
    port map (
            O => \N__26643\,
            I => \N__26640\
        );

    \I__6028\ : CascadeBuf
    port map (
            O => \N__26640\,
            I => \N__26637\
        );

    \I__6027\ : CascadeMux
    port map (
            O => \N__26637\,
            I => \N__26634\
        );

    \I__6026\ : CascadeBuf
    port map (
            O => \N__26634\,
            I => \N__26631\
        );

    \I__6025\ : CascadeMux
    port map (
            O => \N__26631\,
            I => \N__26628\
        );

    \I__6024\ : CascadeBuf
    port map (
            O => \N__26628\,
            I => \N__26625\
        );

    \I__6023\ : CascadeMux
    port map (
            O => \N__26625\,
            I => \N__26622\
        );

    \I__6022\ : CascadeBuf
    port map (
            O => \N__26622\,
            I => \N__26619\
        );

    \I__6021\ : CascadeMux
    port map (
            O => \N__26619\,
            I => \N__26616\
        );

    \I__6020\ : CascadeBuf
    port map (
            O => \N__26616\,
            I => \N__26613\
        );

    \I__6019\ : CascadeMux
    port map (
            O => \N__26613\,
            I => \N__26610\
        );

    \I__6018\ : CascadeBuf
    port map (
            O => \N__26610\,
            I => \N__26607\
        );

    \I__6017\ : CascadeMux
    port map (
            O => \N__26607\,
            I => \N__26604\
        );

    \I__6016\ : CascadeBuf
    port map (
            O => \N__26604\,
            I => \N__26601\
        );

    \I__6015\ : CascadeMux
    port map (
            O => \N__26601\,
            I => \N__26598\
        );

    \I__6014\ : CascadeBuf
    port map (
            O => \N__26598\,
            I => \N__26595\
        );

    \I__6013\ : CascadeMux
    port map (
            O => \N__26595\,
            I => \N__26592\
        );

    \I__6012\ : CascadeBuf
    port map (
            O => \N__26592\,
            I => \N__26589\
        );

    \I__6011\ : CascadeMux
    port map (
            O => \N__26589\,
            I => \N__26586\
        );

    \I__6010\ : CascadeBuf
    port map (
            O => \N__26586\,
            I => \N__26583\
        );

    \I__6009\ : CascadeMux
    port map (
            O => \N__26583\,
            I => \N__26580\
        );

    \I__6008\ : CascadeBuf
    port map (
            O => \N__26580\,
            I => \N__26577\
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__26577\,
            I => \N__26574\
        );

    \I__6006\ : CascadeBuf
    port map (
            O => \N__26574\,
            I => \N__26571\
        );

    \I__6005\ : CascadeMux
    port map (
            O => \N__26571\,
            I => \N__26568\
        );

    \I__6004\ : InMux
    port map (
            O => \N__26568\,
            I => \N__26565\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__26565\,
            I => \N__26562\
        );

    \I__6002\ : Odrv4
    port map (
            O => \N__26562\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__6001\ : CascadeMux
    port map (
            O => \N__26559\,
            I => \N__26556\
        );

    \I__6000\ : CascadeBuf
    port map (
            O => \N__26556\,
            I => \N__26553\
        );

    \I__5999\ : CascadeMux
    port map (
            O => \N__26553\,
            I => \N__26550\
        );

    \I__5998\ : CascadeBuf
    port map (
            O => \N__26550\,
            I => \N__26547\
        );

    \I__5997\ : CascadeMux
    port map (
            O => \N__26547\,
            I => \N__26544\
        );

    \I__5996\ : CascadeBuf
    port map (
            O => \N__26544\,
            I => \N__26541\
        );

    \I__5995\ : CascadeMux
    port map (
            O => \N__26541\,
            I => \N__26538\
        );

    \I__5994\ : CascadeBuf
    port map (
            O => \N__26538\,
            I => \N__26535\
        );

    \I__5993\ : CascadeMux
    port map (
            O => \N__26535\,
            I => \N__26532\
        );

    \I__5992\ : CascadeBuf
    port map (
            O => \N__26532\,
            I => \N__26529\
        );

    \I__5991\ : CascadeMux
    port map (
            O => \N__26529\,
            I => \N__26526\
        );

    \I__5990\ : CascadeBuf
    port map (
            O => \N__26526\,
            I => \N__26523\
        );

    \I__5989\ : CascadeMux
    port map (
            O => \N__26523\,
            I => \N__26520\
        );

    \I__5988\ : CascadeBuf
    port map (
            O => \N__26520\,
            I => \N__26517\
        );

    \I__5987\ : CascadeMux
    port map (
            O => \N__26517\,
            I => \N__26514\
        );

    \I__5986\ : CascadeBuf
    port map (
            O => \N__26514\,
            I => \N__26511\
        );

    \I__5985\ : CascadeMux
    port map (
            O => \N__26511\,
            I => \N__26508\
        );

    \I__5984\ : CascadeBuf
    port map (
            O => \N__26508\,
            I => \N__26505\
        );

    \I__5983\ : CascadeMux
    port map (
            O => \N__26505\,
            I => \N__26502\
        );

    \I__5982\ : CascadeBuf
    port map (
            O => \N__26502\,
            I => \N__26499\
        );

    \I__5981\ : CascadeMux
    port map (
            O => \N__26499\,
            I => \N__26496\
        );

    \I__5980\ : CascadeBuf
    port map (
            O => \N__26496\,
            I => \N__26493\
        );

    \I__5979\ : CascadeMux
    port map (
            O => \N__26493\,
            I => \N__26490\
        );

    \I__5978\ : CascadeBuf
    port map (
            O => \N__26490\,
            I => \N__26487\
        );

    \I__5977\ : CascadeMux
    port map (
            O => \N__26487\,
            I => \N__26484\
        );

    \I__5976\ : CascadeBuf
    port map (
            O => \N__26484\,
            I => \N__26481\
        );

    \I__5975\ : CascadeMux
    port map (
            O => \N__26481\,
            I => \N__26478\
        );

    \I__5974\ : CascadeBuf
    port map (
            O => \N__26478\,
            I => \N__26475\
        );

    \I__5973\ : CascadeMux
    port map (
            O => \N__26475\,
            I => \N__26472\
        );

    \I__5972\ : CascadeBuf
    port map (
            O => \N__26472\,
            I => \N__26469\
        );

    \I__5971\ : CascadeMux
    port map (
            O => \N__26469\,
            I => \N__26466\
        );

    \I__5970\ : InMux
    port map (
            O => \N__26466\,
            I => \N__26463\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__26463\,
            I => \N__26460\
        );

    \I__5968\ : Span4Mux_h
    port map (
            O => \N__26460\,
            I => \N__26454\
        );

    \I__5967\ : CascadeMux
    port map (
            O => \N__26459\,
            I => \N__26451\
        );

    \I__5966\ : CascadeMux
    port map (
            O => \N__26458\,
            I => \N__26448\
        );

    \I__5965\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26445\
        );

    \I__5964\ : Sp12to4
    port map (
            O => \N__26454\,
            I => \N__26442\
        );

    \I__5963\ : InMux
    port map (
            O => \N__26451\,
            I => \N__26439\
        );

    \I__5962\ : InMux
    port map (
            O => \N__26448\,
            I => \N__26436\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__26445\,
            I => \N__26431\
        );

    \I__5960\ : Span12Mux_s8_v
    port map (
            O => \N__26442\,
            I => \N__26431\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__26439\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__26436\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5957\ : Odrv12
    port map (
            O => \N__26431\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5956\ : InMux
    port map (
            O => \N__26424\,
            I => \N__26421\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__26421\,
            I => \N__26418\
        );

    \I__5954\ : Odrv4
    port map (
            O => \N__26418\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_9\
        );

    \I__5953\ : InMux
    port map (
            O => \N__26415\,
            I => \N__26412\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__26412\,
            I => \un1_M_this_sprites_address_q_cry_8_THRU_CO\
        );

    \I__5951\ : CascadeMux
    port map (
            O => \N__26409\,
            I => \N__26406\
        );

    \I__5950\ : CascadeBuf
    port map (
            O => \N__26406\,
            I => \N__26403\
        );

    \I__5949\ : CascadeMux
    port map (
            O => \N__26403\,
            I => \N__26400\
        );

    \I__5948\ : CascadeBuf
    port map (
            O => \N__26400\,
            I => \N__26397\
        );

    \I__5947\ : CascadeMux
    port map (
            O => \N__26397\,
            I => \N__26394\
        );

    \I__5946\ : CascadeBuf
    port map (
            O => \N__26394\,
            I => \N__26391\
        );

    \I__5945\ : CascadeMux
    port map (
            O => \N__26391\,
            I => \N__26388\
        );

    \I__5944\ : CascadeBuf
    port map (
            O => \N__26388\,
            I => \N__26385\
        );

    \I__5943\ : CascadeMux
    port map (
            O => \N__26385\,
            I => \N__26382\
        );

    \I__5942\ : CascadeBuf
    port map (
            O => \N__26382\,
            I => \N__26379\
        );

    \I__5941\ : CascadeMux
    port map (
            O => \N__26379\,
            I => \N__26376\
        );

    \I__5940\ : CascadeBuf
    port map (
            O => \N__26376\,
            I => \N__26373\
        );

    \I__5939\ : CascadeMux
    port map (
            O => \N__26373\,
            I => \N__26370\
        );

    \I__5938\ : CascadeBuf
    port map (
            O => \N__26370\,
            I => \N__26367\
        );

    \I__5937\ : CascadeMux
    port map (
            O => \N__26367\,
            I => \N__26364\
        );

    \I__5936\ : CascadeBuf
    port map (
            O => \N__26364\,
            I => \N__26361\
        );

    \I__5935\ : CascadeMux
    port map (
            O => \N__26361\,
            I => \N__26358\
        );

    \I__5934\ : CascadeBuf
    port map (
            O => \N__26358\,
            I => \N__26355\
        );

    \I__5933\ : CascadeMux
    port map (
            O => \N__26355\,
            I => \N__26352\
        );

    \I__5932\ : CascadeBuf
    port map (
            O => \N__26352\,
            I => \N__26349\
        );

    \I__5931\ : CascadeMux
    port map (
            O => \N__26349\,
            I => \N__26346\
        );

    \I__5930\ : CascadeBuf
    port map (
            O => \N__26346\,
            I => \N__26343\
        );

    \I__5929\ : CascadeMux
    port map (
            O => \N__26343\,
            I => \N__26340\
        );

    \I__5928\ : CascadeBuf
    port map (
            O => \N__26340\,
            I => \N__26337\
        );

    \I__5927\ : CascadeMux
    port map (
            O => \N__26337\,
            I => \N__26334\
        );

    \I__5926\ : CascadeBuf
    port map (
            O => \N__26334\,
            I => \N__26331\
        );

    \I__5925\ : CascadeMux
    port map (
            O => \N__26331\,
            I => \N__26328\
        );

    \I__5924\ : CascadeBuf
    port map (
            O => \N__26328\,
            I => \N__26325\
        );

    \I__5923\ : CascadeMux
    port map (
            O => \N__26325\,
            I => \N__26322\
        );

    \I__5922\ : CascadeBuf
    port map (
            O => \N__26322\,
            I => \N__26319\
        );

    \I__5921\ : CascadeMux
    port map (
            O => \N__26319\,
            I => \N__26316\
        );

    \I__5920\ : InMux
    port map (
            O => \N__26316\,
            I => \N__26313\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__26313\,
            I => \N__26310\
        );

    \I__5918\ : Span4Mux_h
    port map (
            O => \N__26310\,
            I => \N__26305\
        );

    \I__5917\ : CascadeMux
    port map (
            O => \N__26309\,
            I => \N__26302\
        );

    \I__5916\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26298\
        );

    \I__5915\ : Sp12to4
    port map (
            O => \N__26305\,
            I => \N__26295\
        );

    \I__5914\ : InMux
    port map (
            O => \N__26302\,
            I => \N__26292\
        );

    \I__5913\ : InMux
    port map (
            O => \N__26301\,
            I => \N__26289\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__26298\,
            I => \N__26286\
        );

    \I__5911\ : Span12Mux_s7_v
    port map (
            O => \N__26295\,
            I => \N__26283\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__26292\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__26289\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__5908\ : Odrv4
    port map (
            O => \N__26286\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__5907\ : Odrv12
    port map (
            O => \N__26283\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__5906\ : InMux
    port map (
            O => \N__26274\,
            I => \N__26267\
        );

    \I__5905\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26264\
        );

    \I__5904\ : InMux
    port map (
            O => \N__26272\,
            I => \N__26259\
        );

    \I__5903\ : InMux
    port map (
            O => \N__26271\,
            I => \N__26259\
        );

    \I__5902\ : InMux
    port map (
            O => \N__26270\,
            I => \N__26256\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__26267\,
            I => \N__26252\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__26264\,
            I => \N__26245\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__26259\,
            I => \N__26245\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__26256\,
            I => \N__26245\
        );

    \I__5897\ : InMux
    port map (
            O => \N__26255\,
            I => \N__26242\
        );

    \I__5896\ : Span4Mux_h
    port map (
            O => \N__26252\,
            I => \N__26239\
        );

    \I__5895\ : Span4Mux_v
    port map (
            O => \N__26245\,
            I => \N__26236\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__26242\,
            I => \N__26233\
        );

    \I__5893\ : Odrv4
    port map (
            O => \N__26239\,
            I => \this_start_data_delay.N_86_0\
        );

    \I__5892\ : Odrv4
    port map (
            O => \N__26236\,
            I => \this_start_data_delay.N_86_0\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__26233\,
            I => \this_start_data_delay.N_86_0\
        );

    \I__5890\ : CascadeMux
    port map (
            O => \N__26226\,
            I => \N__26219\
        );

    \I__5889\ : CascadeMux
    port map (
            O => \N__26225\,
            I => \N__26215\
        );

    \I__5888\ : InMux
    port map (
            O => \N__26224\,
            I => \N__26175\
        );

    \I__5887\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26175\
        );

    \I__5886\ : InMux
    port map (
            O => \N__26222\,
            I => \N__26172\
        );

    \I__5885\ : InMux
    port map (
            O => \N__26219\,
            I => \N__26169\
        );

    \I__5884\ : InMux
    port map (
            O => \N__26218\,
            I => \N__26166\
        );

    \I__5883\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26161\
        );

    \I__5882\ : InMux
    port map (
            O => \N__26214\,
            I => \N__26161\
        );

    \I__5881\ : InMux
    port map (
            O => \N__26213\,
            I => \N__26156\
        );

    \I__5880\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26156\
        );

    \I__5879\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26153\
        );

    \I__5878\ : InMux
    port map (
            O => \N__26210\,
            I => \N__26148\
        );

    \I__5877\ : InMux
    port map (
            O => \N__26209\,
            I => \N__26148\
        );

    \I__5876\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26143\
        );

    \I__5875\ : InMux
    port map (
            O => \N__26207\,
            I => \N__26143\
        );

    \I__5874\ : InMux
    port map (
            O => \N__26206\,
            I => \N__26140\
        );

    \I__5873\ : InMux
    port map (
            O => \N__26205\,
            I => \N__26137\
        );

    \I__5872\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26134\
        );

    \I__5871\ : InMux
    port map (
            O => \N__26203\,
            I => \N__26131\
        );

    \I__5870\ : InMux
    port map (
            O => \N__26202\,
            I => \N__26126\
        );

    \I__5869\ : InMux
    port map (
            O => \N__26201\,
            I => \N__26126\
        );

    \I__5868\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26123\
        );

    \I__5867\ : InMux
    port map (
            O => \N__26199\,
            I => \N__26120\
        );

    \I__5866\ : InMux
    port map (
            O => \N__26198\,
            I => \N__26115\
        );

    \I__5865\ : InMux
    port map (
            O => \N__26197\,
            I => \N__26115\
        );

    \I__5864\ : InMux
    port map (
            O => \N__26196\,
            I => \N__26112\
        );

    \I__5863\ : InMux
    port map (
            O => \N__26195\,
            I => \N__26107\
        );

    \I__5862\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26107\
        );

    \I__5861\ : InMux
    port map (
            O => \N__26193\,
            I => \N__26102\
        );

    \I__5860\ : InMux
    port map (
            O => \N__26192\,
            I => \N__26102\
        );

    \I__5859\ : InMux
    port map (
            O => \N__26191\,
            I => \N__26097\
        );

    \I__5858\ : InMux
    port map (
            O => \N__26190\,
            I => \N__26097\
        );

    \I__5857\ : InMux
    port map (
            O => \N__26189\,
            I => \N__26090\
        );

    \I__5856\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26090\
        );

    \I__5855\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26090\
        );

    \I__5854\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26085\
        );

    \I__5853\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26085\
        );

    \I__5852\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26082\
        );

    \I__5851\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26077\
        );

    \I__5850\ : InMux
    port map (
            O => \N__26182\,
            I => \N__26077\
        );

    \I__5849\ : InMux
    port map (
            O => \N__26181\,
            I => \N__26072\
        );

    \I__5848\ : InMux
    port map (
            O => \N__26180\,
            I => \N__26072\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__26175\,
            I => \N__26041\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__26172\,
            I => \N__26038\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__26169\,
            I => \N__26035\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__26166\,
            I => \N__26032\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__26161\,
            I => \N__26029\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__26156\,
            I => \N__26026\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__26153\,
            I => \N__26023\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__26148\,
            I => \N__26020\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__26143\,
            I => \N__26017\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__26140\,
            I => \N__26014\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__26137\,
            I => \N__26011\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__26134\,
            I => \N__26008\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__26131\,
            I => \N__26005\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__26126\,
            I => \N__26002\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__26123\,
            I => \N__25999\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__26120\,
            I => \N__25996\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__26115\,
            I => \N__25993\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__26112\,
            I => \N__25990\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__26107\,
            I => \N__25987\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__26102\,
            I => \N__25984\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__26097\,
            I => \N__25981\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__26090\,
            I => \N__25978\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__26085\,
            I => \N__25975\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__26082\,
            I => \N__25972\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__26077\,
            I => \N__25969\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__26072\,
            I => \N__25966\
        );

    \I__5821\ : SRMux
    port map (
            O => \N__26071\,
            I => \N__25857\
        );

    \I__5820\ : SRMux
    port map (
            O => \N__26070\,
            I => \N__25857\
        );

    \I__5819\ : SRMux
    port map (
            O => \N__26069\,
            I => \N__25857\
        );

    \I__5818\ : SRMux
    port map (
            O => \N__26068\,
            I => \N__25857\
        );

    \I__5817\ : SRMux
    port map (
            O => \N__26067\,
            I => \N__25857\
        );

    \I__5816\ : SRMux
    port map (
            O => \N__26066\,
            I => \N__25857\
        );

    \I__5815\ : SRMux
    port map (
            O => \N__26065\,
            I => \N__25857\
        );

    \I__5814\ : SRMux
    port map (
            O => \N__26064\,
            I => \N__25857\
        );

    \I__5813\ : SRMux
    port map (
            O => \N__26063\,
            I => \N__25857\
        );

    \I__5812\ : SRMux
    port map (
            O => \N__26062\,
            I => \N__25857\
        );

    \I__5811\ : SRMux
    port map (
            O => \N__26061\,
            I => \N__25857\
        );

    \I__5810\ : SRMux
    port map (
            O => \N__26060\,
            I => \N__25857\
        );

    \I__5809\ : SRMux
    port map (
            O => \N__26059\,
            I => \N__25857\
        );

    \I__5808\ : SRMux
    port map (
            O => \N__26058\,
            I => \N__25857\
        );

    \I__5807\ : SRMux
    port map (
            O => \N__26057\,
            I => \N__25857\
        );

    \I__5806\ : SRMux
    port map (
            O => \N__26056\,
            I => \N__25857\
        );

    \I__5805\ : SRMux
    port map (
            O => \N__26055\,
            I => \N__25857\
        );

    \I__5804\ : SRMux
    port map (
            O => \N__26054\,
            I => \N__25857\
        );

    \I__5803\ : SRMux
    port map (
            O => \N__26053\,
            I => \N__25857\
        );

    \I__5802\ : SRMux
    port map (
            O => \N__26052\,
            I => \N__25857\
        );

    \I__5801\ : SRMux
    port map (
            O => \N__26051\,
            I => \N__25857\
        );

    \I__5800\ : SRMux
    port map (
            O => \N__26050\,
            I => \N__25857\
        );

    \I__5799\ : SRMux
    port map (
            O => \N__26049\,
            I => \N__25857\
        );

    \I__5798\ : SRMux
    port map (
            O => \N__26048\,
            I => \N__25857\
        );

    \I__5797\ : SRMux
    port map (
            O => \N__26047\,
            I => \N__25857\
        );

    \I__5796\ : SRMux
    port map (
            O => \N__26046\,
            I => \N__25857\
        );

    \I__5795\ : SRMux
    port map (
            O => \N__26045\,
            I => \N__25857\
        );

    \I__5794\ : SRMux
    port map (
            O => \N__26044\,
            I => \N__25857\
        );

    \I__5793\ : Glb2LocalMux
    port map (
            O => \N__26041\,
            I => \N__25857\
        );

    \I__5792\ : Glb2LocalMux
    port map (
            O => \N__26038\,
            I => \N__25857\
        );

    \I__5791\ : Glb2LocalMux
    port map (
            O => \N__26035\,
            I => \N__25857\
        );

    \I__5790\ : Glb2LocalMux
    port map (
            O => \N__26032\,
            I => \N__25857\
        );

    \I__5789\ : Glb2LocalMux
    port map (
            O => \N__26029\,
            I => \N__25857\
        );

    \I__5788\ : Glb2LocalMux
    port map (
            O => \N__26026\,
            I => \N__25857\
        );

    \I__5787\ : Glb2LocalMux
    port map (
            O => \N__26023\,
            I => \N__25857\
        );

    \I__5786\ : Glb2LocalMux
    port map (
            O => \N__26020\,
            I => \N__25857\
        );

    \I__5785\ : Glb2LocalMux
    port map (
            O => \N__26017\,
            I => \N__25857\
        );

    \I__5784\ : Glb2LocalMux
    port map (
            O => \N__26014\,
            I => \N__25857\
        );

    \I__5783\ : Glb2LocalMux
    port map (
            O => \N__26011\,
            I => \N__25857\
        );

    \I__5782\ : Glb2LocalMux
    port map (
            O => \N__26008\,
            I => \N__25857\
        );

    \I__5781\ : Glb2LocalMux
    port map (
            O => \N__26005\,
            I => \N__25857\
        );

    \I__5780\ : Glb2LocalMux
    port map (
            O => \N__26002\,
            I => \N__25857\
        );

    \I__5779\ : Glb2LocalMux
    port map (
            O => \N__25999\,
            I => \N__25857\
        );

    \I__5778\ : Glb2LocalMux
    port map (
            O => \N__25996\,
            I => \N__25857\
        );

    \I__5777\ : Glb2LocalMux
    port map (
            O => \N__25993\,
            I => \N__25857\
        );

    \I__5776\ : Glb2LocalMux
    port map (
            O => \N__25990\,
            I => \N__25857\
        );

    \I__5775\ : Glb2LocalMux
    port map (
            O => \N__25987\,
            I => \N__25857\
        );

    \I__5774\ : Glb2LocalMux
    port map (
            O => \N__25984\,
            I => \N__25857\
        );

    \I__5773\ : Glb2LocalMux
    port map (
            O => \N__25981\,
            I => \N__25857\
        );

    \I__5772\ : Glb2LocalMux
    port map (
            O => \N__25978\,
            I => \N__25857\
        );

    \I__5771\ : Glb2LocalMux
    port map (
            O => \N__25975\,
            I => \N__25857\
        );

    \I__5770\ : Glb2LocalMux
    port map (
            O => \N__25972\,
            I => \N__25857\
        );

    \I__5769\ : Glb2LocalMux
    port map (
            O => \N__25969\,
            I => \N__25857\
        );

    \I__5768\ : Glb2LocalMux
    port map (
            O => \N__25966\,
            I => \N__25857\
        );

    \I__5767\ : GlobalMux
    port map (
            O => \N__25857\,
            I => \N__25854\
        );

    \I__5766\ : gio2CtrlBuf
    port map (
            O => \N__25854\,
            I => \M_this_reset_cond_out_g_0\
        );

    \I__5765\ : InMux
    port map (
            O => \N__25851\,
            I => \N__25848\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__25848\,
            I => \N__25845\
        );

    \I__5763\ : Span4Mux_h
    port map (
            O => \N__25845\,
            I => \N__25842\
        );

    \I__5762\ : Odrv4
    port map (
            O => \N__25842\,
            I => \this_sprites_ram.mem_out_bus5_3\
        );

    \I__5761\ : InMux
    port map (
            O => \N__25839\,
            I => \N__25836\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__25836\,
            I => \N__25833\
        );

    \I__5759\ : Span12Mux_h
    port map (
            O => \N__25833\,
            I => \N__25830\
        );

    \I__5758\ : Span12Mux_v
    port map (
            O => \N__25830\,
            I => \N__25827\
        );

    \I__5757\ : Odrv12
    port map (
            O => \N__25827\,
            I => \this_sprites_ram.mem_out_bus1_3\
        );

    \I__5756\ : CascadeMux
    port map (
            O => \N__25824\,
            I => \N__25821\
        );

    \I__5755\ : CascadeBuf
    port map (
            O => \N__25821\,
            I => \N__25818\
        );

    \I__5754\ : CascadeMux
    port map (
            O => \N__25818\,
            I => \N__25815\
        );

    \I__5753\ : CascadeBuf
    port map (
            O => \N__25815\,
            I => \N__25812\
        );

    \I__5752\ : CascadeMux
    port map (
            O => \N__25812\,
            I => \N__25809\
        );

    \I__5751\ : CascadeBuf
    port map (
            O => \N__25809\,
            I => \N__25806\
        );

    \I__5750\ : CascadeMux
    port map (
            O => \N__25806\,
            I => \N__25803\
        );

    \I__5749\ : CascadeBuf
    port map (
            O => \N__25803\,
            I => \N__25800\
        );

    \I__5748\ : CascadeMux
    port map (
            O => \N__25800\,
            I => \N__25797\
        );

    \I__5747\ : CascadeBuf
    port map (
            O => \N__25797\,
            I => \N__25794\
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__25794\,
            I => \N__25791\
        );

    \I__5745\ : CascadeBuf
    port map (
            O => \N__25791\,
            I => \N__25788\
        );

    \I__5744\ : CascadeMux
    port map (
            O => \N__25788\,
            I => \N__25785\
        );

    \I__5743\ : CascadeBuf
    port map (
            O => \N__25785\,
            I => \N__25782\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__25782\,
            I => \N__25779\
        );

    \I__5741\ : CascadeBuf
    port map (
            O => \N__25779\,
            I => \N__25776\
        );

    \I__5740\ : CascadeMux
    port map (
            O => \N__25776\,
            I => \N__25773\
        );

    \I__5739\ : CascadeBuf
    port map (
            O => \N__25773\,
            I => \N__25770\
        );

    \I__5738\ : CascadeMux
    port map (
            O => \N__25770\,
            I => \N__25767\
        );

    \I__5737\ : CascadeBuf
    port map (
            O => \N__25767\,
            I => \N__25764\
        );

    \I__5736\ : CascadeMux
    port map (
            O => \N__25764\,
            I => \N__25761\
        );

    \I__5735\ : CascadeBuf
    port map (
            O => \N__25761\,
            I => \N__25758\
        );

    \I__5734\ : CascadeMux
    port map (
            O => \N__25758\,
            I => \N__25755\
        );

    \I__5733\ : CascadeBuf
    port map (
            O => \N__25755\,
            I => \N__25752\
        );

    \I__5732\ : CascadeMux
    port map (
            O => \N__25752\,
            I => \N__25749\
        );

    \I__5731\ : CascadeBuf
    port map (
            O => \N__25749\,
            I => \N__25746\
        );

    \I__5730\ : CascadeMux
    port map (
            O => \N__25746\,
            I => \N__25743\
        );

    \I__5729\ : CascadeBuf
    port map (
            O => \N__25743\,
            I => \N__25740\
        );

    \I__5728\ : CascadeMux
    port map (
            O => \N__25740\,
            I => \N__25737\
        );

    \I__5727\ : CascadeBuf
    port map (
            O => \N__25737\,
            I => \N__25734\
        );

    \I__5726\ : CascadeMux
    port map (
            O => \N__25734\,
            I => \N__25731\
        );

    \I__5725\ : InMux
    port map (
            O => \N__25731\,
            I => \N__25728\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__25728\,
            I => \N__25725\
        );

    \I__5723\ : Span4Mux_h
    port map (
            O => \N__25725\,
            I => \N__25722\
        );

    \I__5722\ : Sp12to4
    port map (
            O => \N__25722\,
            I => \N__25716\
        );

    \I__5721\ : InMux
    port map (
            O => \N__25721\,
            I => \N__25713\
        );

    \I__5720\ : InMux
    port map (
            O => \N__25720\,
            I => \N__25708\
        );

    \I__5719\ : InMux
    port map (
            O => \N__25719\,
            I => \N__25708\
        );

    \I__5718\ : Span12Mux_s6_v
    port map (
            O => \N__25716\,
            I => \N__25705\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__25713\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__25708\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__5715\ : Odrv12
    port map (
            O => \N__25705\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__5714\ : InMux
    port map (
            O => \N__25698\,
            I => \N__25695\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__25695\,
            I => \un1_M_this_sprites_address_q_cry_5_THRU_CO\
        );

    \I__5712\ : InMux
    port map (
            O => \N__25692\,
            I => \un1_M_this_sprites_address_q_cry_5\
        );

    \I__5711\ : CascadeMux
    port map (
            O => \N__25689\,
            I => \N__25686\
        );

    \I__5710\ : CascadeBuf
    port map (
            O => \N__25686\,
            I => \N__25683\
        );

    \I__5709\ : CascadeMux
    port map (
            O => \N__25683\,
            I => \N__25680\
        );

    \I__5708\ : CascadeBuf
    port map (
            O => \N__25680\,
            I => \N__25677\
        );

    \I__5707\ : CascadeMux
    port map (
            O => \N__25677\,
            I => \N__25674\
        );

    \I__5706\ : CascadeBuf
    port map (
            O => \N__25674\,
            I => \N__25671\
        );

    \I__5705\ : CascadeMux
    port map (
            O => \N__25671\,
            I => \N__25668\
        );

    \I__5704\ : CascadeBuf
    port map (
            O => \N__25668\,
            I => \N__25665\
        );

    \I__5703\ : CascadeMux
    port map (
            O => \N__25665\,
            I => \N__25662\
        );

    \I__5702\ : CascadeBuf
    port map (
            O => \N__25662\,
            I => \N__25659\
        );

    \I__5701\ : CascadeMux
    port map (
            O => \N__25659\,
            I => \N__25656\
        );

    \I__5700\ : CascadeBuf
    port map (
            O => \N__25656\,
            I => \N__25653\
        );

    \I__5699\ : CascadeMux
    port map (
            O => \N__25653\,
            I => \N__25650\
        );

    \I__5698\ : CascadeBuf
    port map (
            O => \N__25650\,
            I => \N__25647\
        );

    \I__5697\ : CascadeMux
    port map (
            O => \N__25647\,
            I => \N__25644\
        );

    \I__5696\ : CascadeBuf
    port map (
            O => \N__25644\,
            I => \N__25641\
        );

    \I__5695\ : CascadeMux
    port map (
            O => \N__25641\,
            I => \N__25638\
        );

    \I__5694\ : CascadeBuf
    port map (
            O => \N__25638\,
            I => \N__25635\
        );

    \I__5693\ : CascadeMux
    port map (
            O => \N__25635\,
            I => \N__25632\
        );

    \I__5692\ : CascadeBuf
    port map (
            O => \N__25632\,
            I => \N__25629\
        );

    \I__5691\ : CascadeMux
    port map (
            O => \N__25629\,
            I => \N__25626\
        );

    \I__5690\ : CascadeBuf
    port map (
            O => \N__25626\,
            I => \N__25623\
        );

    \I__5689\ : CascadeMux
    port map (
            O => \N__25623\,
            I => \N__25620\
        );

    \I__5688\ : CascadeBuf
    port map (
            O => \N__25620\,
            I => \N__25617\
        );

    \I__5687\ : CascadeMux
    port map (
            O => \N__25617\,
            I => \N__25614\
        );

    \I__5686\ : CascadeBuf
    port map (
            O => \N__25614\,
            I => \N__25611\
        );

    \I__5685\ : CascadeMux
    port map (
            O => \N__25611\,
            I => \N__25608\
        );

    \I__5684\ : CascadeBuf
    port map (
            O => \N__25608\,
            I => \N__25605\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__25605\,
            I => \N__25602\
        );

    \I__5682\ : CascadeBuf
    port map (
            O => \N__25602\,
            I => \N__25599\
        );

    \I__5681\ : CascadeMux
    port map (
            O => \N__25599\,
            I => \N__25596\
        );

    \I__5680\ : InMux
    port map (
            O => \N__25596\,
            I => \N__25593\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__25593\,
            I => \N__25590\
        );

    \I__5678\ : Span4Mux_h
    port map (
            O => \N__25590\,
            I => \N__25585\
        );

    \I__5677\ : CascadeMux
    port map (
            O => \N__25589\,
            I => \N__25582\
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__25588\,
            I => \N__25579\
        );

    \I__5675\ : Sp12to4
    port map (
            O => \N__25585\,
            I => \N__25575\
        );

    \I__5674\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25572\
        );

    \I__5673\ : InMux
    port map (
            O => \N__25579\,
            I => \N__25569\
        );

    \I__5672\ : InMux
    port map (
            O => \N__25578\,
            I => \N__25566\
        );

    \I__5671\ : Span12Mux_s8_v
    port map (
            O => \N__25575\,
            I => \N__25563\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__25572\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__25569\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__25566\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5667\ : Odrv12
    port map (
            O => \N__25563\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5666\ : InMux
    port map (
            O => \N__25554\,
            I => \N__25551\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__25551\,
            I => \un1_M_this_sprites_address_q_cry_6_THRU_CO\
        );

    \I__5664\ : InMux
    port map (
            O => \N__25548\,
            I => \un1_M_this_sprites_address_q_cry_6\
        );

    \I__5663\ : InMux
    port map (
            O => \N__25545\,
            I => \bfn_23_18_0_\
        );

    \I__5662\ : InMux
    port map (
            O => \N__25542\,
            I => \un1_M_this_sprites_address_q_cry_8\
        );

    \I__5661\ : CascadeMux
    port map (
            O => \N__25539\,
            I => \N__25536\
        );

    \I__5660\ : CascadeBuf
    port map (
            O => \N__25536\,
            I => \N__25533\
        );

    \I__5659\ : CascadeMux
    port map (
            O => \N__25533\,
            I => \N__25530\
        );

    \I__5658\ : CascadeBuf
    port map (
            O => \N__25530\,
            I => \N__25527\
        );

    \I__5657\ : CascadeMux
    port map (
            O => \N__25527\,
            I => \N__25524\
        );

    \I__5656\ : CascadeBuf
    port map (
            O => \N__25524\,
            I => \N__25521\
        );

    \I__5655\ : CascadeMux
    port map (
            O => \N__25521\,
            I => \N__25518\
        );

    \I__5654\ : CascadeBuf
    port map (
            O => \N__25518\,
            I => \N__25515\
        );

    \I__5653\ : CascadeMux
    port map (
            O => \N__25515\,
            I => \N__25512\
        );

    \I__5652\ : CascadeBuf
    port map (
            O => \N__25512\,
            I => \N__25509\
        );

    \I__5651\ : CascadeMux
    port map (
            O => \N__25509\,
            I => \N__25506\
        );

    \I__5650\ : CascadeBuf
    port map (
            O => \N__25506\,
            I => \N__25503\
        );

    \I__5649\ : CascadeMux
    port map (
            O => \N__25503\,
            I => \N__25500\
        );

    \I__5648\ : CascadeBuf
    port map (
            O => \N__25500\,
            I => \N__25497\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__25497\,
            I => \N__25494\
        );

    \I__5646\ : CascadeBuf
    port map (
            O => \N__25494\,
            I => \N__25491\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__25491\,
            I => \N__25488\
        );

    \I__5644\ : CascadeBuf
    port map (
            O => \N__25488\,
            I => \N__25485\
        );

    \I__5643\ : CascadeMux
    port map (
            O => \N__25485\,
            I => \N__25482\
        );

    \I__5642\ : CascadeBuf
    port map (
            O => \N__25482\,
            I => \N__25479\
        );

    \I__5641\ : CascadeMux
    port map (
            O => \N__25479\,
            I => \N__25476\
        );

    \I__5640\ : CascadeBuf
    port map (
            O => \N__25476\,
            I => \N__25473\
        );

    \I__5639\ : CascadeMux
    port map (
            O => \N__25473\,
            I => \N__25470\
        );

    \I__5638\ : CascadeBuf
    port map (
            O => \N__25470\,
            I => \N__25467\
        );

    \I__5637\ : CascadeMux
    port map (
            O => \N__25467\,
            I => \N__25464\
        );

    \I__5636\ : CascadeBuf
    port map (
            O => \N__25464\,
            I => \N__25461\
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__25461\,
            I => \N__25458\
        );

    \I__5634\ : CascadeBuf
    port map (
            O => \N__25458\,
            I => \N__25455\
        );

    \I__5633\ : CascadeMux
    port map (
            O => \N__25455\,
            I => \N__25452\
        );

    \I__5632\ : CascadeBuf
    port map (
            O => \N__25452\,
            I => \N__25449\
        );

    \I__5631\ : CascadeMux
    port map (
            O => \N__25449\,
            I => \N__25446\
        );

    \I__5630\ : InMux
    port map (
            O => \N__25446\,
            I => \N__25443\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__25443\,
            I => \N__25440\
        );

    \I__5628\ : Span4Mux_h
    port map (
            O => \N__25440\,
            I => \N__25437\
        );

    \I__5627\ : Sp12to4
    port map (
            O => \N__25437\,
            I => \N__25431\
        );

    \I__5626\ : InMux
    port map (
            O => \N__25436\,
            I => \N__25428\
        );

    \I__5625\ : InMux
    port map (
            O => \N__25435\,
            I => \N__25423\
        );

    \I__5624\ : InMux
    port map (
            O => \N__25434\,
            I => \N__25423\
        );

    \I__5623\ : Span12Mux_s5_v
    port map (
            O => \N__25431\,
            I => \N__25420\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__25428\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__25423\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5620\ : Odrv12
    port map (
            O => \N__25420\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5619\ : InMux
    port map (
            O => \N__25413\,
            I => \N__25410\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__25410\,
            I => \un1_M_this_sprites_address_q_cry_9_THRU_CO\
        );

    \I__5617\ : InMux
    port map (
            O => \N__25407\,
            I => \un1_M_this_sprites_address_q_cry_9\
        );

    \I__5616\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25401\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__25401\,
            I => \un1_M_this_sprites_address_q_cry_10_THRU_CO\
        );

    \I__5614\ : InMux
    port map (
            O => \N__25398\,
            I => \un1_M_this_sprites_address_q_cry_10\
        );

    \I__5613\ : InMux
    port map (
            O => \N__25395\,
            I => \N__25392\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__25392\,
            I => \un1_M_this_sprites_address_q_cry_11_THRU_CO\
        );

    \I__5611\ : InMux
    port map (
            O => \N__25389\,
            I => \un1_M_this_sprites_address_q_cry_11\
        );

    \I__5610\ : InMux
    port map (
            O => \N__25386\,
            I => \N__25383\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__25383\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_13\
        );

    \I__5608\ : InMux
    port map (
            O => \N__25380\,
            I => \un1_M_this_sprites_address_q_cry_12\
        );

    \I__5607\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25374\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__25374\,
            I => \N__25371\
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__25371\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_0\
        );

    \I__5604\ : InMux
    port map (
            O => \N__25368\,
            I => \N__25364\
        );

    \I__5603\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25361\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__25364\,
            I => un30_0
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__25361\,
            I => un30_0
        );

    \I__5600\ : CascadeMux
    port map (
            O => \N__25356\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_1_cascade_\
        );

    \I__5599\ : InMux
    port map (
            O => \N__25353\,
            I => \N__25347\
        );

    \I__5598\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25347\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__25347\,
            I => \N__25340\
        );

    \I__5596\ : InMux
    port map (
            O => \N__25346\,
            I => \N__25331\
        );

    \I__5595\ : InMux
    port map (
            O => \N__25345\,
            I => \N__25331\
        );

    \I__5594\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25331\
        );

    \I__5593\ : InMux
    port map (
            O => \N__25343\,
            I => \N__25331\
        );

    \I__5592\ : Span4Mux_v
    port map (
            O => \N__25340\,
            I => \N__25327\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__25331\,
            I => \N__25324\
        );

    \I__5590\ : InMux
    port map (
            O => \N__25330\,
            I => \N__25321\
        );

    \I__5589\ : Odrv4
    port map (
            O => \N__25327\,
            I => \this_start_data_delay.N_993\
        );

    \I__5588\ : Odrv4
    port map (
            O => \N__25324\,
            I => \this_start_data_delay.N_993\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__25321\,
            I => \this_start_data_delay.N_993\
        );

    \I__5586\ : CascadeMux
    port map (
            O => \N__25314\,
            I => \N__25309\
        );

    \I__5585\ : CascadeMux
    port map (
            O => \N__25313\,
            I => \N__25306\
        );

    \I__5584\ : CascadeMux
    port map (
            O => \N__25312\,
            I => \N__25303\
        );

    \I__5583\ : InMux
    port map (
            O => \N__25309\,
            I => \N__25291\
        );

    \I__5582\ : InMux
    port map (
            O => \N__25306\,
            I => \N__25291\
        );

    \I__5581\ : InMux
    port map (
            O => \N__25303\,
            I => \N__25291\
        );

    \I__5580\ : InMux
    port map (
            O => \N__25302\,
            I => \N__25291\
        );

    \I__5579\ : InMux
    port map (
            O => \N__25301\,
            I => \N__25286\
        );

    \I__5578\ : InMux
    port map (
            O => \N__25300\,
            I => \N__25286\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__25291\,
            I => \N__25283\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__25286\,
            I => \N__25280\
        );

    \I__5575\ : Span4Mux_v
    port map (
            O => \N__25283\,
            I => \N__25277\
        );

    \I__5574\ : Odrv4
    port map (
            O => \N__25280\,
            I => \this_start_data_delay.N_109\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__25277\,
            I => \this_start_data_delay.N_109\
        );

    \I__5572\ : CascadeMux
    port map (
            O => \N__25272\,
            I => \N__25269\
        );

    \I__5571\ : CascadeBuf
    port map (
            O => \N__25269\,
            I => \N__25266\
        );

    \I__5570\ : CascadeMux
    port map (
            O => \N__25266\,
            I => \N__25263\
        );

    \I__5569\ : CascadeBuf
    port map (
            O => \N__25263\,
            I => \N__25260\
        );

    \I__5568\ : CascadeMux
    port map (
            O => \N__25260\,
            I => \N__25257\
        );

    \I__5567\ : CascadeBuf
    port map (
            O => \N__25257\,
            I => \N__25254\
        );

    \I__5566\ : CascadeMux
    port map (
            O => \N__25254\,
            I => \N__25251\
        );

    \I__5565\ : CascadeBuf
    port map (
            O => \N__25251\,
            I => \N__25248\
        );

    \I__5564\ : CascadeMux
    port map (
            O => \N__25248\,
            I => \N__25245\
        );

    \I__5563\ : CascadeBuf
    port map (
            O => \N__25245\,
            I => \N__25242\
        );

    \I__5562\ : CascadeMux
    port map (
            O => \N__25242\,
            I => \N__25239\
        );

    \I__5561\ : CascadeBuf
    port map (
            O => \N__25239\,
            I => \N__25236\
        );

    \I__5560\ : CascadeMux
    port map (
            O => \N__25236\,
            I => \N__25233\
        );

    \I__5559\ : CascadeBuf
    port map (
            O => \N__25233\,
            I => \N__25230\
        );

    \I__5558\ : CascadeMux
    port map (
            O => \N__25230\,
            I => \N__25227\
        );

    \I__5557\ : CascadeBuf
    port map (
            O => \N__25227\,
            I => \N__25224\
        );

    \I__5556\ : CascadeMux
    port map (
            O => \N__25224\,
            I => \N__25221\
        );

    \I__5555\ : CascadeBuf
    port map (
            O => \N__25221\,
            I => \N__25218\
        );

    \I__5554\ : CascadeMux
    port map (
            O => \N__25218\,
            I => \N__25215\
        );

    \I__5553\ : CascadeBuf
    port map (
            O => \N__25215\,
            I => \N__25212\
        );

    \I__5552\ : CascadeMux
    port map (
            O => \N__25212\,
            I => \N__25209\
        );

    \I__5551\ : CascadeBuf
    port map (
            O => \N__25209\,
            I => \N__25206\
        );

    \I__5550\ : CascadeMux
    port map (
            O => \N__25206\,
            I => \N__25203\
        );

    \I__5549\ : CascadeBuf
    port map (
            O => \N__25203\,
            I => \N__25200\
        );

    \I__5548\ : CascadeMux
    port map (
            O => \N__25200\,
            I => \N__25197\
        );

    \I__5547\ : CascadeBuf
    port map (
            O => \N__25197\,
            I => \N__25194\
        );

    \I__5546\ : CascadeMux
    port map (
            O => \N__25194\,
            I => \N__25191\
        );

    \I__5545\ : CascadeBuf
    port map (
            O => \N__25191\,
            I => \N__25188\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__25188\,
            I => \N__25185\
        );

    \I__5543\ : CascadeBuf
    port map (
            O => \N__25185\,
            I => \N__25182\
        );

    \I__5542\ : CascadeMux
    port map (
            O => \N__25182\,
            I => \N__25179\
        );

    \I__5541\ : InMux
    port map (
            O => \N__25179\,
            I => \N__25176\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__25176\,
            I => \N__25172\
        );

    \I__5539\ : CascadeMux
    port map (
            O => \N__25175\,
            I => \N__25169\
        );

    \I__5538\ : Span12Mux_s4_v
    port map (
            O => \N__25172\,
            I => \N__25164\
        );

    \I__5537\ : InMux
    port map (
            O => \N__25169\,
            I => \N__25161\
        );

    \I__5536\ : InMux
    port map (
            O => \N__25168\,
            I => \N__25156\
        );

    \I__5535\ : InMux
    port map (
            O => \N__25167\,
            I => \N__25156\
        );

    \I__5534\ : Span12Mux_v
    port map (
            O => \N__25164\,
            I => \N__25153\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__25161\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__25156\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__5531\ : Odrv12
    port map (
            O => \N__25153\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__5530\ : InMux
    port map (
            O => \N__25146\,
            I => \N__25143\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__25143\,
            I => \un1_M_this_sprites_address_q_cry_0_THRU_CO\
        );

    \I__5528\ : InMux
    port map (
            O => \N__25140\,
            I => \un1_M_this_sprites_address_q_cry_0\
        );

    \I__5527\ : CascadeMux
    port map (
            O => \N__25137\,
            I => \N__25134\
        );

    \I__5526\ : CascadeBuf
    port map (
            O => \N__25134\,
            I => \N__25131\
        );

    \I__5525\ : CascadeMux
    port map (
            O => \N__25131\,
            I => \N__25128\
        );

    \I__5524\ : CascadeBuf
    port map (
            O => \N__25128\,
            I => \N__25125\
        );

    \I__5523\ : CascadeMux
    port map (
            O => \N__25125\,
            I => \N__25122\
        );

    \I__5522\ : CascadeBuf
    port map (
            O => \N__25122\,
            I => \N__25119\
        );

    \I__5521\ : CascadeMux
    port map (
            O => \N__25119\,
            I => \N__25116\
        );

    \I__5520\ : CascadeBuf
    port map (
            O => \N__25116\,
            I => \N__25113\
        );

    \I__5519\ : CascadeMux
    port map (
            O => \N__25113\,
            I => \N__25110\
        );

    \I__5518\ : CascadeBuf
    port map (
            O => \N__25110\,
            I => \N__25107\
        );

    \I__5517\ : CascadeMux
    port map (
            O => \N__25107\,
            I => \N__25104\
        );

    \I__5516\ : CascadeBuf
    port map (
            O => \N__25104\,
            I => \N__25101\
        );

    \I__5515\ : CascadeMux
    port map (
            O => \N__25101\,
            I => \N__25098\
        );

    \I__5514\ : CascadeBuf
    port map (
            O => \N__25098\,
            I => \N__25095\
        );

    \I__5513\ : CascadeMux
    port map (
            O => \N__25095\,
            I => \N__25092\
        );

    \I__5512\ : CascadeBuf
    port map (
            O => \N__25092\,
            I => \N__25089\
        );

    \I__5511\ : CascadeMux
    port map (
            O => \N__25089\,
            I => \N__25086\
        );

    \I__5510\ : CascadeBuf
    port map (
            O => \N__25086\,
            I => \N__25083\
        );

    \I__5509\ : CascadeMux
    port map (
            O => \N__25083\,
            I => \N__25080\
        );

    \I__5508\ : CascadeBuf
    port map (
            O => \N__25080\,
            I => \N__25077\
        );

    \I__5507\ : CascadeMux
    port map (
            O => \N__25077\,
            I => \N__25074\
        );

    \I__5506\ : CascadeBuf
    port map (
            O => \N__25074\,
            I => \N__25071\
        );

    \I__5505\ : CascadeMux
    port map (
            O => \N__25071\,
            I => \N__25068\
        );

    \I__5504\ : CascadeBuf
    port map (
            O => \N__25068\,
            I => \N__25065\
        );

    \I__5503\ : CascadeMux
    port map (
            O => \N__25065\,
            I => \N__25062\
        );

    \I__5502\ : CascadeBuf
    port map (
            O => \N__25062\,
            I => \N__25059\
        );

    \I__5501\ : CascadeMux
    port map (
            O => \N__25059\,
            I => \N__25056\
        );

    \I__5500\ : CascadeBuf
    port map (
            O => \N__25056\,
            I => \N__25053\
        );

    \I__5499\ : CascadeMux
    port map (
            O => \N__25053\,
            I => \N__25050\
        );

    \I__5498\ : CascadeBuf
    port map (
            O => \N__25050\,
            I => \N__25047\
        );

    \I__5497\ : CascadeMux
    port map (
            O => \N__25047\,
            I => \N__25044\
        );

    \I__5496\ : InMux
    port map (
            O => \N__25044\,
            I => \N__25041\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__25041\,
            I => \N__25037\
        );

    \I__5494\ : InMux
    port map (
            O => \N__25040\,
            I => \N__25034\
        );

    \I__5493\ : Span12Mux_s10_h
    port map (
            O => \N__25037\,
            I => \N__25029\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__25034\,
            I => \N__25026\
        );

    \I__5491\ : InMux
    port map (
            O => \N__25033\,
            I => \N__25023\
        );

    \I__5490\ : InMux
    port map (
            O => \N__25032\,
            I => \N__25020\
        );

    \I__5489\ : Span12Mux_v
    port map (
            O => \N__25029\,
            I => \N__25017\
        );

    \I__5488\ : Odrv4
    port map (
            O => \N__25026\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__25023\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__25020\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__5485\ : Odrv12
    port map (
            O => \N__25017\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__5484\ : InMux
    port map (
            O => \N__25008\,
            I => \N__25005\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__25005\,
            I => \N__25002\
        );

    \I__5482\ : Odrv4
    port map (
            O => \N__25002\,
            I => \un1_M_this_sprites_address_q_cry_1_THRU_CO\
        );

    \I__5481\ : InMux
    port map (
            O => \N__24999\,
            I => \un1_M_this_sprites_address_q_cry_1\
        );

    \I__5480\ : CascadeMux
    port map (
            O => \N__24996\,
            I => \N__24993\
        );

    \I__5479\ : CascadeBuf
    port map (
            O => \N__24993\,
            I => \N__24990\
        );

    \I__5478\ : CascadeMux
    port map (
            O => \N__24990\,
            I => \N__24987\
        );

    \I__5477\ : CascadeBuf
    port map (
            O => \N__24987\,
            I => \N__24984\
        );

    \I__5476\ : CascadeMux
    port map (
            O => \N__24984\,
            I => \N__24981\
        );

    \I__5475\ : CascadeBuf
    port map (
            O => \N__24981\,
            I => \N__24978\
        );

    \I__5474\ : CascadeMux
    port map (
            O => \N__24978\,
            I => \N__24975\
        );

    \I__5473\ : CascadeBuf
    port map (
            O => \N__24975\,
            I => \N__24972\
        );

    \I__5472\ : CascadeMux
    port map (
            O => \N__24972\,
            I => \N__24969\
        );

    \I__5471\ : CascadeBuf
    port map (
            O => \N__24969\,
            I => \N__24966\
        );

    \I__5470\ : CascadeMux
    port map (
            O => \N__24966\,
            I => \N__24963\
        );

    \I__5469\ : CascadeBuf
    port map (
            O => \N__24963\,
            I => \N__24960\
        );

    \I__5468\ : CascadeMux
    port map (
            O => \N__24960\,
            I => \N__24957\
        );

    \I__5467\ : CascadeBuf
    port map (
            O => \N__24957\,
            I => \N__24954\
        );

    \I__5466\ : CascadeMux
    port map (
            O => \N__24954\,
            I => \N__24951\
        );

    \I__5465\ : CascadeBuf
    port map (
            O => \N__24951\,
            I => \N__24948\
        );

    \I__5464\ : CascadeMux
    port map (
            O => \N__24948\,
            I => \N__24945\
        );

    \I__5463\ : CascadeBuf
    port map (
            O => \N__24945\,
            I => \N__24942\
        );

    \I__5462\ : CascadeMux
    port map (
            O => \N__24942\,
            I => \N__24939\
        );

    \I__5461\ : CascadeBuf
    port map (
            O => \N__24939\,
            I => \N__24936\
        );

    \I__5460\ : CascadeMux
    port map (
            O => \N__24936\,
            I => \N__24933\
        );

    \I__5459\ : CascadeBuf
    port map (
            O => \N__24933\,
            I => \N__24930\
        );

    \I__5458\ : CascadeMux
    port map (
            O => \N__24930\,
            I => \N__24927\
        );

    \I__5457\ : CascadeBuf
    port map (
            O => \N__24927\,
            I => \N__24924\
        );

    \I__5456\ : CascadeMux
    port map (
            O => \N__24924\,
            I => \N__24921\
        );

    \I__5455\ : CascadeBuf
    port map (
            O => \N__24921\,
            I => \N__24918\
        );

    \I__5454\ : CascadeMux
    port map (
            O => \N__24918\,
            I => \N__24915\
        );

    \I__5453\ : CascadeBuf
    port map (
            O => \N__24915\,
            I => \N__24912\
        );

    \I__5452\ : CascadeMux
    port map (
            O => \N__24912\,
            I => \N__24909\
        );

    \I__5451\ : CascadeBuf
    port map (
            O => \N__24909\,
            I => \N__24906\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__24906\,
            I => \N__24903\
        );

    \I__5449\ : InMux
    port map (
            O => \N__24903\,
            I => \N__24899\
        );

    \I__5448\ : InMux
    port map (
            O => \N__24902\,
            I => \N__24896\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__24899\,
            I => \N__24893\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__24896\,
            I => \N__24890\
        );

    \I__5445\ : Span12Mux_s1_v
    port map (
            O => \N__24893\,
            I => \N__24885\
        );

    \I__5444\ : Span4Mux_h
    port map (
            O => \N__24890\,
            I => \N__24882\
        );

    \I__5443\ : InMux
    port map (
            O => \N__24889\,
            I => \N__24879\
        );

    \I__5442\ : InMux
    port map (
            O => \N__24888\,
            I => \N__24876\
        );

    \I__5441\ : Span12Mux_v
    port map (
            O => \N__24885\,
            I => \N__24873\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__24882\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__24879\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__24876\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5437\ : Odrv12
    port map (
            O => \N__24873\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5436\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24861\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__24861\,
            I => \N__24858\
        );

    \I__5434\ : Odrv4
    port map (
            O => \N__24858\,
            I => \un1_M_this_sprites_address_q_cry_2_THRU_CO\
        );

    \I__5433\ : InMux
    port map (
            O => \N__24855\,
            I => \un1_M_this_sprites_address_q_cry_2\
        );

    \I__5432\ : CascadeMux
    port map (
            O => \N__24852\,
            I => \N__24849\
        );

    \I__5431\ : CascadeBuf
    port map (
            O => \N__24849\,
            I => \N__24846\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__24846\,
            I => \N__24843\
        );

    \I__5429\ : CascadeBuf
    port map (
            O => \N__24843\,
            I => \N__24840\
        );

    \I__5428\ : CascadeMux
    port map (
            O => \N__24840\,
            I => \N__24837\
        );

    \I__5427\ : CascadeBuf
    port map (
            O => \N__24837\,
            I => \N__24834\
        );

    \I__5426\ : CascadeMux
    port map (
            O => \N__24834\,
            I => \N__24831\
        );

    \I__5425\ : CascadeBuf
    port map (
            O => \N__24831\,
            I => \N__24828\
        );

    \I__5424\ : CascadeMux
    port map (
            O => \N__24828\,
            I => \N__24825\
        );

    \I__5423\ : CascadeBuf
    port map (
            O => \N__24825\,
            I => \N__24822\
        );

    \I__5422\ : CascadeMux
    port map (
            O => \N__24822\,
            I => \N__24819\
        );

    \I__5421\ : CascadeBuf
    port map (
            O => \N__24819\,
            I => \N__24816\
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__24816\,
            I => \N__24813\
        );

    \I__5419\ : CascadeBuf
    port map (
            O => \N__24813\,
            I => \N__24810\
        );

    \I__5418\ : CascadeMux
    port map (
            O => \N__24810\,
            I => \N__24807\
        );

    \I__5417\ : CascadeBuf
    port map (
            O => \N__24807\,
            I => \N__24804\
        );

    \I__5416\ : CascadeMux
    port map (
            O => \N__24804\,
            I => \N__24801\
        );

    \I__5415\ : CascadeBuf
    port map (
            O => \N__24801\,
            I => \N__24798\
        );

    \I__5414\ : CascadeMux
    port map (
            O => \N__24798\,
            I => \N__24795\
        );

    \I__5413\ : CascadeBuf
    port map (
            O => \N__24795\,
            I => \N__24792\
        );

    \I__5412\ : CascadeMux
    port map (
            O => \N__24792\,
            I => \N__24789\
        );

    \I__5411\ : CascadeBuf
    port map (
            O => \N__24789\,
            I => \N__24786\
        );

    \I__5410\ : CascadeMux
    port map (
            O => \N__24786\,
            I => \N__24783\
        );

    \I__5409\ : CascadeBuf
    port map (
            O => \N__24783\,
            I => \N__24780\
        );

    \I__5408\ : CascadeMux
    port map (
            O => \N__24780\,
            I => \N__24777\
        );

    \I__5407\ : CascadeBuf
    port map (
            O => \N__24777\,
            I => \N__24774\
        );

    \I__5406\ : CascadeMux
    port map (
            O => \N__24774\,
            I => \N__24771\
        );

    \I__5405\ : CascadeBuf
    port map (
            O => \N__24771\,
            I => \N__24768\
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__24768\,
            I => \N__24765\
        );

    \I__5403\ : CascadeBuf
    port map (
            O => \N__24765\,
            I => \N__24762\
        );

    \I__5402\ : CascadeMux
    port map (
            O => \N__24762\,
            I => \N__24759\
        );

    \I__5401\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24756\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__24756\,
            I => \N__24753\
        );

    \I__5399\ : Span4Mux_s3_v
    port map (
            O => \N__24753\,
            I => \N__24749\
        );

    \I__5398\ : InMux
    port map (
            O => \N__24752\,
            I => \N__24746\
        );

    \I__5397\ : Span4Mux_v
    port map (
            O => \N__24749\,
            I => \N__24741\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__24746\,
            I => \N__24738\
        );

    \I__5395\ : InMux
    port map (
            O => \N__24745\,
            I => \N__24735\
        );

    \I__5394\ : CascadeMux
    port map (
            O => \N__24744\,
            I => \N__24732\
        );

    \I__5393\ : Sp12to4
    port map (
            O => \N__24741\,
            I => \N__24729\
        );

    \I__5392\ : Span4Mux_h
    port map (
            O => \N__24738\,
            I => \N__24726\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__24735\,
            I => \N__24723\
        );

    \I__5390\ : InMux
    port map (
            O => \N__24732\,
            I => \N__24720\
        );

    \I__5389\ : Span12Mux_v
    port map (
            O => \N__24729\,
            I => \N__24717\
        );

    \I__5388\ : Odrv4
    port map (
            O => \N__24726\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__24723\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__24720\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__5385\ : Odrv12
    port map (
            O => \N__24717\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__5384\ : InMux
    port map (
            O => \N__24708\,
            I => \N__24705\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__24705\,
            I => \N__24702\
        );

    \I__5382\ : Span4Mux_h
    port map (
            O => \N__24702\,
            I => \N__24699\
        );

    \I__5381\ : Odrv4
    port map (
            O => \N__24699\,
            I => \un1_M_this_sprites_address_q_cry_3_THRU_CO\
        );

    \I__5380\ : InMux
    port map (
            O => \N__24696\,
            I => \un1_M_this_sprites_address_q_cry_3\
        );

    \I__5379\ : InMux
    port map (
            O => \N__24693\,
            I => \un1_M_this_sprites_address_q_cry_4\
        );

    \I__5378\ : InMux
    port map (
            O => \N__24690\,
            I => \N__24687\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__24687\,
            I => \N__24684\
        );

    \I__5376\ : Span4Mux_h
    port map (
            O => \N__24684\,
            I => \N__24681\
        );

    \I__5375\ : Span4Mux_v
    port map (
            O => \N__24681\,
            I => \N__24677\
        );

    \I__5374\ : InMux
    port map (
            O => \N__24680\,
            I => \N__24674\
        );

    \I__5373\ : Odrv4
    port map (
            O => \N__24677\,
            I => \this_start_data_delay.N_93_0\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__24674\,
            I => \this_start_data_delay.N_93_0\
        );

    \I__5371\ : InMux
    port map (
            O => \N__24669\,
            I => \N__24666\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__24666\,
            I => \N__24663\
        );

    \I__5369\ : Span4Mux_v
    port map (
            O => \N__24663\,
            I => \N__24660\
        );

    \I__5368\ : Span4Mux_v
    port map (
            O => \N__24660\,
            I => \N__24657\
        );

    \I__5367\ : Odrv4
    port map (
            O => \N__24657\,
            I => \this_start_data_delay.N_122\
        );

    \I__5366\ : CascadeMux
    port map (
            O => \N__24654\,
            I => \N__24651\
        );

    \I__5365\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24648\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__24648\,
            I => \N__24644\
        );

    \I__5363\ : InMux
    port map (
            O => \N__24647\,
            I => \N__24641\
        );

    \I__5362\ : Odrv12
    port map (
            O => \N__24644\,
            I => \this_start_data_delay.N_149\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__24641\,
            I => \this_start_data_delay.N_149\
        );

    \I__5360\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24633\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__24633\,
            I => \N__24630\
        );

    \I__5358\ : Span4Mux_v
    port map (
            O => \N__24630\,
            I => \N__24627\
        );

    \I__5357\ : Odrv4
    port map (
            O => \N__24627\,
            I => \this_start_data_delay.N_121\
        );

    \I__5356\ : InMux
    port map (
            O => \N__24624\,
            I => \N__24619\
        );

    \I__5355\ : InMux
    port map (
            O => \N__24623\,
            I => \N__24616\
        );

    \I__5354\ : InMux
    port map (
            O => \N__24622\,
            I => \N__24613\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__24619\,
            I => \N__24610\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__24616\,
            I => \N__24605\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__24613\,
            I => \N__24600\
        );

    \I__5350\ : Span4Mux_h
    port map (
            O => \N__24610\,
            I => \N__24600\
        );

    \I__5349\ : InMux
    port map (
            O => \N__24609\,
            I => \N__24597\
        );

    \I__5348\ : InMux
    port map (
            O => \N__24608\,
            I => \N__24594\
        );

    \I__5347\ : Odrv12
    port map (
            O => \N__24605\,
            I => \this_start_data_delay.N_938_0\
        );

    \I__5346\ : Odrv4
    port map (
            O => \N__24600\,
            I => \this_start_data_delay.N_938_0\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__24597\,
            I => \this_start_data_delay.N_938_0\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__24594\,
            I => \this_start_data_delay.N_938_0\
        );

    \I__5343\ : InMux
    port map (
            O => \N__24585\,
            I => \N__24581\
        );

    \I__5342\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24577\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__24581\,
            I => \N__24573\
        );

    \I__5340\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24570\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__24577\,
            I => \N__24566\
        );

    \I__5338\ : InMux
    port map (
            O => \N__24576\,
            I => \N__24563\
        );

    \I__5337\ : Span4Mux_v
    port map (
            O => \N__24573\,
            I => \N__24557\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__24570\,
            I => \N__24557\
        );

    \I__5335\ : InMux
    port map (
            O => \N__24569\,
            I => \N__24554\
        );

    \I__5334\ : Span4Mux_s2_v
    port map (
            O => \N__24566\,
            I => \N__24548\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__24563\,
            I => \N__24548\
        );

    \I__5332\ : InMux
    port map (
            O => \N__24562\,
            I => \N__24545\
        );

    \I__5331\ : Span4Mux_v
    port map (
            O => \N__24557\,
            I => \N__24541\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__24554\,
            I => \N__24538\
        );

    \I__5329\ : InMux
    port map (
            O => \N__24553\,
            I => \N__24535\
        );

    \I__5328\ : Span4Mux_v
    port map (
            O => \N__24548\,
            I => \N__24530\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__24545\,
            I => \N__24530\
        );

    \I__5326\ : InMux
    port map (
            O => \N__24544\,
            I => \N__24527\
        );

    \I__5325\ : Span4Mux_v
    port map (
            O => \N__24541\,
            I => \N__24520\
        );

    \I__5324\ : Span4Mux_v
    port map (
            O => \N__24538\,
            I => \N__24520\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__24535\,
            I => \N__24520\
        );

    \I__5322\ : Span4Mux_v
    port map (
            O => \N__24530\,
            I => \N__24515\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__24527\,
            I => \N__24515\
        );

    \I__5320\ : Span4Mux_v
    port map (
            O => \N__24520\,
            I => \N__24510\
        );

    \I__5319\ : Span4Mux_v
    port map (
            O => \N__24515\,
            I => \N__24510\
        );

    \I__5318\ : Odrv4
    port map (
            O => \N__24510\,
            I => \N_813_0\
        );

    \I__5317\ : InMux
    port map (
            O => \N__24507\,
            I => \N__24504\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__24504\,
            I => \N__24499\
        );

    \I__5315\ : InMux
    port map (
            O => \N__24503\,
            I => \N__24494\
        );

    \I__5314\ : InMux
    port map (
            O => \N__24502\,
            I => \N__24491\
        );

    \I__5313\ : Span4Mux_v
    port map (
            O => \N__24499\,
            I => \N__24484\
        );

    \I__5312\ : CascadeMux
    port map (
            O => \N__24498\,
            I => \N__24481\
        );

    \I__5311\ : CascadeMux
    port map (
            O => \N__24497\,
            I => \N__24478\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__24494\,
            I => \N__24475\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__24491\,
            I => \N__24470\
        );

    \I__5308\ : InMux
    port map (
            O => \N__24490\,
            I => \N__24467\
        );

    \I__5307\ : InMux
    port map (
            O => \N__24489\,
            I => \N__24464\
        );

    \I__5306\ : InMux
    port map (
            O => \N__24488\,
            I => \N__24459\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__24487\,
            I => \N__24455\
        );

    \I__5304\ : Span4Mux_h
    port map (
            O => \N__24484\,
            I => \N__24452\
        );

    \I__5303\ : InMux
    port map (
            O => \N__24481\,
            I => \N__24449\
        );

    \I__5302\ : InMux
    port map (
            O => \N__24478\,
            I => \N__24446\
        );

    \I__5301\ : Span4Mux_v
    port map (
            O => \N__24475\,
            I => \N__24442\
        );

    \I__5300\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24439\
        );

    \I__5299\ : CascadeMux
    port map (
            O => \N__24473\,
            I => \N__24436\
        );

    \I__5298\ : Span4Mux_h
    port map (
            O => \N__24470\,
            I => \N__24429\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__24467\,
            I => \N__24429\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__24464\,
            I => \N__24429\
        );

    \I__5295\ : InMux
    port map (
            O => \N__24463\,
            I => \N__24426\
        );

    \I__5294\ : CascadeMux
    port map (
            O => \N__24462\,
            I => \N__24423\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__24459\,
            I => \N__24420\
        );

    \I__5292\ : InMux
    port map (
            O => \N__24458\,
            I => \N__24415\
        );

    \I__5291\ : InMux
    port map (
            O => \N__24455\,
            I => \N__24415\
        );

    \I__5290\ : Span4Mux_h
    port map (
            O => \N__24452\,
            I => \N__24412\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__24449\,
            I => \N__24409\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__24446\,
            I => \N__24406\
        );

    \I__5287\ : InMux
    port map (
            O => \N__24445\,
            I => \N__24403\
        );

    \I__5286\ : Span4Mux_v
    port map (
            O => \N__24442\,
            I => \N__24398\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__24439\,
            I => \N__24398\
        );

    \I__5284\ : InMux
    port map (
            O => \N__24436\,
            I => \N__24395\
        );

    \I__5283\ : Span4Mux_v
    port map (
            O => \N__24429\,
            I => \N__24392\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__24426\,
            I => \N__24389\
        );

    \I__5281\ : InMux
    port map (
            O => \N__24423\,
            I => \N__24386\
        );

    \I__5280\ : Span4Mux_h
    port map (
            O => \N__24420\,
            I => \N__24381\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__24415\,
            I => \N__24381\
        );

    \I__5278\ : Span4Mux_h
    port map (
            O => \N__24412\,
            I => \N__24372\
        );

    \I__5277\ : Span4Mux_v
    port map (
            O => \N__24409\,
            I => \N__24372\
        );

    \I__5276\ : Span4Mux_v
    port map (
            O => \N__24406\,
            I => \N__24372\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__24403\,
            I => \N__24372\
        );

    \I__5274\ : Span4Mux_v
    port map (
            O => \N__24398\,
            I => \N__24367\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__24395\,
            I => \N__24367\
        );

    \I__5272\ : Sp12to4
    port map (
            O => \N__24392\,
            I => \N__24364\
        );

    \I__5271\ : Span12Mux_h
    port map (
            O => \N__24389\,
            I => \N__24359\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__24386\,
            I => \N__24359\
        );

    \I__5269\ : Span4Mux_v
    port map (
            O => \N__24381\,
            I => \N__24354\
        );

    \I__5268\ : Span4Mux_v
    port map (
            O => \N__24372\,
            I => \N__24354\
        );

    \I__5267\ : Span4Mux_h
    port map (
            O => \N__24367\,
            I => \N__24351\
        );

    \I__5266\ : Span12Mux_h
    port map (
            O => \N__24364\,
            I => \N__24348\
        );

    \I__5265\ : Span12Mux_h
    port map (
            O => \N__24359\,
            I => \N__24345\
        );

    \I__5264\ : Sp12to4
    port map (
            O => \N__24354\,
            I => \N__24342\
        );

    \I__5263\ : Span4Mux_h
    port map (
            O => \N__24351\,
            I => \N__24339\
        );

    \I__5262\ : Odrv12
    port map (
            O => \N__24348\,
            I => port_data_c_5
        );

    \I__5261\ : Odrv12
    port map (
            O => \N__24345\,
            I => port_data_c_5
        );

    \I__5260\ : Odrv12
    port map (
            O => \N__24342\,
            I => port_data_c_5
        );

    \I__5259\ : Odrv4
    port map (
            O => \N__24339\,
            I => port_data_c_5
        );

    \I__5258\ : CascadeMux
    port map (
            O => \N__24330\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_6_cascade_\
        );

    \I__5257\ : InMux
    port map (
            O => \N__24327\,
            I => \N__24324\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__24324\,
            I => \N__24321\
        );

    \I__5255\ : Odrv12
    port map (
            O => \N__24321\,
            I => \this_start_data_delay.N_68\
        );

    \I__5254\ : CascadeMux
    port map (
            O => \N__24318\,
            I => \N__24314\
        );

    \I__5253\ : CascadeMux
    port map (
            O => \N__24317\,
            I => \N__24310\
        );

    \I__5252\ : InMux
    port map (
            O => \N__24314\,
            I => \N__24305\
        );

    \I__5251\ : CascadeMux
    port map (
            O => \N__24313\,
            I => \N__24302\
        );

    \I__5250\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24298\
        );

    \I__5249\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24295\
        );

    \I__5248\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24292\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__24305\,
            I => \N__24289\
        );

    \I__5246\ : InMux
    port map (
            O => \N__24302\,
            I => \N__24286\
        );

    \I__5245\ : CascadeMux
    port map (
            O => \N__24301\,
            I => \N__24282\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__24298\,
            I => \N__24278\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__24295\,
            I => \N__24275\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__24292\,
            I => \N__24268\
        );

    \I__5241\ : Span4Mux_h
    port map (
            O => \N__24289\,
            I => \N__24268\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__24286\,
            I => \N__24268\
        );

    \I__5239\ : InMux
    port map (
            O => \N__24285\,
            I => \N__24265\
        );

    \I__5238\ : InMux
    port map (
            O => \N__24282\,
            I => \N__24260\
        );

    \I__5237\ : InMux
    port map (
            O => \N__24281\,
            I => \N__24260\
        );

    \I__5236\ : Span4Mux_h
    port map (
            O => \N__24278\,
            I => \N__24257\
        );

    \I__5235\ : Span4Mux_v
    port map (
            O => \N__24275\,
            I => \N__24252\
        );

    \I__5234\ : Span4Mux_h
    port map (
            O => \N__24268\,
            I => \N__24252\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__24265\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__24260\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__5231\ : Odrv4
    port map (
            O => \N__24257\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__5230\ : Odrv4
    port map (
            O => \N__24252\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__5229\ : InMux
    port map (
            O => \N__24243\,
            I => \N__24236\
        );

    \I__5228\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24232\
        );

    \I__5227\ : InMux
    port map (
            O => \N__24241\,
            I => \N__24228\
        );

    \I__5226\ : InMux
    port map (
            O => \N__24240\,
            I => \N__24218\
        );

    \I__5225\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24214\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__24236\,
            I => \N__24211\
        );

    \I__5223\ : InMux
    port map (
            O => \N__24235\,
            I => \N__24208\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__24232\,
            I => \N__24205\
        );

    \I__5221\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24201\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__24228\,
            I => \N__24198\
        );

    \I__5219\ : InMux
    port map (
            O => \N__24227\,
            I => \N__24195\
        );

    \I__5218\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24192\
        );

    \I__5217\ : InMux
    port map (
            O => \N__24225\,
            I => \N__24187\
        );

    \I__5216\ : InMux
    port map (
            O => \N__24224\,
            I => \N__24187\
        );

    \I__5215\ : InMux
    port map (
            O => \N__24223\,
            I => \N__24180\
        );

    \I__5214\ : InMux
    port map (
            O => \N__24222\,
            I => \N__24180\
        );

    \I__5213\ : InMux
    port map (
            O => \N__24221\,
            I => \N__24180\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__24218\,
            I => \N__24175\
        );

    \I__5211\ : InMux
    port map (
            O => \N__24217\,
            I => \N__24172\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__24214\,
            I => \N__24165\
        );

    \I__5209\ : Span4Mux_v
    port map (
            O => \N__24211\,
            I => \N__24165\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__24208\,
            I => \N__24165\
        );

    \I__5207\ : Span4Mux_h
    port map (
            O => \N__24205\,
            I => \N__24154\
        );

    \I__5206\ : InMux
    port map (
            O => \N__24204\,
            I => \N__24151\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__24201\,
            I => \N__24144\
        );

    \I__5204\ : Span4Mux_h
    port map (
            O => \N__24198\,
            I => \N__24144\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__24195\,
            I => \N__24144\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__24192\,
            I => \N__24141\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__24187\,
            I => \N__24136\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__24180\,
            I => \N__24136\
        );

    \I__5199\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24131\
        );

    \I__5198\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24131\
        );

    \I__5197\ : Span4Mux_v
    port map (
            O => \N__24175\,
            I => \N__24118\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__24172\,
            I => \N__24118\
        );

    \I__5195\ : Span4Mux_h
    port map (
            O => \N__24165\,
            I => \N__24118\
        );

    \I__5194\ : InMux
    port map (
            O => \N__24164\,
            I => \N__24115\
        );

    \I__5193\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24110\
        );

    \I__5192\ : InMux
    port map (
            O => \N__24162\,
            I => \N__24110\
        );

    \I__5191\ : InMux
    port map (
            O => \N__24161\,
            I => \N__24107\
        );

    \I__5190\ : InMux
    port map (
            O => \N__24160\,
            I => \N__24098\
        );

    \I__5189\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24098\
        );

    \I__5188\ : InMux
    port map (
            O => \N__24158\,
            I => \N__24098\
        );

    \I__5187\ : InMux
    port map (
            O => \N__24157\,
            I => \N__24098\
        );

    \I__5186\ : Span4Mux_h
    port map (
            O => \N__24154\,
            I => \N__24093\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__24151\,
            I => \N__24093\
        );

    \I__5184\ : Span4Mux_h
    port map (
            O => \N__24144\,
            I => \N__24084\
        );

    \I__5183\ : Span4Mux_v
    port map (
            O => \N__24141\,
            I => \N__24084\
        );

    \I__5182\ : Span4Mux_h
    port map (
            O => \N__24136\,
            I => \N__24084\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__24131\,
            I => \N__24084\
        );

    \I__5180\ : InMux
    port map (
            O => \N__24130\,
            I => \N__24077\
        );

    \I__5179\ : InMux
    port map (
            O => \N__24129\,
            I => \N__24077\
        );

    \I__5178\ : InMux
    port map (
            O => \N__24128\,
            I => \N__24077\
        );

    \I__5177\ : InMux
    port map (
            O => \N__24127\,
            I => \N__24070\
        );

    \I__5176\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24070\
        );

    \I__5175\ : InMux
    port map (
            O => \N__24125\,
            I => \N__24070\
        );

    \I__5174\ : Odrv4
    port map (
            O => \N__24118\,
            I => \N_554_0\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__24115\,
            I => \N_554_0\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__24110\,
            I => \N_554_0\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__24107\,
            I => \N_554_0\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__24098\,
            I => \N_554_0\
        );

    \I__5169\ : Odrv4
    port map (
            O => \N__24093\,
            I => \N_554_0\
        );

    \I__5168\ : Odrv4
    port map (
            O => \N__24084\,
            I => \N_554_0\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__24077\,
            I => \N_554_0\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__24070\,
            I => \N_554_0\
        );

    \I__5165\ : CascadeMux
    port map (
            O => \N__24051\,
            I => \this_start_data_delay_M_this_data_count_q_3_0_a3_0_6_cascade_\
        );

    \I__5164\ : InMux
    port map (
            O => \N__24048\,
            I => \N__24029\
        );

    \I__5163\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24029\
        );

    \I__5162\ : InMux
    port map (
            O => \N__24046\,
            I => \N__24029\
        );

    \I__5161\ : InMux
    port map (
            O => \N__24045\,
            I => \N__24029\
        );

    \I__5160\ : InMux
    port map (
            O => \N__24044\,
            I => \N__24020\
        );

    \I__5159\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24020\
        );

    \I__5158\ : InMux
    port map (
            O => \N__24042\,
            I => \N__24020\
        );

    \I__5157\ : InMux
    port map (
            O => \N__24041\,
            I => \N__24020\
        );

    \I__5156\ : InMux
    port map (
            O => \N__24040\,
            I => \N__24016\
        );

    \I__5155\ : InMux
    port map (
            O => \N__24039\,
            I => \N__24011\
        );

    \I__5154\ : InMux
    port map (
            O => \N__24038\,
            I => \N__24011\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__24029\,
            I => \N__24006\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__24020\,
            I => \N__24006\
        );

    \I__5151\ : InMux
    port map (
            O => \N__24019\,
            I => \N__24003\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__24016\,
            I => \N__24000\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__23994\
        );

    \I__5148\ : Span12Mux_v
    port map (
            O => \N__24006\,
            I => \N__23994\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__24003\,
            I => \N__23991\
        );

    \I__5146\ : Span4Mux_v
    port map (
            O => \N__24000\,
            I => \N__23988\
        );

    \I__5145\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23985\
        );

    \I__5144\ : Span12Mux_h
    port map (
            O => \N__23994\,
            I => \N__23982\
        );

    \I__5143\ : Span4Mux_h
    port map (
            O => \N__23991\,
            I => \N__23979\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__23988\,
            I => \N_911\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__23985\,
            I => \N_911\
        );

    \I__5140\ : Odrv12
    port map (
            O => \N__23982\,
            I => \N_911\
        );

    \I__5139\ : Odrv4
    port map (
            O => \N__23979\,
            I => \N_911\
        );

    \I__5138\ : InMux
    port map (
            O => \N__23970\,
            I => \N__23967\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__23967\,
            I => \N__23964\
        );

    \I__5136\ : Span4Mux_h
    port map (
            O => \N__23964\,
            I => \N__23961\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__23961\,
            I => \M_this_data_count_q_3_0_13\
        );

    \I__5134\ : InMux
    port map (
            O => \N__23958\,
            I => \N__23951\
        );

    \I__5133\ : InMux
    port map (
            O => \N__23957\,
            I => \N__23948\
        );

    \I__5132\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23942\
        );

    \I__5131\ : InMux
    port map (
            O => \N__23955\,
            I => \N__23942\
        );

    \I__5130\ : InMux
    port map (
            O => \N__23954\,
            I => \N__23939\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__23951\,
            I => \N__23936\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__23948\,
            I => \N__23933\
        );

    \I__5127\ : InMux
    port map (
            O => \N__23947\,
            I => \N__23930\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__23942\,
            I => \N__23927\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__23939\,
            I => \N__23922\
        );

    \I__5124\ : Span4Mux_h
    port map (
            O => \N__23936\,
            I => \N__23922\
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__23933\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__23930\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__23927\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5120\ : Odrv4
    port map (
            O => \N__23922\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5119\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23910\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__23910\,
            I => \N__23907\
        );

    \I__5117\ : Span4Mux_h
    port map (
            O => \N__23907\,
            I => \N__23902\
        );

    \I__5116\ : InMux
    port map (
            O => \N__23906\,
            I => \N__23896\
        );

    \I__5115\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23896\
        );

    \I__5114\ : Span4Mux_h
    port map (
            O => \N__23902\,
            I => \N__23893\
        );

    \I__5113\ : InMux
    port map (
            O => \N__23901\,
            I => \N__23890\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__23896\,
            I => \N__23886\
        );

    \I__5111\ : Sp12to4
    port map (
            O => \N__23893\,
            I => \N__23881\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__23890\,
            I => \N__23881\
        );

    \I__5109\ : InMux
    port map (
            O => \N__23889\,
            I => \N__23878\
        );

    \I__5108\ : Span4Mux_v
    port map (
            O => \N__23886\,
            I => \N__23875\
        );

    \I__5107\ : Odrv12
    port map (
            O => \N__23881\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__23878\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__5105\ : Odrv4
    port map (
            O => \N__23875\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__5104\ : CascadeMux
    port map (
            O => \N__23868\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_3_cascade_\
        );

    \I__5103\ : CascadeMux
    port map (
            O => \N__23865\,
            I => \N__23862\
        );

    \I__5102\ : InMux
    port map (
            O => \N__23862\,
            I => \N__23859\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__23859\,
            I => \N__23856\
        );

    \I__5100\ : Span4Mux_h
    port map (
            O => \N__23856\,
            I => \N__23853\
        );

    \I__5099\ : Sp12to4
    port map (
            O => \N__23853\,
            I => \N__23850\
        );

    \I__5098\ : Span12Mux_v
    port map (
            O => \N__23850\,
            I => \N__23847\
        );

    \I__5097\ : Span12Mux_h
    port map (
            O => \N__23847\,
            I => \N__23844\
        );

    \I__5096\ : Odrv12
    port map (
            O => \N__23844\,
            I => \M_this_map_ram_read_data_7\
        );

    \I__5095\ : InMux
    port map (
            O => \N__23841\,
            I => \N__23838\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__23838\,
            I => \N__23835\
        );

    \I__5093\ : Odrv12
    port map (
            O => \N__23835\,
            I => \this_ppu.un10_sprites_addr_cry_4_c_RNIUV9BZ0\
        );

    \I__5092\ : InMux
    port map (
            O => \N__23832\,
            I => \N__23829\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__23829\,
            I => \N__23824\
        );

    \I__5090\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23821\
        );

    \I__5089\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23817\
        );

    \I__5088\ : Span4Mux_v
    port map (
            O => \N__23824\,
            I => \N__23812\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__23821\,
            I => \N__23812\
        );

    \I__5086\ : InMux
    port map (
            O => \N__23820\,
            I => \N__23809\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__23817\,
            I => \this_start_data_delay.N_91_0\
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__23812\,
            I => \this_start_data_delay.N_91_0\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__23809\,
            I => \this_start_data_delay.N_91_0\
        );

    \I__5082\ : CascadeMux
    port map (
            O => \N__23802\,
            I => \this_start_data_delay.N_149_cascade_\
        );

    \I__5081\ : InMux
    port map (
            O => \N__23799\,
            I => \N__23792\
        );

    \I__5080\ : CascadeMux
    port map (
            O => \N__23798\,
            I => \N__23788\
        );

    \I__5079\ : InMux
    port map (
            O => \N__23797\,
            I => \N__23785\
        );

    \I__5078\ : InMux
    port map (
            O => \N__23796\,
            I => \N__23782\
        );

    \I__5077\ : CascadeMux
    port map (
            O => \N__23795\,
            I => \N__23777\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__23792\,
            I => \N__23773\
        );

    \I__5075\ : InMux
    port map (
            O => \N__23791\,
            I => \N__23770\
        );

    \I__5074\ : InMux
    port map (
            O => \N__23788\,
            I => \N__23767\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__23785\,
            I => \N__23762\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__23782\,
            I => \N__23762\
        );

    \I__5071\ : InMux
    port map (
            O => \N__23781\,
            I => \N__23757\
        );

    \I__5070\ : InMux
    port map (
            O => \N__23780\,
            I => \N__23757\
        );

    \I__5069\ : InMux
    port map (
            O => \N__23777\,
            I => \N__23752\
        );

    \I__5068\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23752\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__23773\,
            I => \N__23745\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__23770\,
            I => \N__23745\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__23767\,
            I => \N__23745\
        );

    \I__5064\ : Span4Mux_v
    port map (
            O => \N__23762\,
            I => \N__23740\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__23757\,
            I => \N__23740\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__23752\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__5061\ : Odrv4
    port map (
            O => \N__23745\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__23740\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__5059\ : InMux
    port map (
            O => \N__23733\,
            I => \N__23728\
        );

    \I__5058\ : InMux
    port map (
            O => \N__23732\,
            I => \N__23723\
        );

    \I__5057\ : InMux
    port map (
            O => \N__23731\,
            I => \N__23720\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__23728\,
            I => \N__23717\
        );

    \I__5055\ : InMux
    port map (
            O => \N__23727\,
            I => \N__23714\
        );

    \I__5054\ : InMux
    port map (
            O => \N__23726\,
            I => \N__23711\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__23723\,
            I => \N__23708\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__23720\,
            I => \N__23703\
        );

    \I__5051\ : Span4Mux_h
    port map (
            O => \N__23717\,
            I => \N__23703\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__23714\,
            I => \this_start_data_delay.N_555_0\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__23711\,
            I => \this_start_data_delay.N_555_0\
        );

    \I__5048\ : Odrv4
    port map (
            O => \N__23708\,
            I => \this_start_data_delay.N_555_0\
        );

    \I__5047\ : Odrv4
    port map (
            O => \N__23703\,
            I => \this_start_data_delay.N_555_0\
        );

    \I__5046\ : InMux
    port map (
            O => \N__23694\,
            I => \N__23691\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__23691\,
            I => \N__23688\
        );

    \I__5044\ : Odrv4
    port map (
            O => \N__23688\,
            I => \this_start_data_delay.M_this_data_count_qlde_i_a3_0\
        );

    \I__5043\ : InMux
    port map (
            O => \N__23685\,
            I => \N__23682\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__23682\,
            I => \this_start_data_delay.M_this_data_count_qlde_i_2_tz_0\
        );

    \I__5041\ : CascadeMux
    port map (
            O => \N__23679\,
            I => \this_start_data_delay.N_820_0_cascade_\
        );

    \I__5040\ : InMux
    port map (
            O => \N__23676\,
            I => \N__23673\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__23673\,
            I => \N__23670\
        );

    \I__5038\ : Span4Mux_h
    port map (
            O => \N__23670\,
            I => \N__23667\
        );

    \I__5037\ : Odrv4
    port map (
            O => \N__23667\,
            I => \this_start_data_delay.N_151\
        );

    \I__5036\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23660\
        );

    \I__5035\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23657\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__23660\,
            I => \N__23653\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__23657\,
            I => \N__23649\
        );

    \I__5032\ : InMux
    port map (
            O => \N__23656\,
            I => \N__23646\
        );

    \I__5031\ : Span4Mux_h
    port map (
            O => \N__23653\,
            I => \N__23643\
        );

    \I__5030\ : InMux
    port map (
            O => \N__23652\,
            I => \N__23640\
        );

    \I__5029\ : Span4Mux_v
    port map (
            O => \N__23649\,
            I => \N__23637\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__23646\,
            I => \this_start_data_delay.N_820_0\
        );

    \I__5027\ : Odrv4
    port map (
            O => \N__23643\,
            I => \this_start_data_delay.N_820_0\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__23640\,
            I => \this_start_data_delay.N_820_0\
        );

    \I__5025\ : Odrv4
    port map (
            O => \N__23637\,
            I => \this_start_data_delay.N_820_0\
        );

    \I__5024\ : CascadeMux
    port map (
            O => \N__23628\,
            I => \this_start_data_delay.M_this_data_count_qlde_i_1_cascade_\
        );

    \I__5023\ : InMux
    port map (
            O => \N__23625\,
            I => \N__23622\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__23622\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_11\
        );

    \I__5021\ : CascadeMux
    port map (
            O => \N__23619\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_10_cascade_\
        );

    \I__5020\ : InMux
    port map (
            O => \N__23616\,
            I => \N__23613\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__23613\,
            I => \N__23610\
        );

    \I__5018\ : Span4Mux_v
    port map (
            O => \N__23610\,
            I => \N__23607\
        );

    \I__5017\ : Span4Mux_v
    port map (
            O => \N__23607\,
            I => \N__23604\
        );

    \I__5016\ : Span4Mux_h
    port map (
            O => \N__23604\,
            I => \N__23601\
        );

    \I__5015\ : Odrv4
    port map (
            O => \N__23601\,
            I => \this_sprites_ram.mem_out_bus7_1\
        );

    \I__5014\ : InMux
    port map (
            O => \N__23598\,
            I => \N__23595\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__23595\,
            I => \N__23592\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__23592\,
            I => \N__23589\
        );

    \I__5011\ : Span4Mux_h
    port map (
            O => \N__23589\,
            I => \N__23586\
        );

    \I__5010\ : Odrv4
    port map (
            O => \N__23586\,
            I => \this_sprites_ram.mem_out_bus3_1\
        );

    \I__5009\ : InMux
    port map (
            O => \N__23583\,
            I => \N__23580\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__23580\,
            I => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\
        );

    \I__5007\ : CascadeMux
    port map (
            O => \N__23577\,
            I => \N__23573\
        );

    \I__5006\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23568\
        );

    \I__5005\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23565\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__23572\,
            I => \N__23562\
        );

    \I__5003\ : InMux
    port map (
            O => \N__23571\,
            I => \N__23559\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__23568\,
            I => \N__23556\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__23565\,
            I => \N__23553\
        );

    \I__5000\ : InMux
    port map (
            O => \N__23562\,
            I => \N__23550\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__23559\,
            I => \N__23547\
        );

    \I__4998\ : Span4Mux_v
    port map (
            O => \N__23556\,
            I => \N__23542\
        );

    \I__4997\ : Span4Mux_v
    port map (
            O => \N__23553\,
            I => \N__23542\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__23550\,
            I => \N__23539\
        );

    \I__4995\ : Odrv4
    port map (
            O => \N__23547\,
            I => \this_start_data_delay.N_55_0\
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__23542\,
            I => \this_start_data_delay.N_55_0\
        );

    \I__4993\ : Odrv4
    port map (
            O => \N__23539\,
            I => \this_start_data_delay.N_55_0\
        );

    \I__4992\ : InMux
    port map (
            O => \N__23532\,
            I => \N__23528\
        );

    \I__4991\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23525\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__23528\,
            I => \N__23522\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__23525\,
            I => \N__23519\
        );

    \I__4988\ : Odrv4
    port map (
            O => \N__23522\,
            I => \this_start_data_delay.N_84\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__23519\,
            I => \this_start_data_delay.N_84\
        );

    \I__4986\ : CascadeMux
    port map (
            O => \N__23514\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_2_cascade_\
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__23511\,
            I => \this_start_data_delay.N_913_cascade_\
        );

    \I__4984\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23505\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__23505\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_7\
        );

    \I__4982\ : CascadeMux
    port map (
            O => \N__23502\,
            I => \this_start_data_delay.N_129_cascade_\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__23499\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_12_cascade_\
        );

    \I__4980\ : CascadeMux
    port map (
            O => \N__23496\,
            I => \N__23492\
        );

    \I__4979\ : CascadeMux
    port map (
            O => \N__23495\,
            I => \N__23486\
        );

    \I__4978\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23483\
        );

    \I__4977\ : InMux
    port map (
            O => \N__23491\,
            I => \N__23478\
        );

    \I__4976\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23478\
        );

    \I__4975\ : InMux
    port map (
            O => \N__23489\,
            I => \N__23475\
        );

    \I__4974\ : InMux
    port map (
            O => \N__23486\,
            I => \N__23469\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__23483\,
            I => \N__23464\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__23478\,
            I => \N__23464\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__23475\,
            I => \N__23461\
        );

    \I__4970\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23458\
        );

    \I__4969\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23455\
        );

    \I__4968\ : InMux
    port map (
            O => \N__23472\,
            I => \N__23452\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__23469\,
            I => \N__23447\
        );

    \I__4966\ : Span4Mux_h
    port map (
            O => \N__23464\,
            I => \N__23447\
        );

    \I__4965\ : Odrv4
    port map (
            O => \N__23461\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__23458\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__23455\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__23452\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__4961\ : Odrv4
    port map (
            O => \N__23447\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__4960\ : CascadeMux
    port map (
            O => \N__23436\,
            I => \this_start_data_delay.N_821_0_cascade_\
        );

    \I__4959\ : InMux
    port map (
            O => \N__23433\,
            I => \N__23430\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__23430\,
            I => \N__23425\
        );

    \I__4957\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23420\
        );

    \I__4956\ : InMux
    port map (
            O => \N__23428\,
            I => \N__23420\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__23425\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__23420\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__4953\ : InMux
    port map (
            O => \N__23415\,
            I => \N__23412\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__23412\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__4951\ : CEMux
    port map (
            O => \N__23409\,
            I => \N__23403\
        );

    \I__4950\ : CEMux
    port map (
            O => \N__23408\,
            I => \N__23398\
        );

    \I__4949\ : CEMux
    port map (
            O => \N__23407\,
            I => \N__23394\
        );

    \I__4948\ : CEMux
    port map (
            O => \N__23406\,
            I => \N__23391\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__23403\,
            I => \N__23388\
        );

    \I__4946\ : CEMux
    port map (
            O => \N__23402\,
            I => \N__23385\
        );

    \I__4945\ : CEMux
    port map (
            O => \N__23401\,
            I => \N__23382\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__23398\,
            I => \N__23379\
        );

    \I__4943\ : CEMux
    port map (
            O => \N__23397\,
            I => \N__23376\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__23394\,
            I => \N__23373\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__23391\,
            I => \N__23370\
        );

    \I__4940\ : Span4Mux_h
    port map (
            O => \N__23388\,
            I => \N__23367\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__23385\,
            I => \N__23364\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__23382\,
            I => \N__23361\
        );

    \I__4937\ : Span4Mux_h
    port map (
            O => \N__23379\,
            I => \N__23355\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__23376\,
            I => \N__23355\
        );

    \I__4935\ : Span4Mux_h
    port map (
            O => \N__23373\,
            I => \N__23352\
        );

    \I__4934\ : Span4Mux_v
    port map (
            O => \N__23370\,
            I => \N__23349\
        );

    \I__4933\ : Span4Mux_v
    port map (
            O => \N__23367\,
            I => \N__23342\
        );

    \I__4932\ : Span4Mux_h
    port map (
            O => \N__23364\,
            I => \N__23342\
        );

    \I__4931\ : Span4Mux_h
    port map (
            O => \N__23361\,
            I => \N__23342\
        );

    \I__4930\ : CEMux
    port map (
            O => \N__23360\,
            I => \N__23339\
        );

    \I__4929\ : Span4Mux_h
    port map (
            O => \N__23355\,
            I => \N__23336\
        );

    \I__4928\ : Span4Mux_h
    port map (
            O => \N__23352\,
            I => \N__23333\
        );

    \I__4927\ : Sp12to4
    port map (
            O => \N__23349\,
            I => \N__23326\
        );

    \I__4926\ : Sp12to4
    port map (
            O => \N__23342\,
            I => \N__23326\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__23339\,
            I => \N__23326\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__23336\,
            I => \this_vga_signals.N_1090_0\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__23333\,
            I => \this_vga_signals.N_1090_0\
        );

    \I__4922\ : Odrv12
    port map (
            O => \N__23326\,
            I => \this_vga_signals.N_1090_0\
        );

    \I__4921\ : SRMux
    port map (
            O => \N__23319\,
            I => \N__23292\
        );

    \I__4920\ : SRMux
    port map (
            O => \N__23318\,
            I => \N__23292\
        );

    \I__4919\ : SRMux
    port map (
            O => \N__23317\,
            I => \N__23292\
        );

    \I__4918\ : SRMux
    port map (
            O => \N__23316\,
            I => \N__23292\
        );

    \I__4917\ : SRMux
    port map (
            O => \N__23315\,
            I => \N__23292\
        );

    \I__4916\ : SRMux
    port map (
            O => \N__23314\,
            I => \N__23292\
        );

    \I__4915\ : SRMux
    port map (
            O => \N__23313\,
            I => \N__23292\
        );

    \I__4914\ : SRMux
    port map (
            O => \N__23312\,
            I => \N__23292\
        );

    \I__4913\ : SRMux
    port map (
            O => \N__23311\,
            I => \N__23292\
        );

    \I__4912\ : GlobalMux
    port map (
            O => \N__23292\,
            I => \N__23289\
        );

    \I__4911\ : gio2CtrlBuf
    port map (
            O => \N__23289\,
            I => \this_vga_signals.N_1358_g\
        );

    \I__4910\ : CascadeMux
    port map (
            O => \N__23286\,
            I => \N__23279\
        );

    \I__4909\ : InMux
    port map (
            O => \N__23285\,
            I => \N__23273\
        );

    \I__4908\ : CascadeMux
    port map (
            O => \N__23284\,
            I => \N__23269\
        );

    \I__4907\ : CascadeMux
    port map (
            O => \N__23283\,
            I => \N__23263\
        );

    \I__4906\ : CascadeMux
    port map (
            O => \N__23282\,
            I => \N__23260\
        );

    \I__4905\ : InMux
    port map (
            O => \N__23279\,
            I => \N__23254\
        );

    \I__4904\ : InMux
    port map (
            O => \N__23278\,
            I => \N__23254\
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__23277\,
            I => \N__23251\
        );

    \I__4902\ : InMux
    port map (
            O => \N__23276\,
            I => \N__23245\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__23273\,
            I => \N__23242\
        );

    \I__4900\ : InMux
    port map (
            O => \N__23272\,
            I => \N__23237\
        );

    \I__4899\ : InMux
    port map (
            O => \N__23269\,
            I => \N__23237\
        );

    \I__4898\ : InMux
    port map (
            O => \N__23268\,
            I => \N__23234\
        );

    \I__4897\ : InMux
    port map (
            O => \N__23267\,
            I => \N__23229\
        );

    \I__4896\ : InMux
    port map (
            O => \N__23266\,
            I => \N__23229\
        );

    \I__4895\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23222\
        );

    \I__4894\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23222\
        );

    \I__4893\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23222\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__23254\,
            I => \N__23218\
        );

    \I__4891\ : InMux
    port map (
            O => \N__23251\,
            I => \N__23215\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__23250\,
            I => \N__23210\
        );

    \I__4889\ : CascadeMux
    port map (
            O => \N__23249\,
            I => \N__23207\
        );

    \I__4888\ : InMux
    port map (
            O => \N__23248\,
            I => \N__23204\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__23245\,
            I => \N__23194\
        );

    \I__4886\ : Span4Mux_v
    port map (
            O => \N__23242\,
            I => \N__23194\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__23237\,
            I => \N__23191\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__23234\,
            I => \N__23184\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__23229\,
            I => \N__23184\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__23222\,
            I => \N__23184\
        );

    \I__4881\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23180\
        );

    \I__4880\ : Span4Mux_v
    port map (
            O => \N__23218\,
            I => \N__23175\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__23215\,
            I => \N__23175\
        );

    \I__4878\ : InMux
    port map (
            O => \N__23214\,
            I => \N__23166\
        );

    \I__4877\ : InMux
    port map (
            O => \N__23213\,
            I => \N__23166\
        );

    \I__4876\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23166\
        );

    \I__4875\ : InMux
    port map (
            O => \N__23207\,
            I => \N__23166\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__23204\,
            I => \N__23163\
        );

    \I__4873\ : CascadeMux
    port map (
            O => \N__23203\,
            I => \N__23160\
        );

    \I__4872\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23155\
        );

    \I__4871\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23152\
        );

    \I__4870\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23147\
        );

    \I__4869\ : InMux
    port map (
            O => \N__23199\,
            I => \N__23147\
        );

    \I__4868\ : Span4Mux_v
    port map (
            O => \N__23194\,
            I => \N__23140\
        );

    \I__4867\ : Span4Mux_v
    port map (
            O => \N__23191\,
            I => \N__23140\
        );

    \I__4866\ : Span4Mux_v
    port map (
            O => \N__23184\,
            I => \N__23140\
        );

    \I__4865\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23137\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__23180\,
            I => \N__23134\
        );

    \I__4863\ : Span4Mux_h
    port map (
            O => \N__23175\,
            I => \N__23127\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__23166\,
            I => \N__23127\
        );

    \I__4861\ : Span4Mux_h
    port map (
            O => \N__23163\,
            I => \N__23127\
        );

    \I__4860\ : InMux
    port map (
            O => \N__23160\,
            I => \N__23120\
        );

    \I__4859\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23120\
        );

    \I__4858\ : InMux
    port map (
            O => \N__23158\,
            I => \N__23120\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__23155\,
            I => \N__23115\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__23152\,
            I => \N__23115\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__23147\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__4854\ : Odrv4
    port map (
            O => \N__23140\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__23137\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__4852\ : Odrv12
    port map (
            O => \N__23134\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__4851\ : Odrv4
    port map (
            O => \N__23127\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__23120\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__23115\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__23100\,
            I => \N__23094\
        );

    \I__4847\ : CascadeMux
    port map (
            O => \N__23099\,
            I => \N__23084\
        );

    \I__4846\ : CascadeMux
    port map (
            O => \N__23098\,
            I => \N__23081\
        );

    \I__4845\ : CascadeMux
    port map (
            O => \N__23097\,
            I => \N__23078\
        );

    \I__4844\ : InMux
    port map (
            O => \N__23094\,
            I => \N__23074\
        );

    \I__4843\ : CascadeMux
    port map (
            O => \N__23093\,
            I => \N__23070\
        );

    \I__4842\ : CascadeMux
    port map (
            O => \N__23092\,
            I => \N__23066\
        );

    \I__4841\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23060\
        );

    \I__4840\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23060\
        );

    \I__4839\ : InMux
    port map (
            O => \N__23089\,
            I => \N__23057\
        );

    \I__4838\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23054\
        );

    \I__4837\ : InMux
    port map (
            O => \N__23087\,
            I => \N__23051\
        );

    \I__4836\ : InMux
    port map (
            O => \N__23084\,
            I => \N__23048\
        );

    \I__4835\ : InMux
    port map (
            O => \N__23081\,
            I => \N__23045\
        );

    \I__4834\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23040\
        );

    \I__4833\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23040\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__23074\,
            I => \N__23036\
        );

    \I__4831\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23031\
        );

    \I__4830\ : InMux
    port map (
            O => \N__23070\,
            I => \N__23031\
        );

    \I__4829\ : InMux
    port map (
            O => \N__23069\,
            I => \N__23026\
        );

    \I__4828\ : InMux
    port map (
            O => \N__23066\,
            I => \N__23026\
        );

    \I__4827\ : InMux
    port map (
            O => \N__23065\,
            I => \N__23023\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__23060\,
            I => \N__23020\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__23057\,
            I => \N__23017\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__23054\,
            I => \N__23014\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__23051\,
            I => \N__23011\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__23048\,
            I => \N__23004\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__23045\,
            I => \N__23004\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__23040\,
            I => \N__23004\
        );

    \I__4819\ : CascadeMux
    port map (
            O => \N__23039\,
            I => \N__23001\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__23036\,
            I => \N__22991\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__23031\,
            I => \N__22988\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__23026\,
            I => \N__22983\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__23023\,
            I => \N__22983\
        );

    \I__4814\ : Span4Mux_h
    port map (
            O => \N__23020\,
            I => \N__22980\
        );

    \I__4813\ : Span4Mux_v
    port map (
            O => \N__23017\,
            I => \N__22971\
        );

    \I__4812\ : Span4Mux_v
    port map (
            O => \N__23014\,
            I => \N__22971\
        );

    \I__4811\ : Span4Mux_h
    port map (
            O => \N__23011\,
            I => \N__22971\
        );

    \I__4810\ : Span4Mux_v
    port map (
            O => \N__23004\,
            I => \N__22971\
        );

    \I__4809\ : InMux
    port map (
            O => \N__23001\,
            I => \N__22966\
        );

    \I__4808\ : InMux
    port map (
            O => \N__23000\,
            I => \N__22966\
        );

    \I__4807\ : InMux
    port map (
            O => \N__22999\,
            I => \N__22957\
        );

    \I__4806\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22957\
        );

    \I__4805\ : InMux
    port map (
            O => \N__22997\,
            I => \N__22957\
        );

    \I__4804\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22957\
        );

    \I__4803\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22952\
        );

    \I__4802\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22952\
        );

    \I__4801\ : Odrv4
    port map (
            O => \N__22991\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__4800\ : Odrv4
    port map (
            O => \N__22988\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__4799\ : Odrv4
    port map (
            O => \N__22983\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__22980\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__22971\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__22966\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__22957\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__22952\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__4793\ : InMux
    port map (
            O => \N__22935\,
            I => \N__22930\
        );

    \I__4792\ : InMux
    port map (
            O => \N__22934\,
            I => \N__22925\
        );

    \I__4791\ : InMux
    port map (
            O => \N__22933\,
            I => \N__22922\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__22930\,
            I => \N__22919\
        );

    \I__4789\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22916\
        );

    \I__4788\ : InMux
    port map (
            O => \N__22928\,
            I => \N__22912\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__22925\,
            I => \N__22907\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__22922\,
            I => \N__22907\
        );

    \I__4785\ : Span4Mux_v
    port map (
            O => \N__22919\,
            I => \N__22902\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__22916\,
            I => \N__22902\
        );

    \I__4783\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22899\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__22912\,
            I => \N__22895\
        );

    \I__4781\ : Span4Mux_v
    port map (
            O => \N__22907\,
            I => \N__22890\
        );

    \I__4780\ : Span4Mux_h
    port map (
            O => \N__22902\,
            I => \N__22890\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__22899\,
            I => \N__22887\
        );

    \I__4778\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22884\
        );

    \I__4777\ : Span12Mux_h
    port map (
            O => \N__22895\,
            I => \N__22881\
        );

    \I__4776\ : Span4Mux_h
    port map (
            O => \N__22890\,
            I => \N__22878\
        );

    \I__4775\ : Odrv12
    port map (
            O => \N__22887\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__22884\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__4773\ : Odrv12
    port map (
            O => \N__22881\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__4772\ : Odrv4
    port map (
            O => \N__22878\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__4771\ : CascadeMux
    port map (
            O => \N__22869\,
            I => \N__22862\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__22868\,
            I => \N__22851\
        );

    \I__4769\ : InMux
    port map (
            O => \N__22867\,
            I => \N__22844\
        );

    \I__4768\ : InMux
    port map (
            O => \N__22866\,
            I => \N__22844\
        );

    \I__4767\ : CascadeMux
    port map (
            O => \N__22865\,
            I => \N__22836\
        );

    \I__4766\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22833\
        );

    \I__4765\ : InMux
    port map (
            O => \N__22861\,
            I => \N__22830\
        );

    \I__4764\ : CascadeMux
    port map (
            O => \N__22860\,
            I => \N__22827\
        );

    \I__4763\ : InMux
    port map (
            O => \N__22859\,
            I => \N__22824\
        );

    \I__4762\ : InMux
    port map (
            O => \N__22858\,
            I => \N__22821\
        );

    \I__4761\ : InMux
    port map (
            O => \N__22857\,
            I => \N__22816\
        );

    \I__4760\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22816\
        );

    \I__4759\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22813\
        );

    \I__4758\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22808\
        );

    \I__4757\ : InMux
    port map (
            O => \N__22851\,
            I => \N__22808\
        );

    \I__4756\ : InMux
    port map (
            O => \N__22850\,
            I => \N__22803\
        );

    \I__4755\ : InMux
    port map (
            O => \N__22849\,
            I => \N__22803\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__22844\,
            I => \N__22800\
        );

    \I__4753\ : InMux
    port map (
            O => \N__22843\,
            I => \N__22797\
        );

    \I__4752\ : InMux
    port map (
            O => \N__22842\,
            I => \N__22794\
        );

    \I__4751\ : InMux
    port map (
            O => \N__22841\,
            I => \N__22791\
        );

    \I__4750\ : InMux
    port map (
            O => \N__22840\,
            I => \N__22788\
        );

    \I__4749\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22783\
        );

    \I__4748\ : InMux
    port map (
            O => \N__22836\,
            I => \N__22783\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__22833\,
            I => \N__22778\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__22830\,
            I => \N__22778\
        );

    \I__4745\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22775\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__22824\,
            I => \N__22772\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__22821\,
            I => \N__22760\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__22816\,
            I => \N__22760\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__22813\,
            I => \N__22760\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__22808\,
            I => \N__22760\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__22803\,
            I => \N__22760\
        );

    \I__4738\ : Span4Mux_h
    port map (
            O => \N__22800\,
            I => \N__22755\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__22797\,
            I => \N__22755\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__22794\,
            I => \N__22750\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__22791\,
            I => \N__22750\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__22788\,
            I => \N__22739\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__22783\,
            I => \N__22739\
        );

    \I__4732\ : Span4Mux_v
    port map (
            O => \N__22778\,
            I => \N__22739\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__22775\,
            I => \N__22739\
        );

    \I__4730\ : Span4Mux_h
    port map (
            O => \N__22772\,
            I => \N__22739\
        );

    \I__4729\ : InMux
    port map (
            O => \N__22771\,
            I => \N__22736\
        );

    \I__4728\ : Span4Mux_v
    port map (
            O => \N__22760\,
            I => \N__22733\
        );

    \I__4727\ : Span4Mux_v
    port map (
            O => \N__22755\,
            I => \N__22730\
        );

    \I__4726\ : Span4Mux_v
    port map (
            O => \N__22750\,
            I => \N__22725\
        );

    \I__4725\ : Span4Mux_h
    port map (
            O => \N__22739\,
            I => \N__22725\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__22736\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__4723\ : Odrv4
    port map (
            O => \N__22733\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__4722\ : Odrv4
    port map (
            O => \N__22730\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__4721\ : Odrv4
    port map (
            O => \N__22725\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__4720\ : CascadeMux
    port map (
            O => \N__22716\,
            I => \N__22710\
        );

    \I__4719\ : InMux
    port map (
            O => \N__22715\,
            I => \N__22697\
        );

    \I__4718\ : InMux
    port map (
            O => \N__22714\,
            I => \N__22697\
        );

    \I__4717\ : InMux
    port map (
            O => \N__22713\,
            I => \N__22694\
        );

    \I__4716\ : InMux
    port map (
            O => \N__22710\,
            I => \N__22691\
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__22709\,
            I => \N__22688\
        );

    \I__4714\ : InMux
    port map (
            O => \N__22708\,
            I => \N__22685\
        );

    \I__4713\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22682\
        );

    \I__4712\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22677\
        );

    \I__4711\ : InMux
    port map (
            O => \N__22705\,
            I => \N__22677\
        );

    \I__4710\ : InMux
    port map (
            O => \N__22704\,
            I => \N__22674\
        );

    \I__4709\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22669\
        );

    \I__4708\ : InMux
    port map (
            O => \N__22702\,
            I => \N__22666\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__22697\,
            I => \N__22659\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__22694\,
            I => \N__22659\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__22691\,
            I => \N__22659\
        );

    \I__4704\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22656\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__22685\,
            I => \N__22649\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__22682\,
            I => \N__22649\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__22677\,
            I => \N__22649\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__22674\,
            I => \N__22645\
        );

    \I__4699\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22642\
        );

    \I__4698\ : InMux
    port map (
            O => \N__22672\,
            I => \N__22639\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__22669\,
            I => \N__22636\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__22666\,
            I => \N__22633\
        );

    \I__4695\ : Span4Mux_v
    port map (
            O => \N__22659\,
            I => \N__22630\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__22656\,
            I => \N__22627\
        );

    \I__4693\ : Span4Mux_v
    port map (
            O => \N__22649\,
            I => \N__22624\
        );

    \I__4692\ : InMux
    port map (
            O => \N__22648\,
            I => \N__22621\
        );

    \I__4691\ : Span4Mux_v
    port map (
            O => \N__22645\,
            I => \N__22618\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__22642\,
            I => \N__22613\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__22639\,
            I => \N__22613\
        );

    \I__4688\ : Span4Mux_h
    port map (
            O => \N__22636\,
            I => \N__22610\
        );

    \I__4687\ : Span4Mux_h
    port map (
            O => \N__22633\,
            I => \N__22605\
        );

    \I__4686\ : Span4Mux_h
    port map (
            O => \N__22630\,
            I => \N__22605\
        );

    \I__4685\ : Span4Mux_v
    port map (
            O => \N__22627\,
            I => \N__22600\
        );

    \I__4684\ : Span4Mux_h
    port map (
            O => \N__22624\,
            I => \N__22600\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__22621\,
            I => \N__22593\
        );

    \I__4682\ : Span4Mux_h
    port map (
            O => \N__22618\,
            I => \N__22593\
        );

    \I__4681\ : Span4Mux_v
    port map (
            O => \N__22613\,
            I => \N__22593\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__22610\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__4679\ : Odrv4
    port map (
            O => \N__22605\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__4678\ : Odrv4
    port map (
            O => \N__22600\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__4677\ : Odrv4
    port map (
            O => \N__22593\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__4676\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22575\
        );

    \I__4675\ : InMux
    port map (
            O => \N__22583\,
            I => \N__22572\
        );

    \I__4674\ : InMux
    port map (
            O => \N__22582\,
            I => \N__22566\
        );

    \I__4673\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22559\
        );

    \I__4672\ : InMux
    port map (
            O => \N__22580\,
            I => \N__22559\
        );

    \I__4671\ : InMux
    port map (
            O => \N__22579\,
            I => \N__22559\
        );

    \I__4670\ : InMux
    port map (
            O => \N__22578\,
            I => \N__22556\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__22575\,
            I => \N__22551\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__22572\,
            I => \N__22551\
        );

    \I__4667\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22546\
        );

    \I__4666\ : InMux
    port map (
            O => \N__22570\,
            I => \N__22546\
        );

    \I__4665\ : InMux
    port map (
            O => \N__22569\,
            I => \N__22541\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__22566\,
            I => \N__22538\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__22559\,
            I => \N__22527\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__22556\,
            I => \N__22524\
        );

    \I__4661\ : Span4Mux_v
    port map (
            O => \N__22551\,
            I => \N__22521\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__22546\,
            I => \N__22518\
        );

    \I__4659\ : InMux
    port map (
            O => \N__22545\,
            I => \N__22513\
        );

    \I__4658\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22513\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__22541\,
            I => \N__22510\
        );

    \I__4656\ : Span4Mux_h
    port map (
            O => \N__22538\,
            I => \N__22507\
        );

    \I__4655\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22504\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__22536\,
            I => \N__22498\
        );

    \I__4653\ : CascadeMux
    port map (
            O => \N__22535\,
            I => \N__22495\
        );

    \I__4652\ : InMux
    port map (
            O => \N__22534\,
            I => \N__22492\
        );

    \I__4651\ : InMux
    port map (
            O => \N__22533\,
            I => \N__22489\
        );

    \I__4650\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22482\
        );

    \I__4649\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22482\
        );

    \I__4648\ : InMux
    port map (
            O => \N__22530\,
            I => \N__22482\
        );

    \I__4647\ : Span4Mux_h
    port map (
            O => \N__22527\,
            I => \N__22471\
        );

    \I__4646\ : Span4Mux_v
    port map (
            O => \N__22524\,
            I => \N__22471\
        );

    \I__4645\ : Span4Mux_h
    port map (
            O => \N__22521\,
            I => \N__22471\
        );

    \I__4644\ : Span4Mux_v
    port map (
            O => \N__22518\,
            I => \N__22471\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__22513\,
            I => \N__22471\
        );

    \I__4642\ : Span4Mux_v
    port map (
            O => \N__22510\,
            I => \N__22464\
        );

    \I__4641\ : Span4Mux_h
    port map (
            O => \N__22507\,
            I => \N__22464\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__22504\,
            I => \N__22464\
        );

    \I__4639\ : InMux
    port map (
            O => \N__22503\,
            I => \N__22459\
        );

    \I__4638\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22459\
        );

    \I__4637\ : InMux
    port map (
            O => \N__22501\,
            I => \N__22452\
        );

    \I__4636\ : InMux
    port map (
            O => \N__22498\,
            I => \N__22452\
        );

    \I__4635\ : InMux
    port map (
            O => \N__22495\,
            I => \N__22452\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__22492\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__22489\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__22482\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__4631\ : Odrv4
    port map (
            O => \N__22471\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__22464\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__22459\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__22452\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__4627\ : CascadeMux
    port map (
            O => \N__22437\,
            I => \N__22434\
        );

    \I__4626\ : InMux
    port map (
            O => \N__22434\,
            I => \N__22430\
        );

    \I__4625\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22427\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__22430\,
            I => \N__22424\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__22427\,
            I => \N__22421\
        );

    \I__4622\ : Span4Mux_h
    port map (
            O => \N__22424\,
            I => \N__22418\
        );

    \I__4621\ : Odrv4
    port map (
            O => \N__22421\,
            I => \this_vga_signals.m58_1\
        );

    \I__4620\ : Odrv4
    port map (
            O => \N__22418\,
            I => \this_vga_signals.m58_1\
        );

    \I__4619\ : InMux
    port map (
            O => \N__22413\,
            I => \N__22410\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__22410\,
            I => \this_vga_signals.m58_0\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__22407\,
            I => \this_vga_signals.m58_4_cascade_\
        );

    \I__4616\ : CascadeMux
    port map (
            O => \N__22404\,
            I => \N__22397\
        );

    \I__4615\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22394\
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__22402\,
            I => \N__22388\
        );

    \I__4613\ : InMux
    port map (
            O => \N__22401\,
            I => \N__22383\
        );

    \I__4612\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22380\
        );

    \I__4611\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22377\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__22394\,
            I => \N__22374\
        );

    \I__4609\ : InMux
    port map (
            O => \N__22393\,
            I => \N__22367\
        );

    \I__4608\ : InMux
    port map (
            O => \N__22392\,
            I => \N__22367\
        );

    \I__4607\ : InMux
    port map (
            O => \N__22391\,
            I => \N__22367\
        );

    \I__4606\ : InMux
    port map (
            O => \N__22388\,
            I => \N__22364\
        );

    \I__4605\ : InMux
    port map (
            O => \N__22387\,
            I => \N__22357\
        );

    \I__4604\ : InMux
    port map (
            O => \N__22386\,
            I => \N__22353\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__22383\,
            I => \N__22348\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__22380\,
            I => \N__22345\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__22377\,
            I => \N__22342\
        );

    \I__4600\ : Span4Mux_v
    port map (
            O => \N__22374\,
            I => \N__22335\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__22367\,
            I => \N__22335\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__22364\,
            I => \N__22335\
        );

    \I__4597\ : CascadeMux
    port map (
            O => \N__22363\,
            I => \N__22331\
        );

    \I__4596\ : InMux
    port map (
            O => \N__22362\,
            I => \N__22328\
        );

    \I__4595\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22324\
        );

    \I__4594\ : InMux
    port map (
            O => \N__22360\,
            I => \N__22321\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__22357\,
            I => \N__22317\
        );

    \I__4592\ : InMux
    port map (
            O => \N__22356\,
            I => \N__22313\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__22353\,
            I => \N__22310\
        );

    \I__4590\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22305\
        );

    \I__4589\ : InMux
    port map (
            O => \N__22351\,
            I => \N__22305\
        );

    \I__4588\ : Span4Mux_v
    port map (
            O => \N__22348\,
            I => \N__22296\
        );

    \I__4587\ : Span4Mux_h
    port map (
            O => \N__22345\,
            I => \N__22296\
        );

    \I__4586\ : Span4Mux_v
    port map (
            O => \N__22342\,
            I => \N__22296\
        );

    \I__4585\ : Span4Mux_v
    port map (
            O => \N__22335\,
            I => \N__22296\
        );

    \I__4584\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22291\
        );

    \I__4583\ : InMux
    port map (
            O => \N__22331\,
            I => \N__22291\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__22328\,
            I => \N__22288\
        );

    \I__4581\ : CascadeMux
    port map (
            O => \N__22327\,
            I => \N__22285\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__22324\,
            I => \N__22282\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__22321\,
            I => \N__22279\
        );

    \I__4578\ : InMux
    port map (
            O => \N__22320\,
            I => \N__22276\
        );

    \I__4577\ : Span4Mux_h
    port map (
            O => \N__22317\,
            I => \N__22273\
        );

    \I__4576\ : CascadeMux
    port map (
            O => \N__22316\,
            I => \N__22266\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__22313\,
            I => \N__22257\
        );

    \I__4574\ : Span4Mux_h
    port map (
            O => \N__22310\,
            I => \N__22257\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__22305\,
            I => \N__22257\
        );

    \I__4572\ : Span4Mux_h
    port map (
            O => \N__22296\,
            I => \N__22250\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__22291\,
            I => \N__22250\
        );

    \I__4570\ : Span4Mux_h
    port map (
            O => \N__22288\,
            I => \N__22250\
        );

    \I__4569\ : InMux
    port map (
            O => \N__22285\,
            I => \N__22247\
        );

    \I__4568\ : Span4Mux_v
    port map (
            O => \N__22282\,
            I => \N__22244\
        );

    \I__4567\ : Span4Mux_v
    port map (
            O => \N__22279\,
            I => \N__22237\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__22276\,
            I => \N__22237\
        );

    \I__4565\ : Span4Mux_v
    port map (
            O => \N__22273\,
            I => \N__22237\
        );

    \I__4564\ : InMux
    port map (
            O => \N__22272\,
            I => \N__22228\
        );

    \I__4563\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22228\
        );

    \I__4562\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22228\
        );

    \I__4561\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22228\
        );

    \I__4560\ : InMux
    port map (
            O => \N__22266\,
            I => \N__22225\
        );

    \I__4559\ : InMux
    port map (
            O => \N__22265\,
            I => \N__22220\
        );

    \I__4558\ : InMux
    port map (
            O => \N__22264\,
            I => \N__22220\
        );

    \I__4557\ : Span4Mux_v
    port map (
            O => \N__22257\,
            I => \N__22213\
        );

    \I__4556\ : Span4Mux_v
    port map (
            O => \N__22250\,
            I => \N__22213\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__22247\,
            I => \N__22213\
        );

    \I__4554\ : Odrv4
    port map (
            O => \N__22244\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__4553\ : Odrv4
    port map (
            O => \N__22237\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__22228\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__22225\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__22220\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__4549\ : Odrv4
    port map (
            O => \N__22213\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__4548\ : IoInMux
    port map (
            O => \N__22200\,
            I => \N__22197\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__22197\,
            I => \N__22194\
        );

    \I__4546\ : Span4Mux_s1_v
    port map (
            O => \N__22194\,
            I => \N__22191\
        );

    \I__4545\ : Sp12to4
    port map (
            O => \N__22191\,
            I => \N__22188\
        );

    \I__4544\ : Span12Mux_s8_h
    port map (
            O => \N__22188\,
            I => \N__22185\
        );

    \I__4543\ : Span12Mux_h
    port map (
            O => \N__22185\,
            I => \N__22182\
        );

    \I__4542\ : Odrv12
    port map (
            O => \N__22182\,
            I => this_vga_signals_vsync_1_i
        );

    \I__4541\ : InMux
    port map (
            O => \N__22179\,
            I => \N__22175\
        );

    \I__4540\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22172\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__22175\,
            I => \N__22168\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__22172\,
            I => \N__22164\
        );

    \I__4537\ : InMux
    port map (
            O => \N__22171\,
            I => \N__22160\
        );

    \I__4536\ : Span4Mux_h
    port map (
            O => \N__22168\,
            I => \N__22157\
        );

    \I__4535\ : InMux
    port map (
            O => \N__22167\,
            I => \N__22154\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__22164\,
            I => \N__22151\
        );

    \I__4533\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22148\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__22160\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__22157\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__22154\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__4529\ : Odrv4
    port map (
            O => \N__22151\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__22148\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__4527\ : CascadeMux
    port map (
            O => \N__22137\,
            I => \this_start_data_delay.N_123_cascade_\
        );

    \I__4526\ : InMux
    port map (
            O => \N__22134\,
            I => \N__22130\
        );

    \I__4525\ : InMux
    port map (
            O => \N__22133\,
            I => \N__22126\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__22130\,
            I => \N__22122\
        );

    \I__4523\ : InMux
    port map (
            O => \N__22129\,
            I => \N__22119\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__22126\,
            I => \N__22115\
        );

    \I__4521\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22112\
        );

    \I__4520\ : Span4Mux_h
    port map (
            O => \N__22122\,
            I => \N__22108\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__22119\,
            I => \N__22105\
        );

    \I__4518\ : InMux
    port map (
            O => \N__22118\,
            I => \N__22102\
        );

    \I__4517\ : Span4Mux_v
    port map (
            O => \N__22115\,
            I => \N__22097\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__22112\,
            I => \N__22097\
        );

    \I__4515\ : InMux
    port map (
            O => \N__22111\,
            I => \N__22094\
        );

    \I__4514\ : Span4Mux_v
    port map (
            O => \N__22108\,
            I => \N__22087\
        );

    \I__4513\ : Span4Mux_h
    port map (
            O => \N__22105\,
            I => \N__22087\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__22102\,
            I => \N__22084\
        );

    \I__4511\ : Span4Mux_v
    port map (
            O => \N__22097\,
            I => \N__22079\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__22094\,
            I => \N__22079\
        );

    \I__4509\ : InMux
    port map (
            O => \N__22093\,
            I => \N__22076\
        );

    \I__4508\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22073\
        );

    \I__4507\ : Span4Mux_v
    port map (
            O => \N__22087\,
            I => \N__22068\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__22084\,
            I => \N__22068\
        );

    \I__4505\ : Span4Mux_v
    port map (
            O => \N__22079\,
            I => \N__22063\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__22076\,
            I => \N__22063\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__22073\,
            I => \N__22060\
        );

    \I__4502\ : Span4Mux_v
    port map (
            O => \N__22068\,
            I => \N__22053\
        );

    \I__4501\ : Span4Mux_h
    port map (
            O => \N__22063\,
            I => \N__22053\
        );

    \I__4500\ : Span4Mux_h
    port map (
            O => \N__22060\,
            I => \N__22053\
        );

    \I__4499\ : Odrv4
    port map (
            O => \N__22053\,
            I => \N_812_0\
        );

    \I__4498\ : InMux
    port map (
            O => \N__22050\,
            I => \bfn_21_21_0_\
        );

    \I__4497\ : InMux
    port map (
            O => \N__22047\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__22044\,
            I => \N__22041\
        );

    \I__4495\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22038\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__22038\,
            I => \N__22035\
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__22035\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__4492\ : InMux
    port map (
            O => \N__22032\,
            I => \N__22023\
        );

    \I__4491\ : InMux
    port map (
            O => \N__22031\,
            I => \N__22023\
        );

    \I__4490\ : InMux
    port map (
            O => \N__22030\,
            I => \N__22023\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__22023\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__4488\ : CascadeMux
    port map (
            O => \N__22020\,
            I => \N__22017\
        );

    \I__4487\ : InMux
    port map (
            O => \N__22017\,
            I => \N__22014\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__22014\,
            I => \N__22011\
        );

    \I__4485\ : Span4Mux_v
    port map (
            O => \N__22011\,
            I => \N__22008\
        );

    \I__4484\ : Span4Mux_h
    port map (
            O => \N__22008\,
            I => \N__22005\
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__22005\,
            I => \this_vga_signals.N_4557_0\
        );

    \I__4482\ : InMux
    port map (
            O => \N__22002\,
            I => \N__21994\
        );

    \I__4481\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21994\
        );

    \I__4480\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21991\
        );

    \I__4479\ : InMux
    port map (
            O => \N__21999\,
            I => \N__21986\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__21994\,
            I => \N__21982\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__21991\,
            I => \N__21979\
        );

    \I__4476\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21974\
        );

    \I__4475\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21974\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__21986\,
            I => \N__21971\
        );

    \I__4473\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21968\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__21982\,
            I => \N__21964\
        );

    \I__4471\ : Span4Mux_v
    port map (
            O => \N__21979\,
            I => \N__21957\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__21974\,
            I => \N__21957\
        );

    \I__4469\ : Span4Mux_v
    port map (
            O => \N__21971\,
            I => \N__21952\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__21968\,
            I => \N__21952\
        );

    \I__4467\ : InMux
    port map (
            O => \N__21967\,
            I => \N__21943\
        );

    \I__4466\ : Span4Mux_h
    port map (
            O => \N__21964\,
            I => \N__21940\
        );

    \I__4465\ : InMux
    port map (
            O => \N__21963\,
            I => \N__21935\
        );

    \I__4464\ : InMux
    port map (
            O => \N__21962\,
            I => \N__21935\
        );

    \I__4463\ : Span4Mux_h
    port map (
            O => \N__21957\,
            I => \N__21930\
        );

    \I__4462\ : Span4Mux_v
    port map (
            O => \N__21952\,
            I => \N__21930\
        );

    \I__4461\ : InMux
    port map (
            O => \N__21951\,
            I => \N__21923\
        );

    \I__4460\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21923\
        );

    \I__4459\ : InMux
    port map (
            O => \N__21949\,
            I => \N__21923\
        );

    \I__4458\ : InMux
    port map (
            O => \N__21948\,
            I => \N__21916\
        );

    \I__4457\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21916\
        );

    \I__4456\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21916\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__21943\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__21940\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__21935\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__4452\ : Odrv4
    port map (
            O => \N__21930\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__21923\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__21916\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__4449\ : InMux
    port map (
            O => \N__21903\,
            I => \N__21898\
        );

    \I__4448\ : InMux
    port map (
            O => \N__21902\,
            I => \N__21894\
        );

    \I__4447\ : InMux
    port map (
            O => \N__21901\,
            I => \N__21889\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__21898\,
            I => \N__21886\
        );

    \I__4445\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21883\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__21894\,
            I => \N__21879\
        );

    \I__4443\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21874\
        );

    \I__4442\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21874\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__21889\,
            I => \N__21868\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__21886\,
            I => \N__21863\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__21883\,
            I => \N__21863\
        );

    \I__4438\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21857\
        );

    \I__4437\ : Span12Mux_s11_v
    port map (
            O => \N__21879\,
            I => \N__21852\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__21874\,
            I => \N__21852\
        );

    \I__4435\ : InMux
    port map (
            O => \N__21873\,
            I => \N__21847\
        );

    \I__4434\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21847\
        );

    \I__4433\ : InMux
    port map (
            O => \N__21871\,
            I => \N__21844\
        );

    \I__4432\ : Span4Mux_h
    port map (
            O => \N__21868\,
            I => \N__21839\
        );

    \I__4431\ : Span4Mux_h
    port map (
            O => \N__21863\,
            I => \N__21839\
        );

    \I__4430\ : InMux
    port map (
            O => \N__21862\,
            I => \N__21832\
        );

    \I__4429\ : InMux
    port map (
            O => \N__21861\,
            I => \N__21832\
        );

    \I__4428\ : InMux
    port map (
            O => \N__21860\,
            I => \N__21832\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__21857\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__4426\ : Odrv12
    port map (
            O => \N__21852\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__21847\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__21844\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__4423\ : Odrv4
    port map (
            O => \N__21839\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__21832\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__4421\ : InMux
    port map (
            O => \N__21819\,
            I => \N__21815\
        );

    \I__4420\ : CascadeMux
    port map (
            O => \N__21818\,
            I => \N__21807\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__21815\,
            I => \N__21803\
        );

    \I__4418\ : InMux
    port map (
            O => \N__21814\,
            I => \N__21800\
        );

    \I__4417\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21795\
        );

    \I__4416\ : InMux
    port map (
            O => \N__21812\,
            I => \N__21795\
        );

    \I__4415\ : InMux
    port map (
            O => \N__21811\,
            I => \N__21786\
        );

    \I__4414\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21786\
        );

    \I__4413\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21786\
        );

    \I__4412\ : InMux
    port map (
            O => \N__21806\,
            I => \N__21786\
        );

    \I__4411\ : Odrv4
    port map (
            O => \N__21803\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__21800\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__21795\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__21786\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__21777\,
            I => \N__21771\
        );

    \I__4406\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21765\
        );

    \I__4405\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21762\
        );

    \I__4404\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21759\
        );

    \I__4403\ : InMux
    port map (
            O => \N__21771\,
            I => \N__21756\
        );

    \I__4402\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21751\
        );

    \I__4401\ : InMux
    port map (
            O => \N__21769\,
            I => \N__21751\
        );

    \I__4400\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21748\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__21765\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__21762\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__21759\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__21756\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__21751\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__21748\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__4393\ : InMux
    port map (
            O => \N__21735\,
            I => \N__21729\
        );

    \I__4392\ : InMux
    port map (
            O => \N__21734\,
            I => \N__21729\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__21729\,
            I => \N__21726\
        );

    \I__4390\ : Span4Mux_h
    port map (
            O => \N__21726\,
            I => \N__21723\
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__21723\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_601\
        );

    \I__4388\ : InMux
    port map (
            O => \N__21720\,
            I => \N__21716\
        );

    \I__4387\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21712\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__21716\,
            I => \N__21709\
        );

    \I__4385\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21706\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__21712\,
            I => \N__21703\
        );

    \I__4383\ : Span4Mux_v
    port map (
            O => \N__21709\,
            I => \N__21698\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__21706\,
            I => \N__21698\
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__21703\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__21698\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__4379\ : InMux
    port map (
            O => \N__21693\,
            I => \N__21687\
        );

    \I__4378\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21680\
        );

    \I__4377\ : InMux
    port map (
            O => \N__21691\,
            I => \N__21680\
        );

    \I__4376\ : InMux
    port map (
            O => \N__21690\,
            I => \N__21680\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__21687\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__21680\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__21675\,
            I => \N__21671\
        );

    \I__4372\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21667\
        );

    \I__4371\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21664\
        );

    \I__4370\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21657\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__21667\,
            I => \N__21654\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__21664\,
            I => \N__21651\
        );

    \I__4367\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21648\
        );

    \I__4366\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21643\
        );

    \I__4365\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21643\
        );

    \I__4364\ : InMux
    port map (
            O => \N__21660\,
            I => \N__21640\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__21657\,
            I => \N__21634\
        );

    \I__4362\ : Span4Mux_v
    port map (
            O => \N__21654\,
            I => \N__21631\
        );

    \I__4361\ : Span4Mux_v
    port map (
            O => \N__21651\,
            I => \N__21628\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__21648\,
            I => \N__21623\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__21643\,
            I => \N__21623\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__21640\,
            I => \N__21619\
        );

    \I__4357\ : InMux
    port map (
            O => \N__21639\,
            I => \N__21616\
        );

    \I__4356\ : InMux
    port map (
            O => \N__21638\,
            I => \N__21613\
        );

    \I__4355\ : InMux
    port map (
            O => \N__21637\,
            I => \N__21610\
        );

    \I__4354\ : Span4Mux_h
    port map (
            O => \N__21634\,
            I => \N__21607\
        );

    \I__4353\ : Span4Mux_h
    port map (
            O => \N__21631\,
            I => \N__21602\
        );

    \I__4352\ : Span4Mux_h
    port map (
            O => \N__21628\,
            I => \N__21602\
        );

    \I__4351\ : Span4Mux_h
    port map (
            O => \N__21623\,
            I => \N__21599\
        );

    \I__4350\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21596\
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__21619\,
            I => \this_vga_signals_M_hcounter_d7_0\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__21616\,
            I => \this_vga_signals_M_hcounter_d7_0\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__21613\,
            I => \this_vga_signals_M_hcounter_d7_0\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__21610\,
            I => \this_vga_signals_M_hcounter_d7_0\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__21607\,
            I => \this_vga_signals_M_hcounter_d7_0\
        );

    \I__4344\ : Odrv4
    port map (
            O => \N__21602\,
            I => \this_vga_signals_M_hcounter_d7_0\
        );

    \I__4343\ : Odrv4
    port map (
            O => \N__21599\,
            I => \this_vga_signals_M_hcounter_d7_0\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__21596\,
            I => \this_vga_signals_M_hcounter_d7_0\
        );

    \I__4341\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21575\
        );

    \I__4340\ : InMux
    port map (
            O => \N__21578\,
            I => \N__21572\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__21575\,
            I => \N__21569\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__21572\,
            I => \N__21565\
        );

    \I__4337\ : Span4Mux_h
    port map (
            O => \N__21569\,
            I => \N__21562\
        );

    \I__4336\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21559\
        );

    \I__4335\ : Span12Mux_h
    port map (
            O => \N__21565\,
            I => \N__21556\
        );

    \I__4334\ : Span4Mux_h
    port map (
            O => \N__21562\,
            I => \N__21553\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__21559\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__4332\ : Odrv12
    port map (
            O => \N__21556\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__4331\ : Odrv4
    port map (
            O => \N__21553\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__4330\ : InMux
    port map (
            O => \N__21546\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_0\
        );

    \I__4329\ : InMux
    port map (
            O => \N__21543\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_1\
        );

    \I__4328\ : InMux
    port map (
            O => \N__21540\,
            I => \N__21531\
        );

    \I__4327\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21531\
        );

    \I__4326\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21526\
        );

    \I__4325\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21526\
        );

    \I__4324\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21518\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__21531\,
            I => \N__21515\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__21526\,
            I => \N__21512\
        );

    \I__4321\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21509\
        );

    \I__4320\ : CEMux
    port map (
            O => \N__21524\,
            I => \N__21506\
        );

    \I__4319\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21501\
        );

    \I__4318\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21501\
        );

    \I__4317\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21498\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__21518\,
            I => \N__21485\
        );

    \I__4315\ : Span4Mux_v
    port map (
            O => \N__21515\,
            I => \N__21482\
        );

    \I__4314\ : Span4Mux_v
    port map (
            O => \N__21512\,
            I => \N__21479\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__21509\,
            I => \N__21473\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__21506\,
            I => \N__21466\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__21501\,
            I => \N__21466\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__21498\,
            I => \N__21466\
        );

    \I__4309\ : InMux
    port map (
            O => \N__21497\,
            I => \N__21461\
        );

    \I__4308\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21461\
        );

    \I__4307\ : InMux
    port map (
            O => \N__21495\,
            I => \N__21458\
        );

    \I__4306\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21449\
        );

    \I__4305\ : InMux
    port map (
            O => \N__21493\,
            I => \N__21449\
        );

    \I__4304\ : InMux
    port map (
            O => \N__21492\,
            I => \N__21449\
        );

    \I__4303\ : InMux
    port map (
            O => \N__21491\,
            I => \N__21449\
        );

    \I__4302\ : InMux
    port map (
            O => \N__21490\,
            I => \N__21442\
        );

    \I__4301\ : InMux
    port map (
            O => \N__21489\,
            I => \N__21442\
        );

    \I__4300\ : InMux
    port map (
            O => \N__21488\,
            I => \N__21442\
        );

    \I__4299\ : Span4Mux_v
    port map (
            O => \N__21485\,
            I => \N__21435\
        );

    \I__4298\ : Span4Mux_h
    port map (
            O => \N__21482\,
            I => \N__21435\
        );

    \I__4297\ : Span4Mux_h
    port map (
            O => \N__21479\,
            I => \N__21435\
        );

    \I__4296\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21432\
        );

    \I__4295\ : InMux
    port map (
            O => \N__21477\,
            I => \N__21429\
        );

    \I__4294\ : InMux
    port map (
            O => \N__21476\,
            I => \N__21426\
        );

    \I__4293\ : Span4Mux_h
    port map (
            O => \N__21473\,
            I => \N__21423\
        );

    \I__4292\ : Span4Mux_v
    port map (
            O => \N__21466\,
            I => \N__21420\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__21461\,
            I => \N__21417\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__21458\,
            I => \N__21402\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__21449\,
            I => \N__21402\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__21442\,
            I => \N__21402\
        );

    \I__4287\ : Sp12to4
    port map (
            O => \N__21435\,
            I => \N__21402\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__21432\,
            I => \N__21402\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__21429\,
            I => \N__21402\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__21426\,
            I => \N__21402\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__21423\,
            I => \G_442\
        );

    \I__4282\ : Odrv4
    port map (
            O => \N__21420\,
            I => \G_442\
        );

    \I__4281\ : Odrv4
    port map (
            O => \N__21417\,
            I => \G_442\
        );

    \I__4280\ : Odrv12
    port map (
            O => \N__21402\,
            I => \G_442\
        );

    \I__4279\ : InMux
    port map (
            O => \N__21393\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_2\
        );

    \I__4278\ : InMux
    port map (
            O => \N__21390\,
            I => \N__21386\
        );

    \I__4277\ : InMux
    port map (
            O => \N__21389\,
            I => \N__21382\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__21386\,
            I => \N__21379\
        );

    \I__4275\ : InMux
    port map (
            O => \N__21385\,
            I => \N__21376\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__21382\,
            I => \N__21373\
        );

    \I__4273\ : Span4Mux_v
    port map (
            O => \N__21379\,
            I => \N__21368\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__21376\,
            I => \N__21368\
        );

    \I__4271\ : Span4Mux_h
    port map (
            O => \N__21373\,
            I => \N__21365\
        );

    \I__4270\ : Span4Mux_v
    port map (
            O => \N__21368\,
            I => \N__21362\
        );

    \I__4269\ : Odrv4
    port map (
            O => \N__21365\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__4268\ : Odrv4
    port map (
            O => \N__21362\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__4267\ : InMux
    port map (
            O => \N__21357\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3\
        );

    \I__4266\ : InMux
    port map (
            O => \N__21354\,
            I => \N__21345\
        );

    \I__4265\ : InMux
    port map (
            O => \N__21353\,
            I => \N__21345\
        );

    \I__4264\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21345\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__21345\,
            I => \N__21342\
        );

    \I__4262\ : Span4Mux_h
    port map (
            O => \N__21342\,
            I => \N__21339\
        );

    \I__4261\ : Odrv4
    port map (
            O => \N__21339\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__4260\ : InMux
    port map (
            O => \N__21336\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4\
        );

    \I__4259\ : InMux
    port map (
            O => \N__21333\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5\
        );

    \I__4258\ : InMux
    port map (
            O => \N__21330\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__21327\,
            I => \this_start_data_delay.N_91_0_cascade_\
        );

    \I__4256\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21313\
        );

    \I__4255\ : InMux
    port map (
            O => \N__21323\,
            I => \N__21313\
        );

    \I__4254\ : InMux
    port map (
            O => \N__21322\,
            I => \N__21310\
        );

    \I__4253\ : InMux
    port map (
            O => \N__21321\,
            I => \N__21307\
        );

    \I__4252\ : InMux
    port map (
            O => \N__21320\,
            I => \N__21304\
        );

    \I__4251\ : InMux
    port map (
            O => \N__21319\,
            I => \N__21299\
        );

    \I__4250\ : InMux
    port map (
            O => \N__21318\,
            I => \N__21299\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__21313\,
            I => \N__21292\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__21310\,
            I => \N__21292\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__21307\,
            I => \N__21292\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__21304\,
            I => \N__21289\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__21299\,
            I => \N__21284\
        );

    \I__4244\ : Span4Mux_v
    port map (
            O => \N__21292\,
            I => \N__21284\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__21289\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__4242\ : Odrv4
    port map (
            O => \N__21284\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__4241\ : CascadeMux
    port map (
            O => \N__21279\,
            I => \this_start_data_delay.N_110_cascade_\
        );

    \I__4240\ : CascadeMux
    port map (
            O => \N__21276\,
            I => \N__21273\
        );

    \I__4239\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21267\
        );

    \I__4238\ : InMux
    port map (
            O => \N__21272\,
            I => \N__21267\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__21267\,
            I => \N__21264\
        );

    \I__4236\ : Span4Mux_h
    port map (
            O => \N__21264\,
            I => \N__21259\
        );

    \I__4235\ : InMux
    port map (
            O => \N__21263\,
            I => \N__21254\
        );

    \I__4234\ : InMux
    port map (
            O => \N__21262\,
            I => \N__21254\
        );

    \I__4233\ : Odrv4
    port map (
            O => \N__21259\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__21254\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__4231\ : InMux
    port map (
            O => \N__21249\,
            I => \N__21246\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__21246\,
            I => \N__21243\
        );

    \I__4229\ : Span4Mux_h
    port map (
            O => \N__21243\,
            I => \N__21240\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__21240\,
            I => \this_sprites_ram.mem_out_bus5_1\
        );

    \I__4227\ : InMux
    port map (
            O => \N__21237\,
            I => \N__21234\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__21234\,
            I => \N__21231\
        );

    \I__4225\ : Span4Mux_h
    port map (
            O => \N__21231\,
            I => \N__21228\
        );

    \I__4224\ : Sp12to4
    port map (
            O => \N__21228\,
            I => \N__21225\
        );

    \I__4223\ : Span12Mux_v
    port map (
            O => \N__21225\,
            I => \N__21222\
        );

    \I__4222\ : Odrv12
    port map (
            O => \N__21222\,
            I => \this_sprites_ram.mem_out_bus1_1\
        );

    \I__4221\ : InMux
    port map (
            O => \N__21219\,
            I => \N__21216\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__21216\,
            I => \N__21213\
        );

    \I__4219\ : Span4Mux_h
    port map (
            O => \N__21213\,
            I => \N__21210\
        );

    \I__4218\ : Span4Mux_v
    port map (
            O => \N__21210\,
            I => \N__21207\
        );

    \I__4217\ : Odrv4
    port map (
            O => \N__21207\,
            I => \this_sprites_ram.mem_out_bus6_1\
        );

    \I__4216\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21201\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__21201\,
            I => \N__21198\
        );

    \I__4214\ : Span4Mux_v
    port map (
            O => \N__21198\,
            I => \N__21195\
        );

    \I__4213\ : Span4Mux_h
    port map (
            O => \N__21195\,
            I => \N__21192\
        );

    \I__4212\ : Span4Mux_v
    port map (
            O => \N__21192\,
            I => \N__21189\
        );

    \I__4211\ : Odrv4
    port map (
            O => \N__21189\,
            I => \this_sprites_ram.mem_out_bus2_1\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__21186\,
            I => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0_cascade_\
        );

    \I__4209\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21180\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__21180\,
            I => \N__21177\
        );

    \I__4207\ : Span12Mux_v
    port map (
            O => \N__21177\,
            I => \N__21174\
        );

    \I__4206\ : Odrv12
    port map (
            O => \N__21174\,
            I => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__21171\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\
        );

    \I__4204\ : InMux
    port map (
            O => \N__21168\,
            I => \N__21165\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__21165\,
            I => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\
        );

    \I__4202\ : InMux
    port map (
            O => \N__21162\,
            I => \N__21157\
        );

    \I__4201\ : InMux
    port map (
            O => \N__21161\,
            I => \N__21154\
        );

    \I__4200\ : InMux
    port map (
            O => \N__21160\,
            I => \N__21151\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__21157\,
            I => \N__21148\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__21154\,
            I => \N__21145\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__21151\,
            I => \N__21142\
        );

    \I__4196\ : Span12Mux_s8_h
    port map (
            O => \N__21148\,
            I => \N__21139\
        );

    \I__4195\ : Span4Mux_h
    port map (
            O => \N__21145\,
            I => \N__21136\
        );

    \I__4194\ : Span4Mux_h
    port map (
            O => \N__21142\,
            I => \N__21133\
        );

    \I__4193\ : Span12Mux_h
    port map (
            O => \N__21139\,
            I => \N__21130\
        );

    \I__4192\ : Span4Mux_h
    port map (
            O => \N__21136\,
            I => \N__21127\
        );

    \I__4191\ : Span4Mux_h
    port map (
            O => \N__21133\,
            I => \N__21124\
        );

    \I__4190\ : Odrv12
    port map (
            O => \N__21130\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__4189\ : Odrv4
    port map (
            O => \N__21127\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__21124\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__21117\,
            I => \N__21114\
        );

    \I__4186\ : InMux
    port map (
            O => \N__21114\,
            I => \N__21111\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__21111\,
            I => \this_start_data_delay.M_this_state_q_ns_0_i_2_0\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__21108\,
            I => \N_554_0_cascade_\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__21105\,
            I => \N__21102\
        );

    \I__4182\ : InMux
    port map (
            O => \N__21102\,
            I => \N__21094\
        );

    \I__4181\ : InMux
    port map (
            O => \N__21101\,
            I => \N__21094\
        );

    \I__4180\ : InMux
    port map (
            O => \N__21100\,
            I => \N__21090\
        );

    \I__4179\ : InMux
    port map (
            O => \N__21099\,
            I => \N__21085\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__21094\,
            I => \N__21082\
        );

    \I__4177\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21079\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__21090\,
            I => \N__21076\
        );

    \I__4175\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21073\
        );

    \I__4174\ : InMux
    port map (
            O => \N__21088\,
            I => \N__21070\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__21085\,
            I => \N__21067\
        );

    \I__4172\ : Span4Mux_v
    port map (
            O => \N__21082\,
            I => \N__21064\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__21079\,
            I => \N__21057\
        );

    \I__4170\ : Span4Mux_h
    port map (
            O => \N__21076\,
            I => \N__21057\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__21073\,
            I => \N__21057\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__21070\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4167\ : Odrv12
    port map (
            O => \N__21067\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4166\ : Odrv4
    port map (
            O => \N__21064\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__21057\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4164\ : CascadeMux
    port map (
            O => \N__21048\,
            I => \this_start_data_delay.N_109_cascade_\
        );

    \I__4163\ : InMux
    port map (
            O => \N__21045\,
            I => \N__21042\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__21042\,
            I => \N__21039\
        );

    \I__4161\ : Odrv4
    port map (
            O => \N__21039\,
            I => \this_start_data_delay.M_this_sprites_address_q_0_0_0_4\
        );

    \I__4160\ : InMux
    port map (
            O => \N__21036\,
            I => \N__21033\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__21033\,
            I => \N__21030\
        );

    \I__4158\ : Odrv12
    port map (
            O => \N__21030\,
            I => \this_delay_clk.M_pipe_qZ0Z_3\
        );

    \I__4157\ : InMux
    port map (
            O => \N__21027\,
            I => \N__21020\
        );

    \I__4156\ : InMux
    port map (
            O => \N__21026\,
            I => \N__21020\
        );

    \I__4155\ : InMux
    port map (
            O => \N__21025\,
            I => \N__21017\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__21020\,
            I => \this_start_data_delay.M_last_qZ0\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__21017\,
            I => \this_start_data_delay.M_last_qZ0\
        );

    \I__4152\ : InMux
    port map (
            O => \N__21012\,
            I => \N__21004\
        );

    \I__4151\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21004\
        );

    \I__4150\ : InMux
    port map (
            O => \N__21010\,
            I => \N__20999\
        );

    \I__4149\ : InMux
    port map (
            O => \N__21009\,
            I => \N__20999\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__21004\,
            I => \N__20994\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20994\
        );

    \I__4146\ : Span4Mux_v
    port map (
            O => \N__20994\,
            I => \N__20991\
        );

    \I__4145\ : Span4Mux_h
    port map (
            O => \N__20991\,
            I => \N__20988\
        );

    \I__4144\ : Sp12to4
    port map (
            O => \N__20988\,
            I => \N__20985\
        );

    \I__4143\ : Span12Mux_h
    port map (
            O => \N__20985\,
            I => \N__20982\
        );

    \I__4142\ : Odrv12
    port map (
            O => \N__20982\,
            I => port_enb_c
        );

    \I__4141\ : InMux
    port map (
            O => \N__20979\,
            I => \N__20971\
        );

    \I__4140\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20971\
        );

    \I__4139\ : InMux
    port map (
            O => \N__20977\,
            I => \N__20966\
        );

    \I__4138\ : InMux
    port map (
            O => \N__20976\,
            I => \N__20966\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__20971\,
            I => \M_this_delay_clk_out_0\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__20966\,
            I => \M_this_delay_clk_out_0\
        );

    \I__4135\ : InMux
    port map (
            O => \N__20961\,
            I => \N__20958\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__20958\,
            I => \this_vga_signals.vaddress_1_6\
        );

    \I__4133\ : InMux
    port map (
            O => \N__20955\,
            I => \N__20952\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__20952\,
            I => \N__20949\
        );

    \I__4131\ : Span12Mux_h
    port map (
            O => \N__20949\,
            I => \N__20946\
        );

    \I__4130\ : Span12Mux_v
    port map (
            O => \N__20946\,
            I => \N__20943\
        );

    \I__4129\ : Odrv12
    port map (
            O => \N__20943\,
            I => \this_ppu.un3_sprites_addr_cry_0_c_RNIRLAZ0Z8\
        );

    \I__4128\ : CascadeMux
    port map (
            O => \N__20940\,
            I => \N__20937\
        );

    \I__4127\ : InMux
    port map (
            O => \N__20937\,
            I => \N__20934\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__20934\,
            I => \N__20930\
        );

    \I__4125\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20927\
        );

    \I__4124\ : Span4Mux_v
    port map (
            O => \N__20930\,
            I => \N__20923\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__20927\,
            I => \N__20920\
        );

    \I__4122\ : CascadeMux
    port map (
            O => \N__20926\,
            I => \N__20917\
        );

    \I__4121\ : Span4Mux_h
    port map (
            O => \N__20923\,
            I => \N__20914\
        );

    \I__4120\ : Span12Mux_h
    port map (
            O => \N__20920\,
            I => \N__20907\
        );

    \I__4119\ : InMux
    port map (
            O => \N__20917\,
            I => \N__20904\
        );

    \I__4118\ : Span4Mux_v
    port map (
            O => \N__20914\,
            I => \N__20901\
        );

    \I__4117\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20894\
        );

    \I__4116\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20894\
        );

    \I__4115\ : InMux
    port map (
            O => \N__20911\,
            I => \N__20894\
        );

    \I__4114\ : InMux
    port map (
            O => \N__20910\,
            I => \N__20891\
        );

    \I__4113\ : Span12Mux_v
    port map (
            O => \N__20907\,
            I => \N__20886\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__20904\,
            I => \N__20886\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__20901\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__20894\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__20891\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__4108\ : Odrv12
    port map (
            O => \N__20886\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__4107\ : CascadeMux
    port map (
            O => \N__20877\,
            I => \N__20874\
        );

    \I__4106\ : CascadeBuf
    port map (
            O => \N__20874\,
            I => \N__20871\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__20871\,
            I => \N__20868\
        );

    \I__4104\ : CascadeBuf
    port map (
            O => \N__20868\,
            I => \N__20865\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__20865\,
            I => \N__20862\
        );

    \I__4102\ : CascadeBuf
    port map (
            O => \N__20862\,
            I => \N__20859\
        );

    \I__4101\ : CascadeMux
    port map (
            O => \N__20859\,
            I => \N__20856\
        );

    \I__4100\ : CascadeBuf
    port map (
            O => \N__20856\,
            I => \N__20853\
        );

    \I__4099\ : CascadeMux
    port map (
            O => \N__20853\,
            I => \N__20850\
        );

    \I__4098\ : CascadeBuf
    port map (
            O => \N__20850\,
            I => \N__20847\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__20847\,
            I => \N__20844\
        );

    \I__4096\ : CascadeBuf
    port map (
            O => \N__20844\,
            I => \N__20841\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__20841\,
            I => \N__20838\
        );

    \I__4094\ : CascadeBuf
    port map (
            O => \N__20838\,
            I => \N__20835\
        );

    \I__4093\ : CascadeMux
    port map (
            O => \N__20835\,
            I => \N__20832\
        );

    \I__4092\ : CascadeBuf
    port map (
            O => \N__20832\,
            I => \N__20829\
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__20829\,
            I => \N__20826\
        );

    \I__4090\ : CascadeBuf
    port map (
            O => \N__20826\,
            I => \N__20823\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__20823\,
            I => \N__20820\
        );

    \I__4088\ : CascadeBuf
    port map (
            O => \N__20820\,
            I => \N__20817\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__20817\,
            I => \N__20814\
        );

    \I__4086\ : CascadeBuf
    port map (
            O => \N__20814\,
            I => \N__20811\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__20811\,
            I => \N__20808\
        );

    \I__4084\ : CascadeBuf
    port map (
            O => \N__20808\,
            I => \N__20805\
        );

    \I__4083\ : CascadeMux
    port map (
            O => \N__20805\,
            I => \N__20802\
        );

    \I__4082\ : CascadeBuf
    port map (
            O => \N__20802\,
            I => \N__20799\
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__20799\,
            I => \N__20796\
        );

    \I__4080\ : CascadeBuf
    port map (
            O => \N__20796\,
            I => \N__20793\
        );

    \I__4079\ : CascadeMux
    port map (
            O => \N__20793\,
            I => \N__20790\
        );

    \I__4078\ : CascadeBuf
    port map (
            O => \N__20790\,
            I => \N__20787\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__20787\,
            I => \N__20784\
        );

    \I__4076\ : InMux
    port map (
            O => \N__20784\,
            I => \N__20781\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__20781\,
            I => \N__20778\
        );

    \I__4074\ : Odrv12
    port map (
            O => \N__20778\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__4073\ : InMux
    port map (
            O => \N__20775\,
            I => \N__20772\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__20772\,
            I => \N__20769\
        );

    \I__4071\ : Span4Mux_h
    port map (
            O => \N__20769\,
            I => \N__20766\
        );

    \I__4070\ : Span4Mux_v
    port map (
            O => \N__20766\,
            I => \N__20763\
        );

    \I__4069\ : Odrv4
    port map (
            O => \N__20763\,
            I => \this_sprites_ram.mem_out_bus4_1\
        );

    \I__4068\ : InMux
    port map (
            O => \N__20760\,
            I => \N__20757\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__20757\,
            I => \N__20754\
        );

    \I__4066\ : Span4Mux_v
    port map (
            O => \N__20754\,
            I => \N__20751\
        );

    \I__4065\ : Span4Mux_h
    port map (
            O => \N__20751\,
            I => \N__20748\
        );

    \I__4064\ : Span4Mux_v
    port map (
            O => \N__20748\,
            I => \N__20745\
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__20745\,
            I => \this_sprites_ram.mem_out_bus0_1\
        );

    \I__4062\ : InMux
    port map (
            O => \N__20742\,
            I => \N__20738\
        );

    \I__4061\ : CascadeMux
    port map (
            O => \N__20741\,
            I => \N__20735\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__20738\,
            I => \N__20732\
        );

    \I__4059\ : InMux
    port map (
            O => \N__20735\,
            I => \N__20726\
        );

    \I__4058\ : Span4Mux_h
    port map (
            O => \N__20732\,
            I => \N__20723\
        );

    \I__4057\ : InMux
    port map (
            O => \N__20731\,
            I => \N__20716\
        );

    \I__4056\ : InMux
    port map (
            O => \N__20730\,
            I => \N__20716\
        );

    \I__4055\ : InMux
    port map (
            O => \N__20729\,
            I => \N__20716\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__20726\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__20723\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__20716\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__4051\ : CascadeMux
    port map (
            O => \N__20709\,
            I => \N__20706\
        );

    \I__4050\ : InMux
    port map (
            O => \N__20706\,
            I => \N__20703\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__20703\,
            I => \this_start_data_delay.N_125\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__20700\,
            I => \this_start_data_delay.un30_0_0_cascade_\
        );

    \I__4047\ : InMux
    port map (
            O => \N__20697\,
            I => \N__20694\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__20694\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_3_x1\
        );

    \I__4045\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20688\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__20688\,
            I => \N__20684\
        );

    \I__4043\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20681\
        );

    \I__4042\ : Span4Mux_h
    port map (
            O => \N__20684\,
            I => \N__20678\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__20681\,
            I => \N__20675\
        );

    \I__4040\ : Odrv4
    port map (
            O => \N__20678\,
            I => \this_vga_signals.N_4_0\
        );

    \I__4039\ : Odrv4
    port map (
            O => \N__20675\,
            I => \this_vga_signals.N_4_0\
        );

    \I__4038\ : CascadeMux
    port map (
            O => \N__20670\,
            I => \this_vga_signals.g0_6_1_cascade_\
        );

    \I__4037\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20663\
        );

    \I__4036\ : InMux
    port map (
            O => \N__20666\,
            I => \N__20657\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__20663\,
            I => \N__20648\
        );

    \I__4034\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20645\
        );

    \I__4033\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20640\
        );

    \I__4032\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20640\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__20657\,
            I => \N__20637\
        );

    \I__4030\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20632\
        );

    \I__4029\ : InMux
    port map (
            O => \N__20655\,
            I => \N__20632\
        );

    \I__4028\ : InMux
    port map (
            O => \N__20654\,
            I => \N__20623\
        );

    \I__4027\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20623\
        );

    \I__4026\ : InMux
    port map (
            O => \N__20652\,
            I => \N__20623\
        );

    \I__4025\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20623\
        );

    \I__4024\ : Odrv4
    port map (
            O => \N__20648\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__20645\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__20640\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__4021\ : Odrv12
    port map (
            O => \N__20637\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__20632\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__20623\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__4018\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20607\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__20607\,
            I => \N__20604\
        );

    \I__4016\ : Odrv4
    port map (
            O => \N__20604\,
            I => \this_vga_signals.N_4_0_0_1\
        );

    \I__4015\ : InMux
    port map (
            O => \N__20601\,
            I => \N__20598\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__20598\,
            I => \N__20595\
        );

    \I__4013\ : Odrv4
    port map (
            O => \N__20595\,
            I => \this_vga_signals.vaddress_0_5\
        );

    \I__4012\ : CascadeMux
    port map (
            O => \N__20592\,
            I => \this_vga_signals.vaddress_0_6_cascade_\
        );

    \I__4011\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20586\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__20586\,
            I => \N__20583\
        );

    \I__4009\ : Odrv4
    port map (
            O => \N__20583\,
            I => \this_vga_signals.mult1_un47_sum_c3_0\
        );

    \I__4008\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20576\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__20579\,
            I => \N__20573\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__20576\,
            I => \N__20566\
        );

    \I__4005\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20560\
        );

    \I__4004\ : InMux
    port map (
            O => \N__20572\,
            I => \N__20560\
        );

    \I__4003\ : InMux
    port map (
            O => \N__20571\,
            I => \N__20553\
        );

    \I__4002\ : InMux
    port map (
            O => \N__20570\,
            I => \N__20553\
        );

    \I__4001\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20553\
        );

    \I__4000\ : Span4Mux_h
    port map (
            O => \N__20566\,
            I => \N__20548\
        );

    \I__3999\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20545\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__20560\,
            I => \N__20542\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__20553\,
            I => \N__20539\
        );

    \I__3996\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20536\
        );

    \I__3995\ : InMux
    port map (
            O => \N__20551\,
            I => \N__20533\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__20548\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__20545\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__20542\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__20539\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__20536\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__20533\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__3988\ : InMux
    port map (
            O => \N__20520\,
            I => \N__20515\
        );

    \I__3987\ : CascadeMux
    port map (
            O => \N__20519\,
            I => \N__20510\
        );

    \I__3986\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20505\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__20515\,
            I => \N__20499\
        );

    \I__3984\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20496\
        );

    \I__3983\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20489\
        );

    \I__3982\ : InMux
    port map (
            O => \N__20510\,
            I => \N__20489\
        );

    \I__3981\ : InMux
    port map (
            O => \N__20509\,
            I => \N__20489\
        );

    \I__3980\ : InMux
    port map (
            O => \N__20508\,
            I => \N__20486\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__20505\,
            I => \N__20483\
        );

    \I__3978\ : InMux
    port map (
            O => \N__20504\,
            I => \N__20478\
        );

    \I__3977\ : InMux
    port map (
            O => \N__20503\,
            I => \N__20478\
        );

    \I__3976\ : InMux
    port map (
            O => \N__20502\,
            I => \N__20475\
        );

    \I__3975\ : Span4Mux_h
    port map (
            O => \N__20499\,
            I => \N__20466\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__20496\,
            I => \N__20466\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__20489\,
            I => \N__20466\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__20486\,
            I => \N__20466\
        );

    \I__3971\ : Odrv12
    port map (
            O => \N__20483\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__20478\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__20475\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__3968\ : Odrv4
    port map (
            O => \N__20466\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__3967\ : CascadeMux
    port map (
            O => \N__20457\,
            I => \N__20451\
        );

    \I__3966\ : CascadeMux
    port map (
            O => \N__20456\,
            I => \N__20447\
        );

    \I__3965\ : CascadeMux
    port map (
            O => \N__20455\,
            I => \N__20444\
        );

    \I__3964\ : InMux
    port map (
            O => \N__20454\,
            I => \N__20439\
        );

    \I__3963\ : InMux
    port map (
            O => \N__20451\,
            I => \N__20439\
        );

    \I__3962\ : InMux
    port map (
            O => \N__20450\,
            I => \N__20436\
        );

    \I__3961\ : InMux
    port map (
            O => \N__20447\,
            I => \N__20431\
        );

    \I__3960\ : InMux
    port map (
            O => \N__20444\,
            I => \N__20431\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__20439\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__20436\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__20431\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__3956\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20420\
        );

    \I__3955\ : InMux
    port map (
            O => \N__20423\,
            I => \N__20415\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__20420\,
            I => \N__20406\
        );

    \I__3953\ : InMux
    port map (
            O => \N__20419\,
            I => \N__20401\
        );

    \I__3952\ : InMux
    port map (
            O => \N__20418\,
            I => \N__20401\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__20415\,
            I => \N__20398\
        );

    \I__3950\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20393\
        );

    \I__3949\ : InMux
    port map (
            O => \N__20413\,
            I => \N__20393\
        );

    \I__3948\ : InMux
    port map (
            O => \N__20412\,
            I => \N__20384\
        );

    \I__3947\ : InMux
    port map (
            O => \N__20411\,
            I => \N__20384\
        );

    \I__3946\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20384\
        );

    \I__3945\ : InMux
    port map (
            O => \N__20409\,
            I => \N__20384\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__20406\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__20401\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__3942\ : Odrv4
    port map (
            O => \N__20398\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__20393\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__20384\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__3939\ : CascadeMux
    port map (
            O => \N__20373\,
            I => \N__20367\
        );

    \I__3938\ : InMux
    port map (
            O => \N__20372\,
            I => \N__20363\
        );

    \I__3937\ : InMux
    port map (
            O => \N__20371\,
            I => \N__20360\
        );

    \I__3936\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20355\
        );

    \I__3935\ : InMux
    port map (
            O => \N__20367\,
            I => \N__20355\
        );

    \I__3934\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20352\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__20363\,
            I => \N__20348\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__20360\,
            I => \N__20343\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__20355\,
            I => \N__20343\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__20352\,
            I => \N__20338\
        );

    \I__3929\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20335\
        );

    \I__3928\ : Span4Mux_v
    port map (
            O => \N__20348\,
            I => \N__20328\
        );

    \I__3927\ : Span4Mux_v
    port map (
            O => \N__20343\,
            I => \N__20328\
        );

    \I__3926\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20323\
        );

    \I__3925\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20323\
        );

    \I__3924\ : Span4Mux_h
    port map (
            O => \N__20338\,
            I => \N__20320\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__20335\,
            I => \N__20317\
        );

    \I__3922\ : InMux
    port map (
            O => \N__20334\,
            I => \N__20312\
        );

    \I__3921\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20312\
        );

    \I__3920\ : Odrv4
    port map (
            O => \N__20328\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__20323\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__20320\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__20317\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__20312\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__3915\ : CascadeMux
    port map (
            O => \N__20301\,
            I => \this_vga_signals.g2_1_cascade_\
        );

    \I__3914\ : InMux
    port map (
            O => \N__20298\,
            I => \N__20294\
        );

    \I__3913\ : InMux
    port map (
            O => \N__20297\,
            I => \N__20291\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__20294\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_2\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__20291\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_2\
        );

    \I__3910\ : InMux
    port map (
            O => \N__20286\,
            I => \N__20283\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__20283\,
            I => \N__20280\
        );

    \I__3908\ : Span4Mux_h
    port map (
            O => \N__20280\,
            I => \N__20277\
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__20277\,
            I => \this_vga_signals.g0_i_x4_0_0\
        );

    \I__3906\ : CascadeMux
    port map (
            O => \N__20274\,
            I => \N__20271\
        );

    \I__3905\ : InMux
    port map (
            O => \N__20271\,
            I => \N__20268\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__20268\,
            I => \N__20265\
        );

    \I__3903\ : Odrv12
    port map (
            O => \N__20265\,
            I => \this_vga_signals.g0_3_0_a3_1\
        );

    \I__3902\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20259\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__20259\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_602_x0\
        );

    \I__3900\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20252\
        );

    \I__3899\ : InMux
    port map (
            O => \N__20255\,
            I => \N__20249\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__20252\,
            I => \N__20240\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__20249\,
            I => \N__20240\
        );

    \I__3896\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20234\
        );

    \I__3895\ : CascadeMux
    port map (
            O => \N__20247\,
            I => \N__20230\
        );

    \I__3894\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20227\
        );

    \I__3893\ : InMux
    port map (
            O => \N__20245\,
            I => \N__20224\
        );

    \I__3892\ : Span4Mux_v
    port map (
            O => \N__20240\,
            I => \N__20221\
        );

    \I__3891\ : InMux
    port map (
            O => \N__20239\,
            I => \N__20216\
        );

    \I__3890\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20216\
        );

    \I__3889\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20213\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__20234\,
            I => \N__20210\
        );

    \I__3887\ : InMux
    port map (
            O => \N__20233\,
            I => \N__20205\
        );

    \I__3886\ : InMux
    port map (
            O => \N__20230\,
            I => \N__20205\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__20227\,
            I => \N__20202\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__20224\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__3883\ : Odrv4
    port map (
            O => \N__20221\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__20216\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__20213\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__20210\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__20205\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__20202\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__20187\,
            I => \N__20184\
        );

    \I__3876\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20180\
        );

    \I__3875\ : CascadeMux
    port map (
            O => \N__20183\,
            I => \N__20177\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__20180\,
            I => \N__20174\
        );

    \I__3873\ : InMux
    port map (
            O => \N__20177\,
            I => \N__20171\
        );

    \I__3872\ : Span4Mux_v
    port map (
            O => \N__20174\,
            I => \N__20168\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__20171\,
            I => \N__20165\
        );

    \I__3870\ : Span4Mux_h
    port map (
            O => \N__20168\,
            I => \N__20162\
        );

    \I__3869\ : Span4Mux_v
    port map (
            O => \N__20165\,
            I => \N__20159\
        );

    \I__3868\ : Odrv4
    port map (
            O => \N__20162\,
            I => \this_vga_signals.r_N_4_mux\
        );

    \I__3867\ : Odrv4
    port map (
            O => \N__20159\,
            I => \this_vga_signals.r_N_4_mux\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__20154\,
            I => \this_vga_signals.r_N_4_mux_cascade_\
        );

    \I__3865\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20148\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__20148\,
            I => \N__20144\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__20147\,
            I => \N__20141\
        );

    \I__3862\ : Span4Mux_v
    port map (
            O => \N__20144\,
            I => \N__20138\
        );

    \I__3861\ : InMux
    port map (
            O => \N__20141\,
            I => \N__20135\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__20138\,
            I => \this_vga_signals.SUM_2\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__20135\,
            I => \this_vga_signals.SUM_2\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__20130\,
            I => \N__20127\
        );

    \I__3857\ : InMux
    port map (
            O => \N__20127\,
            I => \N__20121\
        );

    \I__3856\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20118\
        );

    \I__3855\ : InMux
    port map (
            O => \N__20125\,
            I => \N__20113\
        );

    \I__3854\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20113\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__20121\,
            I => \N__20110\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__20118\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__20113\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__3850\ : Odrv4
    port map (
            O => \N__20110\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__3849\ : CascadeMux
    port map (
            O => \N__20103\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a1_x1_cascade_\
        );

    \I__3848\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20097\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__20097\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a1_ns\
        );

    \I__3846\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20091\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__20091\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a1_x0\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__20088\,
            I => \N__20080\
        );

    \I__3843\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20077\
        );

    \I__3842\ : CascadeMux
    port map (
            O => \N__20086\,
            I => \N__20074\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__20085\,
            I => \N__20067\
        );

    \I__3840\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20064\
        );

    \I__3839\ : InMux
    port map (
            O => \N__20083\,
            I => \N__20059\
        );

    \I__3838\ : InMux
    port map (
            O => \N__20080\,
            I => \N__20059\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__20077\,
            I => \N__20056\
        );

    \I__3836\ : InMux
    port map (
            O => \N__20074\,
            I => \N__20049\
        );

    \I__3835\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20049\
        );

    \I__3834\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20049\
        );

    \I__3833\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20044\
        );

    \I__3832\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20044\
        );

    \I__3831\ : InMux
    port map (
            O => \N__20067\,
            I => \N__20041\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__20064\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__20059\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__3828\ : Odrv4
    port map (
            O => \N__20056\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__20049\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__20044\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__20041\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__3824\ : InMux
    port map (
            O => \N__20028\,
            I => \N__20022\
        );

    \I__3823\ : InMux
    port map (
            O => \N__20027\,
            I => \N__20015\
        );

    \I__3822\ : InMux
    port map (
            O => \N__20026\,
            I => \N__20015\
        );

    \I__3821\ : InMux
    port map (
            O => \N__20025\,
            I => \N__20015\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__20022\,
            I => \N__20012\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__20015\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__3818\ : Odrv4
    port map (
            O => \N__20012\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__3817\ : CascadeMux
    port map (
            O => \N__20007\,
            I => \N__20004\
        );

    \I__3816\ : InMux
    port map (
            O => \N__20004\,
            I => \N__20001\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__20001\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_602_x1\
        );

    \I__3814\ : InMux
    port map (
            O => \N__19998\,
            I => \N__19995\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__19995\,
            I => \this_start_data_delay.N_67\
        );

    \I__3812\ : InMux
    port map (
            O => \N__19992\,
            I => \N__19989\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__19989\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_2_1_0\
        );

    \I__3810\ : InMux
    port map (
            O => \N__19986\,
            I => \N__19983\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__19983\,
            I => \this_vga_signals.N_4558_0\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__19980\,
            I => \this_vga_signals.g0_4_i_a3_1_cascade_\
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__19977\,
            I => \this_vga_signals.g0_4_i_1_cascade_\
        );

    \I__3806\ : InMux
    port map (
            O => \N__19974\,
            I => \N__19971\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__19971\,
            I => \this_vga_signals.N_6_2\
        );

    \I__3804\ : InMux
    port map (
            O => \N__19968\,
            I => \N__19964\
        );

    \I__3803\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19961\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__19964\,
            I => \this_start_data_delay.N_47_0\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__19961\,
            I => \this_start_data_delay.N_47_0\
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__19956\,
            I => \this_start_data_delay.N_909_0_cascade_\
        );

    \I__3799\ : IoInMux
    port map (
            O => \N__19953\,
            I => \N__19950\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__19950\,
            I => \N__19947\
        );

    \I__3797\ : IoSpan4Mux
    port map (
            O => \N__19947\,
            I => \N__19944\
        );

    \I__3796\ : Span4Mux_s0_h
    port map (
            O => \N__19944\,
            I => \N__19941\
        );

    \I__3795\ : Span4Mux_v
    port map (
            O => \N__19941\,
            I => \N__19938\
        );

    \I__3794\ : Sp12to4
    port map (
            O => \N__19938\,
            I => \N__19935\
        );

    \I__3793\ : Span12Mux_h
    port map (
            O => \N__19935\,
            I => \N__19929\
        );

    \I__3792\ : InMux
    port map (
            O => \N__19934\,
            I => \N__19926\
        );

    \I__3791\ : InMux
    port map (
            O => \N__19933\,
            I => \N__19921\
        );

    \I__3790\ : InMux
    port map (
            O => \N__19932\,
            I => \N__19921\
        );

    \I__3789\ : Odrv12
    port map (
            O => \N__19929\,
            I => led_c_1
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__19926\,
            I => led_c_1
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__19921\,
            I => led_c_1
        );

    \I__3786\ : InMux
    port map (
            O => \N__19914\,
            I => \N__19911\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__19911\,
            I => \N__19908\
        );

    \I__3784\ : Odrv4
    port map (
            O => \N__19908\,
            I => \this_start_data_delay.M_this_state_q_ns_0_i_0_0\
        );

    \I__3783\ : InMux
    port map (
            O => \N__19905\,
            I => \N__19902\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__19902\,
            I => \this_start_data_delay.M_this_state_q_ns_0_i_2_0_0\
        );

    \I__3781\ : CEMux
    port map (
            O => \N__19899\,
            I => \N__19893\
        );

    \I__3780\ : CEMux
    port map (
            O => \N__19898\,
            I => \N__19888\
        );

    \I__3779\ : InMux
    port map (
            O => \N__19897\,
            I => \N__19884\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__19896\,
            I => \N__19880\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__19893\,
            I => \N__19877\
        );

    \I__3776\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19873\
        );

    \I__3775\ : InMux
    port map (
            O => \N__19891\,
            I => \N__19869\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__19888\,
            I => \N__19865\
        );

    \I__3773\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19862\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__19884\,
            I => \N__19859\
        );

    \I__3771\ : InMux
    port map (
            O => \N__19883\,
            I => \N__19856\
        );

    \I__3770\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19853\
        );

    \I__3769\ : Span4Mux_h
    port map (
            O => \N__19877\,
            I => \N__19850\
        );

    \I__3768\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19847\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__19873\,
            I => \N__19844\
        );

    \I__3766\ : InMux
    port map (
            O => \N__19872\,
            I => \N__19841\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__19869\,
            I => \N__19838\
        );

    \I__3764\ : InMux
    port map (
            O => \N__19868\,
            I => \N__19835\
        );

    \I__3763\ : Span4Mux_h
    port map (
            O => \N__19865\,
            I => \N__19824\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__19862\,
            I => \N__19824\
        );

    \I__3761\ : Span4Mux_v
    port map (
            O => \N__19859\,
            I => \N__19824\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__19856\,
            I => \N__19824\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__19853\,
            I => \N__19824\
        );

    \I__3758\ : Span4Mux_v
    port map (
            O => \N__19850\,
            I => \N__19818\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__19847\,
            I => \N__19818\
        );

    \I__3756\ : Span4Mux_h
    port map (
            O => \N__19844\,
            I => \N__19813\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__19841\,
            I => \N__19813\
        );

    \I__3754\ : Span4Mux_h
    port map (
            O => \N__19838\,
            I => \N__19806\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__19835\,
            I => \N__19806\
        );

    \I__3752\ : Span4Mux_v
    port map (
            O => \N__19824\,
            I => \N__19806\
        );

    \I__3751\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19803\
        );

    \I__3750\ : Span4Mux_h
    port map (
            O => \N__19818\,
            I => \N__19800\
        );

    \I__3749\ : Span4Mux_v
    port map (
            O => \N__19813\,
            I => \N__19795\
        );

    \I__3748\ : Span4Mux_h
    port map (
            O => \N__19806\,
            I => \N__19795\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__19803\,
            I => \N__19791\
        );

    \I__3746\ : Span4Mux_h
    port map (
            O => \N__19800\,
            I => \N__19788\
        );

    \I__3745\ : Span4Mux_h
    port map (
            O => \N__19795\,
            I => \N__19785\
        );

    \I__3744\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19782\
        );

    \I__3743\ : Span12Mux_h
    port map (
            O => \N__19791\,
            I => \N__19777\
        );

    \I__3742\ : Sp12to4
    port map (
            O => \N__19788\,
            I => \N__19777\
        );

    \I__3741\ : Span4Mux_v
    port map (
            O => \N__19785\,
            I => \N__19774\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__19782\,
            I => \N_822_0\
        );

    \I__3739\ : Odrv12
    port map (
            O => \N__19777\,
            I => \N_822_0\
        );

    \I__3738\ : Odrv4
    port map (
            O => \N__19774\,
            I => \N_822_0\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__19767\,
            I => \this_start_data_delay.N_910_cascade_\
        );

    \I__3736\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19760\
        );

    \I__3735\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19757\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__19760\,
            I => \N__19749\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__19757\,
            I => \N__19749\
        );

    \I__3732\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19746\
        );

    \I__3731\ : InMux
    port map (
            O => \N__19755\,
            I => \N__19743\
        );

    \I__3730\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19740\
        );

    \I__3729\ : Odrv4
    port map (
            O => \N__19749\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__19746\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__19743\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__19740\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__19731\,
            I => \N__19728\
        );

    \I__3724\ : InMux
    port map (
            O => \N__19728\,
            I => \N__19724\
        );

    \I__3723\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19720\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__19724\,
            I => \N__19717\
        );

    \I__3721\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19714\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__19720\,
            I => \this_start_data_delay.N_90_0\
        );

    \I__3719\ : Odrv4
    port map (
            O => \N__19717\,
            I => \this_start_data_delay.N_90_0\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__19714\,
            I => \this_start_data_delay.N_90_0\
        );

    \I__3717\ : CascadeMux
    port map (
            O => \N__19707\,
            I => \N__19700\
        );

    \I__3716\ : CascadeMux
    port map (
            O => \N__19706\,
            I => \N__19697\
        );

    \I__3715\ : CascadeMux
    port map (
            O => \N__19705\,
            I => \N__19693\
        );

    \I__3714\ : InMux
    port map (
            O => \N__19704\,
            I => \N__19688\
        );

    \I__3713\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19688\
        );

    \I__3712\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19681\
        );

    \I__3711\ : InMux
    port map (
            O => \N__19697\,
            I => \N__19681\
        );

    \I__3710\ : InMux
    port map (
            O => \N__19696\,
            I => \N__19678\
        );

    \I__3709\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19675\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__19688\,
            I => \N__19672\
        );

    \I__3707\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19667\
        );

    \I__3706\ : InMux
    port map (
            O => \N__19686\,
            I => \N__19667\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__19681\,
            I => \N__19662\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__19678\,
            I => \N__19662\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__19675\,
            I => \N__19655\
        );

    \I__3702\ : Span4Mux_v
    port map (
            O => \N__19672\,
            I => \N__19655\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__19667\,
            I => \N__19655\
        );

    \I__3700\ : Span4Mux_v
    port map (
            O => \N__19662\,
            I => \N__19652\
        );

    \I__3699\ : Span4Mux_h
    port map (
            O => \N__19655\,
            I => \N__19649\
        );

    \I__3698\ : Span4Mux_v
    port map (
            O => \N__19652\,
            I => \N__19646\
        );

    \I__3697\ : Span4Mux_h
    port map (
            O => \N__19649\,
            I => \N__19643\
        );

    \I__3696\ : Sp12to4
    port map (
            O => \N__19646\,
            I => \N__19640\
        );

    \I__3695\ : Sp12to4
    port map (
            O => \N__19643\,
            I => \N__19637\
        );

    \I__3694\ : Span12Mux_h
    port map (
            O => \N__19640\,
            I => \N__19634\
        );

    \I__3693\ : Odrv12
    port map (
            O => \N__19637\,
            I => port_address_in_1
        );

    \I__3692\ : Odrv12
    port map (
            O => \N__19634\,
            I => port_address_in_1
        );

    \I__3691\ : InMux
    port map (
            O => \N__19629\,
            I => \N__19621\
        );

    \I__3690\ : InMux
    port map (
            O => \N__19628\,
            I => \N__19616\
        );

    \I__3689\ : InMux
    port map (
            O => \N__19627\,
            I => \N__19611\
        );

    \I__3688\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19611\
        );

    \I__3687\ : InMux
    port map (
            O => \N__19625\,
            I => \N__19606\
        );

    \I__3686\ : InMux
    port map (
            O => \N__19624\,
            I => \N__19606\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__19621\,
            I => \N__19603\
        );

    \I__3684\ : InMux
    port map (
            O => \N__19620\,
            I => \N__19598\
        );

    \I__3683\ : InMux
    port map (
            O => \N__19619\,
            I => \N__19598\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__19616\,
            I => \N__19593\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__19611\,
            I => \N__19593\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__19606\,
            I => \N__19586\
        );

    \I__3679\ : Span4Mux_v
    port map (
            O => \N__19603\,
            I => \N__19586\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__19598\,
            I => \N__19586\
        );

    \I__3677\ : Span4Mux_v
    port map (
            O => \N__19593\,
            I => \N__19583\
        );

    \I__3676\ : Span4Mux_h
    port map (
            O => \N__19586\,
            I => \N__19580\
        );

    \I__3675\ : Sp12to4
    port map (
            O => \N__19583\,
            I => \N__19577\
        );

    \I__3674\ : Sp12to4
    port map (
            O => \N__19580\,
            I => \N__19572\
        );

    \I__3673\ : Span12Mux_h
    port map (
            O => \N__19577\,
            I => \N__19572\
        );

    \I__3672\ : Odrv12
    port map (
            O => \N__19572\,
            I => port_address_in_0
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__19569\,
            I => \N__19564\
        );

    \I__3670\ : CascadeMux
    port map (
            O => \N__19568\,
            I => \N__19561\
        );

    \I__3669\ : CascadeMux
    port map (
            O => \N__19567\,
            I => \N__19556\
        );

    \I__3668\ : InMux
    port map (
            O => \N__19564\,
            I => \N__19551\
        );

    \I__3667\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19551\
        );

    \I__3666\ : InMux
    port map (
            O => \N__19560\,
            I => \N__19544\
        );

    \I__3665\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19544\
        );

    \I__3664\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19541\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__19551\,
            I => \N__19538\
        );

    \I__3662\ : InMux
    port map (
            O => \N__19550\,
            I => \N__19533\
        );

    \I__3661\ : InMux
    port map (
            O => \N__19549\,
            I => \N__19533\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__19544\,
            I => \N__19530\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__19541\,
            I => \N__19527\
        );

    \I__3658\ : Span4Mux_v
    port map (
            O => \N__19538\,
            I => \N__19522\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__19533\,
            I => \N__19522\
        );

    \I__3656\ : Span4Mux_v
    port map (
            O => \N__19530\,
            I => \N__19519\
        );

    \I__3655\ : Span4Mux_v
    port map (
            O => \N__19527\,
            I => \N__19516\
        );

    \I__3654\ : Span4Mux_h
    port map (
            O => \N__19522\,
            I => \N__19513\
        );

    \I__3653\ : Span4Mux_v
    port map (
            O => \N__19519\,
            I => \N__19508\
        );

    \I__3652\ : Span4Mux_v
    port map (
            O => \N__19516\,
            I => \N__19508\
        );

    \I__3651\ : Sp12to4
    port map (
            O => \N__19513\,
            I => \N__19505\
        );

    \I__3650\ : Span4Mux_v
    port map (
            O => \N__19508\,
            I => \N__19502\
        );

    \I__3649\ : Span12Mux_v
    port map (
            O => \N__19505\,
            I => \N__19499\
        );

    \I__3648\ : IoSpan4Mux
    port map (
            O => \N__19502\,
            I => \N__19496\
        );

    \I__3647\ : Odrv12
    port map (
            O => \N__19499\,
            I => port_address_in_2
        );

    \I__3646\ : Odrv4
    port map (
            O => \N__19496\,
            I => port_address_in_2
        );

    \I__3645\ : InMux
    port map (
            O => \N__19491\,
            I => \N__19483\
        );

    \I__3644\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19483\
        );

    \I__3643\ : InMux
    port map (
            O => \N__19489\,
            I => \N__19480\
        );

    \I__3642\ : InMux
    port map (
            O => \N__19488\,
            I => \N__19477\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__19483\,
            I => \this_start_data_delay.N_48_0\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__19480\,
            I => \this_start_data_delay.N_48_0\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__19477\,
            I => \this_start_data_delay.N_48_0\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__19470\,
            I => \N__19467\
        );

    \I__3637\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19464\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__19464\,
            I => \this_start_data_delay.N_71\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__19461\,
            I => \this_start_data_delay.N_127_cascade_\
        );

    \I__3634\ : InMux
    port map (
            O => \N__19458\,
            I => \N__19452\
        );

    \I__3633\ : InMux
    port map (
            O => \N__19457\,
            I => \N__19449\
        );

    \I__3632\ : InMux
    port map (
            O => \N__19456\,
            I => \N__19444\
        );

    \I__3631\ : InMux
    port map (
            O => \N__19455\,
            I => \N__19444\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__19452\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__19449\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__19444\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__19437\,
            I => \this_start_data_delay.N_844_0_cascade_\
        );

    \I__3626\ : CascadeMux
    port map (
            O => \N__19434\,
            I => \this_start_data_delay.N_151_cascade_\
        );

    \I__3625\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19428\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__19428\,
            I => \N__19424\
        );

    \I__3623\ : InMux
    port map (
            O => \N__19427\,
            I => \N__19419\
        );

    \I__3622\ : Span4Mux_v
    port map (
            O => \N__19424\,
            I => \N__19416\
        );

    \I__3621\ : InMux
    port map (
            O => \N__19423\,
            I => \N__19411\
        );

    \I__3620\ : InMux
    port map (
            O => \N__19422\,
            I => \N__19411\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__19419\,
            I => \this_start_data_delay.N_89_0\
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__19416\,
            I => \this_start_data_delay.N_89_0\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__19411\,
            I => \this_start_data_delay.N_89_0\
        );

    \I__3616\ : InMux
    port map (
            O => \N__19404\,
            I => \N__19400\
        );

    \I__3615\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19396\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__19400\,
            I => \N__19391\
        );

    \I__3613\ : InMux
    port map (
            O => \N__19399\,
            I => \N__19387\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__19396\,
            I => \N__19384\
        );

    \I__3611\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19381\
        );

    \I__3610\ : InMux
    port map (
            O => \N__19394\,
            I => \N__19378\
        );

    \I__3609\ : Span4Mux_v
    port map (
            O => \N__19391\,
            I => \N__19375\
        );

    \I__3608\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19372\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__19387\,
            I => \N__19369\
        );

    \I__3606\ : Span4Mux_h
    port map (
            O => \N__19384\,
            I => \N__19364\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__19381\,
            I => \N__19364\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__19378\,
            I => \M_this_state_qZ0Z_16\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__19375\,
            I => \M_this_state_qZ0Z_16\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__19372\,
            I => \M_this_state_qZ0Z_16\
        );

    \I__3601\ : Odrv4
    port map (
            O => \N__19369\,
            I => \M_this_state_qZ0Z_16\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__19364\,
            I => \M_this_state_qZ0Z_16\
        );

    \I__3599\ : InMux
    port map (
            O => \N__19353\,
            I => \N__19350\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__19350\,
            I => \N__19347\
        );

    \I__3597\ : Span4Mux_v
    port map (
            O => \N__19347\,
            I => \N__19344\
        );

    \I__3596\ : Sp12to4
    port map (
            O => \N__19344\,
            I => \N__19341\
        );

    \I__3595\ : Span12Mux_h
    port map (
            O => \N__19341\,
            I => \N__19338\
        );

    \I__3594\ : Odrv12
    port map (
            O => \N__19338\,
            I => \this_ppu.un3_sprites_addr_axb_0\
        );

    \I__3593\ : CascadeMux
    port map (
            O => \N__19335\,
            I => \N__19331\
        );

    \I__3592\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19328\
        );

    \I__3591\ : InMux
    port map (
            O => \N__19331\,
            I => \N__19325\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__19328\,
            I => \N__19322\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__19325\,
            I => \N__19319\
        );

    \I__3588\ : Span4Mux_h
    port map (
            O => \N__19322\,
            I => \N__19315\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__19319\,
            I => \N__19312\
        );

    \I__3586\ : CascadeMux
    port map (
            O => \N__19318\,
            I => \N__19308\
        );

    \I__3585\ : Span4Mux_v
    port map (
            O => \N__19315\,
            I => \N__19303\
        );

    \I__3584\ : Span4Mux_v
    port map (
            O => \N__19312\,
            I => \N__19300\
        );

    \I__3583\ : InMux
    port map (
            O => \N__19311\,
            I => \N__19297\
        );

    \I__3582\ : InMux
    port map (
            O => \N__19308\,
            I => \N__19294\
        );

    \I__3581\ : CascadeMux
    port map (
            O => \N__19307\,
            I => \N__19291\
        );

    \I__3580\ : CascadeMux
    port map (
            O => \N__19306\,
            I => \N__19287\
        );

    \I__3579\ : Span4Mux_v
    port map (
            O => \N__19303\,
            I => \N__19282\
        );

    \I__3578\ : Span4Mux_v
    port map (
            O => \N__19300\,
            I => \N__19275\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__19297\,
            I => \N__19275\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__19294\,
            I => \N__19275\
        );

    \I__3575\ : InMux
    port map (
            O => \N__19291\,
            I => \N__19266\
        );

    \I__3574\ : InMux
    port map (
            O => \N__19290\,
            I => \N__19266\
        );

    \I__3573\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19266\
        );

    \I__3572\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19266\
        );

    \I__3571\ : InMux
    port map (
            O => \N__19285\,
            I => \N__19263\
        );

    \I__3570\ : Span4Mux_v
    port map (
            O => \N__19282\,
            I => \N__19258\
        );

    \I__3569\ : Span4Mux_h
    port map (
            O => \N__19275\,
            I => \N__19258\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__19266\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__19263\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__19258\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__3565\ : CascadeMux
    port map (
            O => \N__19251\,
            I => \N__19248\
        );

    \I__3564\ : CascadeBuf
    port map (
            O => \N__19248\,
            I => \N__19245\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__19245\,
            I => \N__19242\
        );

    \I__3562\ : CascadeBuf
    port map (
            O => \N__19242\,
            I => \N__19239\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__19239\,
            I => \N__19236\
        );

    \I__3560\ : CascadeBuf
    port map (
            O => \N__19236\,
            I => \N__19233\
        );

    \I__3559\ : CascadeMux
    port map (
            O => \N__19233\,
            I => \N__19230\
        );

    \I__3558\ : CascadeBuf
    port map (
            O => \N__19230\,
            I => \N__19227\
        );

    \I__3557\ : CascadeMux
    port map (
            O => \N__19227\,
            I => \N__19224\
        );

    \I__3556\ : CascadeBuf
    port map (
            O => \N__19224\,
            I => \N__19221\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__19221\,
            I => \N__19218\
        );

    \I__3554\ : CascadeBuf
    port map (
            O => \N__19218\,
            I => \N__19215\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__19215\,
            I => \N__19212\
        );

    \I__3552\ : CascadeBuf
    port map (
            O => \N__19212\,
            I => \N__19209\
        );

    \I__3551\ : CascadeMux
    port map (
            O => \N__19209\,
            I => \N__19206\
        );

    \I__3550\ : CascadeBuf
    port map (
            O => \N__19206\,
            I => \N__19203\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__19203\,
            I => \N__19200\
        );

    \I__3548\ : CascadeBuf
    port map (
            O => \N__19200\,
            I => \N__19197\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__19197\,
            I => \N__19194\
        );

    \I__3546\ : CascadeBuf
    port map (
            O => \N__19194\,
            I => \N__19191\
        );

    \I__3545\ : CascadeMux
    port map (
            O => \N__19191\,
            I => \N__19188\
        );

    \I__3544\ : CascadeBuf
    port map (
            O => \N__19188\,
            I => \N__19185\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__19185\,
            I => \N__19182\
        );

    \I__3542\ : CascadeBuf
    port map (
            O => \N__19182\,
            I => \N__19179\
        );

    \I__3541\ : CascadeMux
    port map (
            O => \N__19179\,
            I => \N__19176\
        );

    \I__3540\ : CascadeBuf
    port map (
            O => \N__19176\,
            I => \N__19173\
        );

    \I__3539\ : CascadeMux
    port map (
            O => \N__19173\,
            I => \N__19170\
        );

    \I__3538\ : CascadeBuf
    port map (
            O => \N__19170\,
            I => \N__19167\
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__19167\,
            I => \N__19164\
        );

    \I__3536\ : CascadeBuf
    port map (
            O => \N__19164\,
            I => \N__19161\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__19161\,
            I => \N__19158\
        );

    \I__3534\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19155\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__19155\,
            I => \N__19152\
        );

    \I__3532\ : Span4Mux_h
    port map (
            O => \N__19152\,
            I => \N__19149\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__19149\,
            I => \M_this_ppu_sprites_addr_0\
        );

    \I__3530\ : InMux
    port map (
            O => \N__19146\,
            I => \N__19141\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__19145\,
            I => \N__19138\
        );

    \I__3528\ : InMux
    port map (
            O => \N__19144\,
            I => \N__19134\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__19141\,
            I => \N__19131\
        );

    \I__3526\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19126\
        );

    \I__3525\ : InMux
    port map (
            O => \N__19137\,
            I => \N__19126\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__19134\,
            I => \M_this_state_qZ0Z_15\
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__19131\,
            I => \M_this_state_qZ0Z_15\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__19126\,
            I => \M_this_state_qZ0Z_15\
        );

    \I__3521\ : InMux
    port map (
            O => \N__19119\,
            I => \N__19116\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__19116\,
            I => \N__19112\
        );

    \I__3519\ : InMux
    port map (
            O => \N__19115\,
            I => \N__19107\
        );

    \I__3518\ : Span4Mux_h
    port map (
            O => \N__19112\,
            I => \N__19104\
        );

    \I__3517\ : InMux
    port map (
            O => \N__19111\,
            I => \N__19099\
        );

    \I__3516\ : InMux
    port map (
            O => \N__19110\,
            I => \N__19099\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__19107\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__3514\ : Odrv4
    port map (
            O => \N__19104\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__19099\,
            I => \M_this_state_qZ0Z_14\
        );

    \I__3512\ : InMux
    port map (
            O => \N__19092\,
            I => \N__19088\
        );

    \I__3511\ : InMux
    port map (
            O => \N__19091\,
            I => \N__19083\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__19088\,
            I => \N__19080\
        );

    \I__3509\ : InMux
    port map (
            O => \N__19087\,
            I => \N__19075\
        );

    \I__3508\ : InMux
    port map (
            O => \N__19086\,
            I => \N__19075\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__19083\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__19080\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__19075\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__3504\ : InMux
    port map (
            O => \N__19068\,
            I => \N__19065\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__19065\,
            I => \N__19062\
        );

    \I__3502\ : Odrv4
    port map (
            O => \N__19062\,
            I => \this_start_data_delay.N_112_0\
        );

    \I__3501\ : InMux
    port map (
            O => \N__19059\,
            I => \N__19053\
        );

    \I__3500\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19053\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__19053\,
            I => \this_start_data_delay.N_80_0\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__19050\,
            I => \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_aZ0Z2_cascade_\
        );

    \I__3497\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19043\
        );

    \I__3496\ : InMux
    port map (
            O => \N__19046\,
            I => \N__19040\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__19043\,
            I => \N__19037\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__19040\,
            I => \N__19034\
        );

    \I__3493\ : Span4Mux_h
    port map (
            O => \N__19037\,
            I => \N__19031\
        );

    \I__3492\ : Span4Mux_h
    port map (
            O => \N__19034\,
            I => \N__19028\
        );

    \I__3491\ : Odrv4
    port map (
            O => \N__19031\,
            I => \this_start_data_delay.N_76_1\
        );

    \I__3490\ : Odrv4
    port map (
            O => \N__19028\,
            I => \this_start_data_delay.N_76_1\
        );

    \I__3489\ : InMux
    port map (
            O => \N__19023\,
            I => \N__19020\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__19020\,
            I => \this_vga_signals.mult1_un54_sum_ac0_4_x1\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__19017\,
            I => \this_vga_signals.mult1_un47_sum_c3_cascade_\
        );

    \I__3486\ : InMux
    port map (
            O => \N__19014\,
            I => \N__19011\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__19011\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1\
        );

    \I__3484\ : InMux
    port map (
            O => \N__19008\,
            I => \N__19005\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__19005\,
            I => \N__19001\
        );

    \I__3482\ : InMux
    port map (
            O => \N__19004\,
            I => \N__18997\
        );

    \I__3481\ : Span4Mux_h
    port map (
            O => \N__19001\,
            I => \N__18994\
        );

    \I__3480\ : InMux
    port map (
            O => \N__19000\,
            I => \N__18991\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__18997\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__18994\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__18991\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__3476\ : InMux
    port map (
            O => \N__18984\,
            I => \N__18981\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__18981\,
            I => \this_vga_signals.i1_mux\
        );

    \I__3474\ : InMux
    port map (
            O => \N__18978\,
            I => \N__18974\
        );

    \I__3473\ : InMux
    port map (
            O => \N__18977\,
            I => \N__18971\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__18974\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1_0\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__18971\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1_0\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__18966\,
            I => \N__18963\
        );

    \I__3469\ : InMux
    port map (
            O => \N__18963\,
            I => \N__18954\
        );

    \I__3468\ : InMux
    port map (
            O => \N__18962\,
            I => \N__18954\
        );

    \I__3467\ : InMux
    port map (
            O => \N__18961\,
            I => \N__18954\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__18954\,
            I => \N__18948\
        );

    \I__3465\ : InMux
    port map (
            O => \N__18953\,
            I => \N__18941\
        );

    \I__3464\ : InMux
    port map (
            O => \N__18952\,
            I => \N__18941\
        );

    \I__3463\ : InMux
    port map (
            O => \N__18951\,
            I => \N__18941\
        );

    \I__3462\ : Span4Mux_h
    port map (
            O => \N__18948\,
            I => \N__18936\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__18941\,
            I => \N__18936\
        );

    \I__3460\ : Odrv4
    port map (
            O => \N__18936\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__18933\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1_0_cascade_\
        );

    \I__3458\ : InMux
    port map (
            O => \N__18930\,
            I => \N__18927\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__18927\,
            I => \this_vga_signals.mult1_un54_sum_ac0_4_x0\
        );

    \I__3456\ : InMux
    port map (
            O => \N__18924\,
            I => \N__18921\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__18921\,
            I => \N__18917\
        );

    \I__3454\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18914\
        );

    \I__3453\ : Odrv4
    port map (
            O => \N__18917\,
            I => \this_vga_signals.g1_7\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__18914\,
            I => \this_vga_signals.g1_7\
        );

    \I__3451\ : CascadeMux
    port map (
            O => \N__18909\,
            I => \N__18906\
        );

    \I__3450\ : InMux
    port map (
            O => \N__18906\,
            I => \N__18903\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__18903\,
            I => \N__18900\
        );

    \I__3448\ : Odrv4
    port map (
            O => \N__18900\,
            I => \this_vga_signals.vaddress_3_6\
        );

    \I__3447\ : InMux
    port map (
            O => \N__18897\,
            I => \N__18894\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__18894\,
            I => \N__18891\
        );

    \I__3445\ : Span4Mux_h
    port map (
            O => \N__18891\,
            I => \N__18888\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__18888\,
            I => \this_vga_signals.g2_1_0\
        );

    \I__3443\ : InMux
    port map (
            O => \N__18885\,
            I => \N__18879\
        );

    \I__3442\ : InMux
    port map (
            O => \N__18884\,
            I => \N__18874\
        );

    \I__3441\ : InMux
    port map (
            O => \N__18883\,
            I => \N__18874\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__18882\,
            I => \N__18871\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__18879\,
            I => \N__18868\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__18874\,
            I => \N__18865\
        );

    \I__3437\ : InMux
    port map (
            O => \N__18871\,
            I => \N__18862\
        );

    \I__3436\ : Odrv12
    port map (
            O => \N__18868\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0\
        );

    \I__3435\ : Odrv4
    port map (
            O => \N__18865\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__18862\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__18855\,
            I => \N__18851\
        );

    \I__3432\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18846\
        );

    \I__3431\ : InMux
    port map (
            O => \N__18851\,
            I => \N__18846\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__18846\,
            I => \N__18843\
        );

    \I__3429\ : Odrv4
    port map (
            O => \N__18843\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_2_1\
        );

    \I__3428\ : InMux
    port map (
            O => \N__18840\,
            I => \N__18834\
        );

    \I__3427\ : InMux
    port map (
            O => \N__18839\,
            I => \N__18834\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__18834\,
            I => \N__18831\
        );

    \I__3425\ : Odrv4
    port map (
            O => \N__18831\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_a4\
        );

    \I__3424\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18825\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__18825\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_1\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__18822\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_3_cascade_\
        );

    \I__3421\ : InMux
    port map (
            O => \N__18819\,
            I => \N__18810\
        );

    \I__3420\ : InMux
    port map (
            O => \N__18818\,
            I => \N__18810\
        );

    \I__3419\ : InMux
    port map (
            O => \N__18817\,
            I => \N__18810\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__18810\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_602_ns\
        );

    \I__3417\ : CascadeMux
    port map (
            O => \N__18807\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\
        );

    \I__3416\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18801\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__18801\,
            I => \this_vga_signals.g0_1_0\
        );

    \I__3414\ : InMux
    port map (
            O => \N__18798\,
            I => \N__18794\
        );

    \I__3413\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18791\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__18794\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__18791\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__3410\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18778\
        );

    \I__3409\ : InMux
    port map (
            O => \N__18785\,
            I => \N__18773\
        );

    \I__3408\ : InMux
    port map (
            O => \N__18784\,
            I => \N__18769\
        );

    \I__3407\ : InMux
    port map (
            O => \N__18783\,
            I => \N__18755\
        );

    \I__3406\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18755\
        );

    \I__3405\ : InMux
    port map (
            O => \N__18781\,
            I => \N__18755\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__18778\,
            I => \N__18752\
        );

    \I__3403\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18747\
        );

    \I__3402\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18747\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__18773\,
            I => \N__18744\
        );

    \I__3400\ : InMux
    port map (
            O => \N__18772\,
            I => \N__18741\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__18769\,
            I => \N__18738\
        );

    \I__3398\ : InMux
    port map (
            O => \N__18768\,
            I => \N__18731\
        );

    \I__3397\ : InMux
    port map (
            O => \N__18767\,
            I => \N__18731\
        );

    \I__3396\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18731\
        );

    \I__3395\ : InMux
    port map (
            O => \N__18765\,
            I => \N__18726\
        );

    \I__3394\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18726\
        );

    \I__3393\ : InMux
    port map (
            O => \N__18763\,
            I => \N__18721\
        );

    \I__3392\ : InMux
    port map (
            O => \N__18762\,
            I => \N__18721\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__18755\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__3390\ : Odrv4
    port map (
            O => \N__18752\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__18747\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__3388\ : Odrv4
    port map (
            O => \N__18744\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__18741\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__18738\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__18731\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__18726\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__18721\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__3382\ : InMux
    port map (
            O => \N__18702\,
            I => \N__18699\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__18699\,
            I => \N__18696\
        );

    \I__3380\ : Span4Mux_h
    port map (
            O => \N__18696\,
            I => \N__18693\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__18693\,
            I => \this_vga_signals.g0_5_2_0\
        );

    \I__3378\ : InMux
    port map (
            O => \N__18690\,
            I => \N__18687\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__18687\,
            I => \N_28_0\
        );

    \I__3376\ : InMux
    port map (
            O => \N__18684\,
            I => \N__18681\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__18681\,
            I => \this_start_data_delay.N_82\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__18678\,
            I => \this_start_data_delay.N_82_cascade_\
        );

    \I__3373\ : InMux
    port map (
            O => \N__18675\,
            I => \N__18670\
        );

    \I__3372\ : InMux
    port map (
            O => \N__18674\,
            I => \N__18665\
        );

    \I__3371\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18665\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__18670\,
            I => \M_this_substate_qZ0\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__18665\,
            I => \M_this_substate_qZ0\
        );

    \I__3368\ : InMux
    port map (
            O => \N__18660\,
            I => \N__18657\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__18657\,
            I => \N__18654\
        );

    \I__3366\ : Span4Mux_v
    port map (
            O => \N__18654\,
            I => \N__18651\
        );

    \I__3365\ : Odrv4
    port map (
            O => \N__18651\,
            I => \this_vga_signals.g0_0_x4_0_0\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__18648\,
            I => \this_vga_signals.vaddress_c2_cascade_\
        );

    \I__3363\ : CascadeMux
    port map (
            O => \N__18645\,
            I => \this_vga_signals.N_5_2_1_cascade_\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__18642\,
            I => \this_vga_signals.g0_5_0_cascade_\
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__18639\,
            I => \this_vga_signals.g0_1_1_cascade_\
        );

    \I__3360\ : InMux
    port map (
            O => \N__18636\,
            I => \N__18633\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__18633\,
            I => \N__18630\
        );

    \I__3358\ : Span4Mux_v
    port map (
            O => \N__18630\,
            I => \N__18627\
        );

    \I__3357\ : Odrv4
    port map (
            O => \N__18627\,
            I => \this_vga_signals.N_3_2\
        );

    \I__3356\ : CascadeMux
    port map (
            O => \N__18624\,
            I => \N__18614\
        );

    \I__3355\ : InMux
    port map (
            O => \N__18623\,
            I => \N__18611\
        );

    \I__3354\ : CEMux
    port map (
            O => \N__18622\,
            I => \N__18605\
        );

    \I__3353\ : CEMux
    port map (
            O => \N__18621\,
            I => \N__18602\
        );

    \I__3352\ : InMux
    port map (
            O => \N__18620\,
            I => \N__18593\
        );

    \I__3351\ : InMux
    port map (
            O => \N__18619\,
            I => \N__18572\
        );

    \I__3350\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18567\
        );

    \I__3349\ : InMux
    port map (
            O => \N__18617\,
            I => \N__18567\
        );

    \I__3348\ : InMux
    port map (
            O => \N__18614\,
            I => \N__18564\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__18611\,
            I => \N__18561\
        );

    \I__3346\ : InMux
    port map (
            O => \N__18610\,
            I => \N__18554\
        );

    \I__3345\ : InMux
    port map (
            O => \N__18609\,
            I => \N__18554\
        );

    \I__3344\ : InMux
    port map (
            O => \N__18608\,
            I => \N__18554\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__18605\,
            I => \N__18549\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__18602\,
            I => \N__18549\
        );

    \I__3341\ : InMux
    port map (
            O => \N__18601\,
            I => \N__18536\
        );

    \I__3340\ : InMux
    port map (
            O => \N__18600\,
            I => \N__18536\
        );

    \I__3339\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18536\
        );

    \I__3338\ : InMux
    port map (
            O => \N__18598\,
            I => \N__18536\
        );

    \I__3337\ : InMux
    port map (
            O => \N__18597\,
            I => \N__18536\
        );

    \I__3336\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18536\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__18593\,
            I => \N__18533\
        );

    \I__3334\ : InMux
    port map (
            O => \N__18592\,
            I => \N__18528\
        );

    \I__3333\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18528\
        );

    \I__3332\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18518\
        );

    \I__3331\ : InMux
    port map (
            O => \N__18589\,
            I => \N__18518\
        );

    \I__3330\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18518\
        );

    \I__3329\ : InMux
    port map (
            O => \N__18587\,
            I => \N__18518\
        );

    \I__3328\ : InMux
    port map (
            O => \N__18586\,
            I => \N__18509\
        );

    \I__3327\ : InMux
    port map (
            O => \N__18585\,
            I => \N__18509\
        );

    \I__3326\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18509\
        );

    \I__3325\ : InMux
    port map (
            O => \N__18583\,
            I => \N__18509\
        );

    \I__3324\ : InMux
    port map (
            O => \N__18582\,
            I => \N__18496\
        );

    \I__3323\ : InMux
    port map (
            O => \N__18581\,
            I => \N__18496\
        );

    \I__3322\ : InMux
    port map (
            O => \N__18580\,
            I => \N__18496\
        );

    \I__3321\ : InMux
    port map (
            O => \N__18579\,
            I => \N__18496\
        );

    \I__3320\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18496\
        );

    \I__3319\ : InMux
    port map (
            O => \N__18577\,
            I => \N__18496\
        );

    \I__3318\ : InMux
    port map (
            O => \N__18576\,
            I => \N__18491\
        );

    \I__3317\ : InMux
    port map (
            O => \N__18575\,
            I => \N__18491\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__18572\,
            I => \N__18484\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__18567\,
            I => \N__18484\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__18564\,
            I => \N__18484\
        );

    \I__3313\ : Span4Mux_v
    port map (
            O => \N__18561\,
            I => \N__18477\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__18554\,
            I => \N__18477\
        );

    \I__3311\ : Span4Mux_v
    port map (
            O => \N__18549\,
            I => \N__18472\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__18536\,
            I => \N__18472\
        );

    \I__3309\ : Span4Mux_v
    port map (
            O => \N__18533\,
            I => \N__18467\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__18528\,
            I => \N__18467\
        );

    \I__3307\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18464\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__18518\,
            I => \N__18457\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__18509\,
            I => \N__18457\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__18496\,
            I => \N__18457\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__18491\,
            I => \N__18452\
        );

    \I__3302\ : Span4Mux_v
    port map (
            O => \N__18484\,
            I => \N__18452\
        );

    \I__3301\ : InMux
    port map (
            O => \N__18483\,
            I => \N__18449\
        );

    \I__3300\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18446\
        );

    \I__3299\ : Span4Mux_v
    port map (
            O => \N__18477\,
            I => \N__18443\
        );

    \I__3298\ : Span4Mux_h
    port map (
            O => \N__18472\,
            I => \N__18440\
        );

    \I__3297\ : Span4Mux_h
    port map (
            O => \N__18467\,
            I => \N__18437\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__18464\,
            I => \N__18434\
        );

    \I__3295\ : Span4Mux_v
    port map (
            O => \N__18457\,
            I => \N__18429\
        );

    \I__3294\ : Span4Mux_h
    port map (
            O => \N__18452\,
            I => \N__18429\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__18449\,
            I => \N__18424\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__18446\,
            I => \N__18424\
        );

    \I__3291\ : Span4Mux_h
    port map (
            O => \N__18443\,
            I => \N__18421\
        );

    \I__3290\ : Span4Mux_h
    port map (
            O => \N__18440\,
            I => \N__18418\
        );

    \I__3289\ : Span4Mux_h
    port map (
            O => \N__18437\,
            I => \N__18415\
        );

    \I__3288\ : Span4Mux_v
    port map (
            O => \N__18434\,
            I => \N__18408\
        );

    \I__3287\ : Span4Mux_h
    port map (
            O => \N__18429\,
            I => \N__18408\
        );

    \I__3286\ : Span4Mux_v
    port map (
            O => \N__18424\,
            I => \N__18408\
        );

    \I__3285\ : Odrv4
    port map (
            O => \N__18421\,
            I => led23
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__18418\,
            I => led23
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__18415\,
            I => led23
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__18408\,
            I => led23
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__18399\,
            I => \N__18396\
        );

    \I__3280\ : InMux
    port map (
            O => \N__18396\,
            I => \N__18393\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__18393\,
            I => \N__18390\
        );

    \I__3278\ : Odrv4
    port map (
            O => \N__18390\,
            I => \this_start_data_delay.dmalto4_0_a2Z0Z_1\
        );

    \I__3277\ : InMux
    port map (
            O => \N__18387\,
            I => \N__18384\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__18384\,
            I => \this_start_data_delay.N_115\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__18381\,
            I => \N__18378\
        );

    \I__3274\ : InMux
    port map (
            O => \N__18378\,
            I => \N__18375\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__18375\,
            I => \this_start_data_delay.N_69\
        );

    \I__3272\ : InMux
    port map (
            O => \N__18372\,
            I => \N__18369\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__18369\,
            I => \N__18366\
        );

    \I__3270\ : Span4Mux_v
    port map (
            O => \N__18366\,
            I => \N__18363\
        );

    \I__3269\ : Sp12to4
    port map (
            O => \N__18363\,
            I => \N__18360\
        );

    \I__3268\ : Span12Mux_h
    port map (
            O => \N__18360\,
            I => \N__18357\
        );

    \I__3267\ : Odrv12
    port map (
            O => \N__18357\,
            I => port_address_in_5
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__18354\,
            I => \N__18351\
        );

    \I__3265\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18348\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__18348\,
            I => \N__18345\
        );

    \I__3263\ : Sp12to4
    port map (
            O => \N__18345\,
            I => \N__18342\
        );

    \I__3262\ : Span12Mux_v
    port map (
            O => \N__18342\,
            I => \N__18339\
        );

    \I__3261\ : Span12Mux_h
    port map (
            O => \N__18339\,
            I => \N__18336\
        );

    \I__3260\ : Odrv12
    port map (
            O => \N__18336\,
            I => port_address_in_6
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__18333\,
            I => \this_start_data_delay.N_47_0_cascade_\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__18330\,
            I => \this_start_data_delay.N_48_0_cascade_\
        );

    \I__3257\ : CascadeMux
    port map (
            O => \N__18327\,
            I => \this_vga_signals.mult1_un54_sum_axb1_cascade_\
        );

    \I__3256\ : InMux
    port map (
            O => \N__18324\,
            I => \N__18320\
        );

    \I__3255\ : InMux
    port map (
            O => \N__18323\,
            I => \N__18317\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__18320\,
            I => \N__18313\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__18317\,
            I => \N__18310\
        );

    \I__3252\ : InMux
    port map (
            O => \N__18316\,
            I => \N__18307\
        );

    \I__3251\ : Span4Mux_v
    port map (
            O => \N__18313\,
            I => \N__18304\
        );

    \I__3250\ : Odrv4
    port map (
            O => \N__18310\,
            I => \this_vga_signals.if_N_9_i\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__18307\,
            I => \this_vga_signals.if_N_9_i\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__18304\,
            I => \this_vga_signals.if_N_9_i\
        );

    \I__3247\ : InMux
    port map (
            O => \N__18297\,
            I => \N__18294\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__18294\,
            I => \N__18289\
        );

    \I__3245\ : InMux
    port map (
            O => \N__18293\,
            I => \N__18286\
        );

    \I__3244\ : InMux
    port map (
            O => \N__18292\,
            I => \N__18283\
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__18289\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__18286\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__18283\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__3240\ : InMux
    port map (
            O => \N__18276\,
            I => \N__18273\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__18273\,
            I => \this_vga_signals.SUM_2_0_1\
        );

    \I__3238\ : InMux
    port map (
            O => \N__18270\,
            I => \N__18267\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__18267\,
            I => \this_vga_signals.mult1_un47_sum_c3_1_0\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__18264\,
            I => \this_vga_signals.mult1_un47_sum_c3_1_0_cascade_\
        );

    \I__3235\ : InMux
    port map (
            O => \N__18261\,
            I => \N__18252\
        );

    \I__3234\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18252\
        );

    \I__3233\ : InMux
    port map (
            O => \N__18259\,
            I => \N__18244\
        );

    \I__3232\ : InMux
    port map (
            O => \N__18258\,
            I => \N__18237\
        );

    \I__3231\ : InMux
    port map (
            O => \N__18257\,
            I => \N__18237\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__18252\,
            I => \N__18226\
        );

    \I__3229\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18215\
        );

    \I__3228\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18215\
        );

    \I__3227\ : InMux
    port map (
            O => \N__18249\,
            I => \N__18215\
        );

    \I__3226\ : InMux
    port map (
            O => \N__18248\,
            I => \N__18215\
        );

    \I__3225\ : InMux
    port map (
            O => \N__18247\,
            I => \N__18215\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__18244\,
            I => \N__18212\
        );

    \I__3223\ : InMux
    port map (
            O => \N__18243\,
            I => \N__18207\
        );

    \I__3222\ : InMux
    port map (
            O => \N__18242\,
            I => \N__18207\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__18237\,
            I => \N__18204\
        );

    \I__3220\ : InMux
    port map (
            O => \N__18236\,
            I => \N__18201\
        );

    \I__3219\ : InMux
    port map (
            O => \N__18235\,
            I => \N__18194\
        );

    \I__3218\ : InMux
    port map (
            O => \N__18234\,
            I => \N__18194\
        );

    \I__3217\ : InMux
    port map (
            O => \N__18233\,
            I => \N__18194\
        );

    \I__3216\ : InMux
    port map (
            O => \N__18232\,
            I => \N__18185\
        );

    \I__3215\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18185\
        );

    \I__3214\ : InMux
    port map (
            O => \N__18230\,
            I => \N__18185\
        );

    \I__3213\ : InMux
    port map (
            O => \N__18229\,
            I => \N__18185\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__18226\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__18215\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__18212\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__18207\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__18204\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__18201\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__18194\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__18185\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__3204\ : InMux
    port map (
            O => \N__18168\,
            I => \N__18165\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__18165\,
            I => \this_vga_signals.g2_4\
        );

    \I__3202\ : InMux
    port map (
            O => \N__18162\,
            I => \N__18159\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__18159\,
            I => \N__18156\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__18156\,
            I => \this_vga_signals.m12_0_1\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__18153\,
            I => \N__18150\
        );

    \I__3198\ : InMux
    port map (
            O => \N__18150\,
            I => \N__18147\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__18147\,
            I => \N__18144\
        );

    \I__3196\ : Odrv4
    port map (
            O => \N__18144\,
            I => \this_start_data_delay.N_400\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__18141\,
            I => \this_vga_signals.N_4_3_0_cascade_\
        );

    \I__3194\ : InMux
    port map (
            O => \N__18138\,
            I => \N__18135\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__18135\,
            I => \this_vga_signals.N_14_0\
        );

    \I__3192\ : InMux
    port map (
            O => \N__18132\,
            I => \N__18129\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__18129\,
            I => \this_vga_signals.g1\
        );

    \I__3190\ : InMux
    port map (
            O => \N__18126\,
            I => \N__18123\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__18123\,
            I => \this_vga_signals.g0_10_1\
        );

    \I__3188\ : InMux
    port map (
            O => \N__18120\,
            I => \N__18117\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__18117\,
            I => \this_vga_signals.N_24_mux\
        );

    \I__3186\ : InMux
    port map (
            O => \N__18114\,
            I => \N__18111\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__18111\,
            I => \this_vga_signals.g1_2\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__18108\,
            I => \N__18105\
        );

    \I__3183\ : InMux
    port map (
            O => \N__18105\,
            I => \N__18102\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__18102\,
            I => \this_vga_signals.g0_3_0_a3_3\
        );

    \I__3181\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18095\
        );

    \I__3180\ : InMux
    port map (
            O => \N__18098\,
            I => \N__18092\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__18095\,
            I => \N__18089\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__18092\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__18089\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__18084\,
            I => \this_vga_signals.mult1_un61_sum_axb2_0_cascade_\
        );

    \I__3175\ : InMux
    port map (
            O => \N__18081\,
            I => \N__18075\
        );

    \I__3174\ : InMux
    port map (
            O => \N__18080\,
            I => \N__18068\
        );

    \I__3173\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18068\
        );

    \I__3172\ : InMux
    port map (
            O => \N__18078\,
            I => \N__18068\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__18075\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__18068\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d
        );

    \I__3169\ : InMux
    port map (
            O => \N__18063\,
            I => \N__18060\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__18060\,
            I => \this_vga_signals.g2_0\
        );

    \I__3167\ : CascadeMux
    port map (
            O => \N__18057\,
            I => \N__18054\
        );

    \I__3166\ : InMux
    port map (
            O => \N__18054\,
            I => \N__18051\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__18051\,
            I => \N__18048\
        );

    \I__3164\ : Span4Mux_h
    port map (
            O => \N__18048\,
            I => \N__18044\
        );

    \I__3163\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18041\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__18044\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__18041\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__18036\,
            I => \this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d_cascade_\
        );

    \I__3159\ : InMux
    port map (
            O => \N__18033\,
            I => \N__18030\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__18030\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_0\
        );

    \I__3157\ : InMux
    port map (
            O => \N__18027\,
            I => \N__18023\
        );

    \I__3156\ : InMux
    port map (
            O => \N__18026\,
            I => \N__18020\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__18023\,
            I => \N__18017\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__18020\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_0\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__18017\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_0\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__18012\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_0_cascade_\
        );

    \I__3151\ : CascadeMux
    port map (
            O => \N__18009\,
            I => \N__18004\
        );

    \I__3150\ : InMux
    port map (
            O => \N__18008\,
            I => \N__18000\
        );

    \I__3149\ : InMux
    port map (
            O => \N__18007\,
            I => \N__17995\
        );

    \I__3148\ : InMux
    port map (
            O => \N__18004\,
            I => \N__17995\
        );

    \I__3147\ : InMux
    port map (
            O => \N__18003\,
            I => \N__17992\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__18000\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__17995\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__17992\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__3143\ : InMux
    port map (
            O => \N__17985\,
            I => \N__17982\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__17982\,
            I => \this_vga_signals.mult1_un75_sum_axb1_i_0\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__17979\,
            I => \this_vga_signals.N_4_2_cascade_\
        );

    \I__3140\ : InMux
    port map (
            O => \N__17976\,
            I => \N__17970\
        );

    \I__3139\ : InMux
    port map (
            O => \N__17975\,
            I => \N__17970\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__17970\,
            I => \this_vga_signals.if_m1_0_0\
        );

    \I__3137\ : InMux
    port map (
            O => \N__17967\,
            I => \N__17964\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__17964\,
            I => \N__17961\
        );

    \I__3135\ : Odrv12
    port map (
            O => \N__17961\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_d_0_0\
        );

    \I__3134\ : CascadeMux
    port map (
            O => \N__17958\,
            I => \N__17954\
        );

    \I__3133\ : InMux
    port map (
            O => \N__17957\,
            I => \N__17950\
        );

    \I__3132\ : InMux
    port map (
            O => \N__17954\,
            I => \N__17947\
        );

    \I__3131\ : InMux
    port map (
            O => \N__17953\,
            I => \N__17944\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__17950\,
            I => \N__17939\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__17947\,
            I => \N__17939\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__17944\,
            I => \this_vga_signals.mult1_un61_sum_axb2_0\
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__17939\,
            I => \this_vga_signals.mult1_un61_sum_axb2_0\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__17934\,
            I => \N__17930\
        );

    \I__3125\ : InMux
    port map (
            O => \N__17933\,
            I => \N__17925\
        );

    \I__3124\ : InMux
    port map (
            O => \N__17930\,
            I => \N__17920\
        );

    \I__3123\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17920\
        );

    \I__3122\ : InMux
    port map (
            O => \N__17928\,
            I => \N__17917\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__17925\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__17920\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__17917\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__17910\,
            I => \N__17907\
        );

    \I__3117\ : InMux
    port map (
            O => \N__17907\,
            I => \N__17903\
        );

    \I__3116\ : InMux
    port map (
            O => \N__17906\,
            I => \N__17900\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__17903\,
            I => \this_vga_signals.mult1_un75_sum_axb1_1\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__17900\,
            I => \this_vga_signals.mult1_un75_sum_axb1_1\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__17895\,
            I => \this_vga_signals.mult1_un54_sum_ac0_4_cascade_\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__17892\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__17889\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_0_2_cascade_\
        );

    \I__3110\ : InMux
    port map (
            O => \N__17886\,
            I => \N__17877\
        );

    \I__3109\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17877\
        );

    \I__3108\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17877\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__17877\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__17874\,
            I => \this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3_cascade_\
        );

    \I__3105\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17868\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__17868\,
            I => \this_vga_signals.mult1_un61_sum_c3_0\
        );

    \I__3103\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17862\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__17862\,
            I => \N__17859\
        );

    \I__3101\ : Span4Mux_h
    port map (
            O => \N__17859\,
            I => \N__17856\
        );

    \I__3100\ : Span4Mux_h
    port map (
            O => \N__17856\,
            I => \N__17853\
        );

    \I__3099\ : Span4Mux_h
    port map (
            O => \N__17853\,
            I => \N__17850\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__17850\,
            I => \this_vga_signals.if_m2\
        );

    \I__3097\ : InMux
    port map (
            O => \N__17847\,
            I => \N__17844\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__17844\,
            I => \this_vga_signals.if_m1_9_0\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__17841\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_cascade_\
        );

    \I__3094\ : InMux
    port map (
            O => \N__17838\,
            I => \N__17834\
        );

    \I__3093\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17831\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__17834\,
            I => \this_vga_signals.if_m2_3_1\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__17831\,
            I => \this_vga_signals.if_m2_3_1\
        );

    \I__3090\ : InMux
    port map (
            O => \N__17826\,
            I => \N__17823\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__17823\,
            I => \this_vga_signals.if_i4_mux\
        );

    \I__3088\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17817\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__17817\,
            I => \this_vga_signals.g0_1\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__17814\,
            I => \N__17811\
        );

    \I__3085\ : InMux
    port map (
            O => \N__17811\,
            I => \N__17808\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__17808\,
            I => \N__17805\
        );

    \I__3083\ : Span4Mux_h
    port map (
            O => \N__17805\,
            I => \N__17802\
        );

    \I__3082\ : Odrv4
    port map (
            O => \N__17802\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_a1_0\
        );

    \I__3081\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17796\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__17796\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_0_2_1\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__17793\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_0_2_1_cascade_\
        );

    \I__3078\ : CascadeMux
    port map (
            O => \N__17790\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1_cascade_\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__17787\,
            I => \N__17784\
        );

    \I__3076\ : InMux
    port map (
            O => \N__17784\,
            I => \N__17781\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__17781\,
            I => \M_this_state_d_0_sqmuxa_2\
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__17778\,
            I => \this_start_data_delay.N_65_cascade_\
        );

    \I__3073\ : InMux
    port map (
            O => \N__17775\,
            I => \N__17772\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__17772\,
            I => \N__17769\
        );

    \I__3071\ : Odrv4
    port map (
            O => \N__17769\,
            I => \this_start_data_delay.N_42_0\
        );

    \I__3070\ : InMux
    port map (
            O => \N__17766\,
            I => \N__17763\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__17763\,
            I => \N__17759\
        );

    \I__3068\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17756\
        );

    \I__3067\ : Span4Mux_v
    port map (
            O => \N__17759\,
            I => \N__17753\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__17756\,
            I => \N__17750\
        );

    \I__3065\ : Odrv4
    port map (
            O => \N__17753\,
            I => \this_start_data_delay.N_43_0\
        );

    \I__3064\ : Odrv4
    port map (
            O => \N__17750\,
            I => \this_start_data_delay.N_43_0\
        );

    \I__3063\ : IoInMux
    port map (
            O => \N__17745\,
            I => \N__17742\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__17742\,
            I => \N__17739\
        );

    \I__3061\ : Span4Mux_s1_h
    port map (
            O => \N__17739\,
            I => \N__17736\
        );

    \I__3060\ : Span4Mux_h
    port map (
            O => \N__17736\,
            I => \N__17731\
        );

    \I__3059\ : InMux
    port map (
            O => \N__17735\,
            I => \N__17728\
        );

    \I__3058\ : InMux
    port map (
            O => \N__17734\,
            I => \N__17725\
        );

    \I__3057\ : Sp12to4
    port map (
            O => \N__17731\,
            I => \N__17721\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__17728\,
            I => \N__17718\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__17725\,
            I => \N__17715\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__17724\,
            I => \N__17712\
        );

    \I__3053\ : Span12Mux_v
    port map (
            O => \N__17721\,
            I => \N__17707\
        );

    \I__3052\ : Span12Mux_s5_h
    port map (
            O => \N__17718\,
            I => \N__17707\
        );

    \I__3051\ : Span4Mux_h
    port map (
            O => \N__17715\,
            I => \N__17704\
        );

    \I__3050\ : InMux
    port map (
            O => \N__17712\,
            I => \N__17701\
        );

    \I__3049\ : Span12Mux_h
    port map (
            O => \N__17707\,
            I => \N__17698\
        );

    \I__3048\ : Span4Mux_v
    port map (
            O => \N__17704\,
            I => \N__17693\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__17701\,
            I => \N__17693\
        );

    \I__3046\ : Odrv12
    port map (
            O => \N__17698\,
            I => dma_0
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__17693\,
            I => dma_0
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__17688\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2_cascade_\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__17685\,
            I => \this_vga_signals.g0_i_x4_1_cascade_\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__17682\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_1_0_0_cascade_\
        );

    \I__3041\ : InMux
    port map (
            O => \N__17679\,
            I => \N__17676\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__17676\,
            I => \this_vga_signals.g0_9_N_3L3\
        );

    \I__3039\ : InMux
    port map (
            O => \N__17673\,
            I => \N__17670\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__17670\,
            I => \N__17667\
        );

    \I__3037\ : Odrv4
    port map (
            O => \N__17667\,
            I => \this_vga_signals.g0_i_a4_4_0_0\
        );

    \I__3036\ : CEMux
    port map (
            O => \N__17664\,
            I => \N__17660\
        );

    \I__3035\ : CEMux
    port map (
            O => \N__17663\,
            I => \N__17656\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__17660\,
            I => \N__17653\
        );

    \I__3033\ : CEMux
    port map (
            O => \N__17659\,
            I => \N__17650\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__17656\,
            I => \N__17646\
        );

    \I__3031\ : Span4Mux_v
    port map (
            O => \N__17653\,
            I => \N__17642\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__17650\,
            I => \N__17639\
        );

    \I__3029\ : CEMux
    port map (
            O => \N__17649\,
            I => \N__17636\
        );

    \I__3028\ : Span4Mux_v
    port map (
            O => \N__17646\,
            I => \N__17633\
        );

    \I__3027\ : CEMux
    port map (
            O => \N__17645\,
            I => \N__17630\
        );

    \I__3026\ : Span4Mux_h
    port map (
            O => \N__17642\,
            I => \N__17625\
        );

    \I__3025\ : Span4Mux_v
    port map (
            O => \N__17639\,
            I => \N__17625\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__17636\,
            I => \N__17622\
        );

    \I__3023\ : Span4Mux_h
    port map (
            O => \N__17633\,
            I => \N__17617\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__17630\,
            I => \N__17617\
        );

    \I__3021\ : Span4Mux_h
    port map (
            O => \N__17625\,
            I => \N__17612\
        );

    \I__3020\ : Span4Mux_h
    port map (
            O => \N__17622\,
            I => \N__17612\
        );

    \I__3019\ : Sp12to4
    port map (
            O => \N__17617\,
            I => \N__17609\
        );

    \I__3018\ : Span4Mux_h
    port map (
            O => \N__17612\,
            I => \N__17606\
        );

    \I__3017\ : Odrv12
    port map (
            O => \N__17609\,
            I => \N_1422_0\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__17606\,
            I => \N_1422_0\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__17601\,
            I => \M_this_state_d_0_sqmuxa_2_cascade_\
        );

    \I__3014\ : InMux
    port map (
            O => \N__17598\,
            I => \N__17594\
        );

    \I__3013\ : InMux
    port map (
            O => \N__17597\,
            I => \N__17591\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__17594\,
            I => \this_vga_signals.if_m1_0\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__17591\,
            I => \this_vga_signals.if_m1_0\
        );

    \I__3010\ : InMux
    port map (
            O => \N__17586\,
            I => \N__17583\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__17583\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__17580\,
            I => \N__17577\
        );

    \I__3007\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17574\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__17574\,
            I => \this_vga_signals.g0_3_0_a3\
        );

    \I__3005\ : InMux
    port map (
            O => \N__17571\,
            I => \N__17568\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__17568\,
            I => \this_vga_signals.g1_0\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__17565\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_1_0_cascade_\
        );

    \I__3002\ : InMux
    port map (
            O => \N__17562\,
            I => \N__17559\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__17559\,
            I => \this_vga_signals.g0_i_x4_7_0_0\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__17556\,
            I => \this_vga_signals.g0_9_N_2L1_cascade_\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__17553\,
            I => \this_vga_signals.mult1_un68_sum_c3_cascade_\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__17550\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_0_cascade_\
        );

    \I__2997\ : InMux
    port map (
            O => \N__17547\,
            I => \N__17543\
        );

    \I__2996\ : InMux
    port map (
            O => \N__17546\,
            I => \N__17540\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__17543\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__17540\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__17535\,
            I => \this_vga_signals.if_m2_3_1_cascade_\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__17532\,
            I => \this_vga_signals.g2_cascade_\
        );

    \I__2991\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17526\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__17526\,
            I => \this_vga_signals.g0_4\
        );

    \I__2989\ : InMux
    port map (
            O => \N__17523\,
            I => \N__17520\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__17520\,
            I => \this_vga_signals.g1_0_0\
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__17517\,
            I => \this_vga_signals.if_m1_0_cascade_\
        );

    \I__2986\ : InMux
    port map (
            O => \N__17514\,
            I => \N__17511\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__17511\,
            I => \N__17508\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__17508\,
            I => \this_vga_signals.N_129_i\
        );

    \I__2983\ : InMux
    port map (
            O => \N__17505\,
            I => \N__17502\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__17502\,
            I => \N__17499\
        );

    \I__2981\ : Sp12to4
    port map (
            O => \N__17499\,
            I => \N__17496\
        );

    \I__2980\ : Span12Mux_v
    port map (
            O => \N__17496\,
            I => \N__17493\
        );

    \I__2979\ : Odrv12
    port map (
            O => \N__17493\,
            I => \this_sprites_ram.mem_out_bus7_2\
        );

    \I__2978\ : InMux
    port map (
            O => \N__17490\,
            I => \N__17487\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__17487\,
            I => \N__17484\
        );

    \I__2976\ : Span4Mux_h
    port map (
            O => \N__17484\,
            I => \N__17481\
        );

    \I__2975\ : Span4Mux_h
    port map (
            O => \N__17481\,
            I => \N__17478\
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__17478\,
            I => \this_sprites_ram.mem_out_bus3_2\
        );

    \I__2973\ : InMux
    port map (
            O => \N__17475\,
            I => \N__17472\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__17472\,
            I => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\
        );

    \I__2971\ : InMux
    port map (
            O => \N__17469\,
            I => \N__17463\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__17468\,
            I => \N__17460\
        );

    \I__2969\ : InMux
    port map (
            O => \N__17467\,
            I => \N__17456\
        );

    \I__2968\ : InMux
    port map (
            O => \N__17466\,
            I => \N__17453\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__17463\,
            I => \N__17450\
        );

    \I__2966\ : InMux
    port map (
            O => \N__17460\,
            I => \N__17447\
        );

    \I__2965\ : InMux
    port map (
            O => \N__17459\,
            I => \N__17444\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__17456\,
            I => \N__17439\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__17453\,
            I => \N__17439\
        );

    \I__2962\ : Span4Mux_h
    port map (
            O => \N__17450\,
            I => \N__17430\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__17447\,
            I => \N__17430\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__17444\,
            I => \N__17430\
        );

    \I__2959\ : Span4Mux_v
    port map (
            O => \N__17439\,
            I => \N__17430\
        );

    \I__2958\ : Odrv4
    port map (
            O => \N__17430\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__2957\ : InMux
    port map (
            O => \N__17427\,
            I => \N__17424\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__17424\,
            I => \N__17421\
        );

    \I__2955\ : Span4Mux_h
    port map (
            O => \N__17421\,
            I => \N__17417\
        );

    \I__2954\ : InMux
    port map (
            O => \N__17420\,
            I => \N__17414\
        );

    \I__2953\ : Odrv4
    port map (
            O => \N__17417\,
            I => \this_ppu.M_state_q_srsts_i_a3_5_2\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__17414\,
            I => \this_ppu.M_state_q_srsts_i_a3_5_2\
        );

    \I__2951\ : InMux
    port map (
            O => \N__17409\,
            I => \N__17406\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__17406\,
            I => \N__17403\
        );

    \I__2949\ : Span4Mux_h
    port map (
            O => \N__17403\,
            I => \N__17399\
        );

    \I__2948\ : InMux
    port map (
            O => \N__17402\,
            I => \N__17396\
        );

    \I__2947\ : Odrv4
    port map (
            O => \N__17399\,
            I => \this_ppu.M_state_q_srsts_i_a3_4_2\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__17396\,
            I => \this_ppu.M_state_q_srsts_i_a3_4_2\
        );

    \I__2945\ : CascadeMux
    port map (
            O => \N__17391\,
            I => \N_2_cascade_\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__17388\,
            I => \this_vga_signals.N_6_1_cascade_\
        );

    \I__2943\ : InMux
    port map (
            O => \N__17385\,
            I => \N__17382\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__17382\,
            I => \this_vga_signals.vaddress_N_4_0\
        );

    \I__2941\ : InMux
    port map (
            O => \N__17379\,
            I => \N__17376\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__17376\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0\
        );

    \I__2939\ : InMux
    port map (
            O => \N__17373\,
            I => \N__17370\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__17370\,
            I => \this_vga_signals.mult1_un75_sum_axb1_i_1\
        );

    \I__2937\ : InMux
    port map (
            O => \N__17367\,
            I => \N__17364\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__17364\,
            I => \this_vga_signals.N_7_0\
        );

    \I__2935\ : CEMux
    port map (
            O => \N__17361\,
            I => \N__17358\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__17358\,
            I => \N__17354\
        );

    \I__2933\ : CEMux
    port map (
            O => \N__17357\,
            I => \N__17349\
        );

    \I__2932\ : Span4Mux_v
    port map (
            O => \N__17354\,
            I => \N__17346\
        );

    \I__2931\ : CEMux
    port map (
            O => \N__17353\,
            I => \N__17343\
        );

    \I__2930\ : CEMux
    port map (
            O => \N__17352\,
            I => \N__17340\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__17349\,
            I => \N__17336\
        );

    \I__2928\ : Span4Mux_h
    port map (
            O => \N__17346\,
            I => \N__17331\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__17343\,
            I => \N__17331\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__17340\,
            I => \N__17328\
        );

    \I__2925\ : CEMux
    port map (
            O => \N__17339\,
            I => \N__17325\
        );

    \I__2924\ : Span4Mux_h
    port map (
            O => \N__17336\,
            I => \N__17322\
        );

    \I__2923\ : Span4Mux_h
    port map (
            O => \N__17331\,
            I => \N__17315\
        );

    \I__2922\ : Span4Mux_v
    port map (
            O => \N__17328\,
            I => \N__17315\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__17325\,
            I => \N__17315\
        );

    \I__2920\ : Span4Mux_h
    port map (
            O => \N__17322\,
            I => \N__17312\
        );

    \I__2919\ : Sp12to4
    port map (
            O => \N__17315\,
            I => \N__17309\
        );

    \I__2918\ : Odrv4
    port map (
            O => \N__17312\,
            I => \N_1438_0\
        );

    \I__2917\ : Odrv12
    port map (
            O => \N__17309\,
            I => \N_1438_0\
        );

    \I__2916\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17301\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__17301\,
            I => \this_start_data_delay.port_data_rw_0_a2Z0Z_1\
        );

    \I__2914\ : IoInMux
    port map (
            O => \N__17298\,
            I => \N__17295\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__17295\,
            I => \N__17292\
        );

    \I__2912\ : Span4Mux_s1_h
    port map (
            O => \N__17292\,
            I => \N__17289\
        );

    \I__2911\ : Span4Mux_h
    port map (
            O => \N__17289\,
            I => \N__17286\
        );

    \I__2910\ : Span4Mux_h
    port map (
            O => \N__17286\,
            I => \N__17283\
        );

    \I__2909\ : Sp12to4
    port map (
            O => \N__17283\,
            I => \N__17280\
        );

    \I__2908\ : Span12Mux_v
    port map (
            O => \N__17280\,
            I => \N__17277\
        );

    \I__2907\ : Odrv12
    port map (
            O => \N__17277\,
            I => port_data_rw_0_i
        );

    \I__2906\ : InMux
    port map (
            O => \N__17274\,
            I => \N__17271\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__17271\,
            I => \N__17268\
        );

    \I__2904\ : Span12Mux_v
    port map (
            O => \N__17268\,
            I => \N__17265\
        );

    \I__2903\ : Odrv12
    port map (
            O => \N__17265\,
            I => \this_sprites_ram.mem_out_bus5_2\
        );

    \I__2902\ : InMux
    port map (
            O => \N__17262\,
            I => \N__17259\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__17259\,
            I => \N__17256\
        );

    \I__2900\ : Span12Mux_v
    port map (
            O => \N__17256\,
            I => \N__17253\
        );

    \I__2899\ : Odrv12
    port map (
            O => \N__17253\,
            I => \this_sprites_ram.mem_out_bus1_2\
        );

    \I__2898\ : InMux
    port map (
            O => \N__17250\,
            I => \N__17247\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__17247\,
            I => \N__17244\
        );

    \I__2896\ : Span4Mux_h
    port map (
            O => \N__17244\,
            I => \N__17241\
        );

    \I__2895\ : Span4Mux_h
    port map (
            O => \N__17241\,
            I => \N__17238\
        );

    \I__2894\ : Span4Mux_h
    port map (
            O => \N__17238\,
            I => \N__17235\
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__17235\,
            I => \this_delay_clk.M_pipe_qZ0Z_2\
        );

    \I__2892\ : InMux
    port map (
            O => \N__17232\,
            I => \N__17229\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__17229\,
            I => \N__17226\
        );

    \I__2890\ : Span4Mux_h
    port map (
            O => \N__17226\,
            I => \N__17223\
        );

    \I__2889\ : Span4Mux_h
    port map (
            O => \N__17223\,
            I => \N__17220\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__17220\,
            I => \this_sprites_ram.mem_out_bus4_2\
        );

    \I__2887\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17214\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__17214\,
            I => \N__17211\
        );

    \I__2885\ : Span12Mux_v
    port map (
            O => \N__17211\,
            I => \N__17208\
        );

    \I__2884\ : Span12Mux_v
    port map (
            O => \N__17208\,
            I => \N__17205\
        );

    \I__2883\ : Odrv12
    port map (
            O => \N__17205\,
            I => \this_sprites_ram.mem_out_bus0_2\
        );

    \I__2882\ : CascadeMux
    port map (
            O => \N__17202\,
            I => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_\
        );

    \I__2881\ : InMux
    port map (
            O => \N__17199\,
            I => \N__17196\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__17196\,
            I => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__17193\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\
        );

    \I__2878\ : InMux
    port map (
            O => \N__17190\,
            I => \N__17186\
        );

    \I__2877\ : InMux
    port map (
            O => \N__17189\,
            I => \N__17183\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__17186\,
            I => \N__17179\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__17183\,
            I => \N__17176\
        );

    \I__2874\ : InMux
    port map (
            O => \N__17182\,
            I => \N__17173\
        );

    \I__2873\ : Span12Mux_h
    port map (
            O => \N__17179\,
            I => \N__17170\
        );

    \I__2872\ : Span4Mux_h
    port map (
            O => \N__17176\,
            I => \N__17167\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__17173\,
            I => \N__17164\
        );

    \I__2870\ : Odrv12
    port map (
            O => \N__17170\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__2869\ : Odrv4
    port map (
            O => \N__17167\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__2868\ : Odrv12
    port map (
            O => \N__17164\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__2867\ : InMux
    port map (
            O => \N__17157\,
            I => \N__17154\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__17154\,
            I => \this_ppu.un10_sprites_addr_cry_2_c_RNIQP7BZ0\
        );

    \I__2865\ : InMux
    port map (
            O => \N__17151\,
            I => \N__17148\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__17148\,
            I => \N__17145\
        );

    \I__2863\ : Span4Mux_v
    port map (
            O => \N__17145\,
            I => \N__17142\
        );

    \I__2862\ : Span4Mux_v
    port map (
            O => \N__17142\,
            I => \N__17139\
        );

    \I__2861\ : Span4Mux_h
    port map (
            O => \N__17139\,
            I => \N__17136\
        );

    \I__2860\ : Span4Mux_h
    port map (
            O => \N__17136\,
            I => \N__17133\
        );

    \I__2859\ : Odrv4
    port map (
            O => \N__17133\,
            I => \M_this_map_ram_read_data_5\
        );

    \I__2858\ : InMux
    port map (
            O => \N__17130\,
            I => \N__17125\
        );

    \I__2857\ : InMux
    port map (
            O => \N__17129\,
            I => \N__17122\
        );

    \I__2856\ : InMux
    port map (
            O => \N__17128\,
            I => \N__17115\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__17125\,
            I => \N__17112\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__17122\,
            I => \N__17109\
        );

    \I__2853\ : InMux
    port map (
            O => \N__17121\,
            I => \N__17106\
        );

    \I__2852\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17103\
        );

    \I__2851\ : InMux
    port map (
            O => \N__17119\,
            I => \N__17098\
        );

    \I__2850\ : InMux
    port map (
            O => \N__17118\,
            I => \N__17098\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__17115\,
            I => \N__17095\
        );

    \I__2848\ : Span4Mux_h
    port map (
            O => \N__17112\,
            I => \N__17092\
        );

    \I__2847\ : Span4Mux_h
    port map (
            O => \N__17109\,
            I => \N__17089\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__17106\,
            I => \N__17086\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__17103\,
            I => \N__17083\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__17098\,
            I => \N__17080\
        );

    \I__2843\ : Span4Mux_h
    port map (
            O => \N__17095\,
            I => \N__17071\
        );

    \I__2842\ : Span4Mux_v
    port map (
            O => \N__17092\,
            I => \N__17071\
        );

    \I__2841\ : Span4Mux_v
    port map (
            O => \N__17089\,
            I => \N__17071\
        );

    \I__2840\ : Span4Mux_h
    port map (
            O => \N__17086\,
            I => \N__17068\
        );

    \I__2839\ : Span4Mux_v
    port map (
            O => \N__17083\,
            I => \N__17063\
        );

    \I__2838\ : Span4Mux_h
    port map (
            O => \N__17080\,
            I => \N__17063\
        );

    \I__2837\ : InMux
    port map (
            O => \N__17079\,
            I => \N__17058\
        );

    \I__2836\ : InMux
    port map (
            O => \N__17078\,
            I => \N__17058\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__17071\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__2834\ : Odrv4
    port map (
            O => \N__17068\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__17063\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__17058\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__17049\,
            I => \this_vga_signals.mult1_un75_sum_c3_0_0_0_0_cascade_\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__17046\,
            I => \N__17043\
        );

    \I__2829\ : InMux
    port map (
            O => \N__17043\,
            I => \N__17040\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__17040\,
            I => \N__17037\
        );

    \I__2827\ : Span4Mux_v
    port map (
            O => \N__17037\,
            I => \N__17034\
        );

    \I__2826\ : Span4Mux_h
    port map (
            O => \N__17034\,
            I => \N__17031\
        );

    \I__2825\ : Span4Mux_h
    port map (
            O => \N__17031\,
            I => \N__17028\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__17028\,
            I => \M_this_vga_signals_address_7\
        );

    \I__2823\ : InMux
    port map (
            O => \N__17025\,
            I => \N__17022\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__17022\,
            I => \this_vga_signals.un6_vvisibilitylt9_0\
        );

    \I__2821\ : InMux
    port map (
            O => \N__17019\,
            I => \N__17016\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__17016\,
            I => \this_vga_signals.g2_2\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__17013\,
            I => \this_vga_signals.SUM_2_1_cascade_\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__17010\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_1_1_cascade_\
        );

    \I__2817\ : InMux
    port map (
            O => \N__17007\,
            I => \N__17004\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__17004\,
            I => \this_vga_signals.N_4_0_0_0\
        );

    \I__2815\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16998\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__16998\,
            I => \this_vga_signals.g3_2_0\
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__16995\,
            I => \this_vga_signals.N_6_cascade_\
        );

    \I__2812\ : InMux
    port map (
            O => \N__16992\,
            I => \N__16989\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__16989\,
            I => \this_vga_signals.g4\
        );

    \I__2810\ : InMux
    port map (
            O => \N__16986\,
            I => \N__16983\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__16983\,
            I => \N__16979\
        );

    \I__2808\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16975\
        );

    \I__2807\ : Span4Mux_v
    port map (
            O => \N__16979\,
            I => \N__16969\
        );

    \I__2806\ : InMux
    port map (
            O => \N__16978\,
            I => \N__16966\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__16975\,
            I => \N__16963\
        );

    \I__2804\ : InMux
    port map (
            O => \N__16974\,
            I => \N__16956\
        );

    \I__2803\ : InMux
    port map (
            O => \N__16973\,
            I => \N__16956\
        );

    \I__2802\ : InMux
    port map (
            O => \N__16972\,
            I => \N__16956\
        );

    \I__2801\ : Odrv4
    port map (
            O => \N__16969\,
            I => \this_ppu.M_last_q\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__16966\,
            I => \this_ppu.M_last_q\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__16963\,
            I => \this_ppu.M_last_q\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__16956\,
            I => \this_ppu.M_last_q\
        );

    \I__2797\ : InMux
    port map (
            O => \N__16947\,
            I => \N__16940\
        );

    \I__2796\ : InMux
    port map (
            O => \N__16946\,
            I => \N__16937\
        );

    \I__2795\ : InMux
    port map (
            O => \N__16945\,
            I => \N__16930\
        );

    \I__2794\ : InMux
    port map (
            O => \N__16944\,
            I => \N__16930\
        );

    \I__2793\ : InMux
    port map (
            O => \N__16943\,
            I => \N__16930\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__16940\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__16937\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__16930\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__2789\ : InMux
    port map (
            O => \N__16923\,
            I => \N__16918\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__16922\,
            I => \N__16913\
        );

    \I__2787\ : InMux
    port map (
            O => \N__16921\,
            I => \N__16910\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__16918\,
            I => \N__16907\
        );

    \I__2785\ : InMux
    port map (
            O => \N__16917\,
            I => \N__16904\
        );

    \I__2784\ : InMux
    port map (
            O => \N__16916\,
            I => \N__16901\
        );

    \I__2783\ : InMux
    port map (
            O => \N__16913\,
            I => \N__16898\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__16910\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__16907\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__16904\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__16901\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__16898\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__16887\,
            I => \N__16882\
        );

    \I__2776\ : InMux
    port map (
            O => \N__16886\,
            I => \N__16877\
        );

    \I__2775\ : InMux
    port map (
            O => \N__16885\,
            I => \N__16877\
        );

    \I__2774\ : InMux
    port map (
            O => \N__16882\,
            I => \N__16873\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__16877\,
            I => \N__16868\
        );

    \I__2772\ : InMux
    port map (
            O => \N__16876\,
            I => \N__16865\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__16873\,
            I => \N__16862\
        );

    \I__2770\ : InMux
    port map (
            O => \N__16872\,
            I => \N__16857\
        );

    \I__2769\ : InMux
    port map (
            O => \N__16871\,
            I => \N__16857\
        );

    \I__2768\ : Odrv4
    port map (
            O => \N__16868\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__16865\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__2766\ : Odrv4
    port map (
            O => \N__16862\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__16857\,
            I => \this_ppu.M_state_d_0_sqmuxa\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__16848\,
            I => \N__16845\
        );

    \I__2763\ : InMux
    port map (
            O => \N__16845\,
            I => \N__16842\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__16842\,
            I => \N__16839\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__16839\,
            I => \N__16836\
        );

    \I__2760\ : Sp12to4
    port map (
            O => \N__16836\,
            I => \N__16829\
        );

    \I__2759\ : CascadeMux
    port map (
            O => \N__16835\,
            I => \N__16826\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__16834\,
            I => \N__16822\
        );

    \I__2757\ : InMux
    port map (
            O => \N__16833\,
            I => \N__16817\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__16832\,
            I => \N__16814\
        );

    \I__2755\ : Span12Mux_v
    port map (
            O => \N__16829\,
            I => \N__16811\
        );

    \I__2754\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16804\
        );

    \I__2753\ : InMux
    port map (
            O => \N__16825\,
            I => \N__16804\
        );

    \I__2752\ : InMux
    port map (
            O => \N__16822\,
            I => \N__16804\
        );

    \I__2751\ : InMux
    port map (
            O => \N__16821\,
            I => \N__16799\
        );

    \I__2750\ : InMux
    port map (
            O => \N__16820\,
            I => \N__16799\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__16817\,
            I => \N__16796\
        );

    \I__2748\ : InMux
    port map (
            O => \N__16814\,
            I => \N__16793\
        );

    \I__2747\ : Odrv12
    port map (
            O => \N__16811\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__16804\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__16799\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__16796\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__16793\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__16782\,
            I => \N__16779\
        );

    \I__2741\ : CascadeBuf
    port map (
            O => \N__16779\,
            I => \N__16776\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__16776\,
            I => \N__16772\
        );

    \I__2739\ : InMux
    port map (
            O => \N__16775\,
            I => \N__16768\
        );

    \I__2738\ : InMux
    port map (
            O => \N__16772\,
            I => \N__16765\
        );

    \I__2737\ : InMux
    port map (
            O => \N__16771\,
            I => \N__16762\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__16768\,
            I => \N__16759\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__16765\,
            I => \N__16756\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__16762\,
            I => \N__16752\
        );

    \I__2733\ : Span4Mux_v
    port map (
            O => \N__16759\,
            I => \N__16748\
        );

    \I__2732\ : Sp12to4
    port map (
            O => \N__16756\,
            I => \N__16745\
        );

    \I__2731\ : InMux
    port map (
            O => \N__16755\,
            I => \N__16742\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__16752\,
            I => \N__16739\
        );

    \I__2729\ : InMux
    port map (
            O => \N__16751\,
            I => \N__16736\
        );

    \I__2728\ : Sp12to4
    port map (
            O => \N__16748\,
            I => \N__16731\
        );

    \I__2727\ : Span12Mux_v
    port map (
            O => \N__16745\,
            I => \N__16731\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__16742\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__16739\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__16736\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__2723\ : Odrv12
    port map (
            O => \N__16731\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__2722\ : InMux
    port map (
            O => \N__16722\,
            I => \N__16713\
        );

    \I__2721\ : InMux
    port map (
            O => \N__16721\,
            I => \N__16713\
        );

    \I__2720\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16713\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__16713\,
            I => \N__16709\
        );

    \I__2718\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16706\
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__16709\,
            I => \this_ppu.un1_M_vaddress_q_c3\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__16706\,
            I => \this_ppu.un1_M_vaddress_q_c3\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__16701\,
            I => \N__16698\
        );

    \I__2714\ : CascadeBuf
    port map (
            O => \N__16698\,
            I => \N__16695\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__16695\,
            I => \N__16692\
        );

    \I__2712\ : InMux
    port map (
            O => \N__16692\,
            I => \N__16688\
        );

    \I__2711\ : InMux
    port map (
            O => \N__16691\,
            I => \N__16683\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__16688\,
            I => \N__16679\
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__16687\,
            I => \N__16676\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__16686\,
            I => \N__16673\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__16683\,
            I => \N__16669\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__16682\,
            I => \N__16666\
        );

    \I__2705\ : Sp12to4
    port map (
            O => \N__16679\,
            I => \N__16663\
        );

    \I__2704\ : InMux
    port map (
            O => \N__16676\,
            I => \N__16656\
        );

    \I__2703\ : InMux
    port map (
            O => \N__16673\,
            I => \N__16656\
        );

    \I__2702\ : InMux
    port map (
            O => \N__16672\,
            I => \N__16656\
        );

    \I__2701\ : Span4Mux_v
    port map (
            O => \N__16669\,
            I => \N__16653\
        );

    \I__2700\ : InMux
    port map (
            O => \N__16666\,
            I => \N__16650\
        );

    \I__2699\ : Span12Mux_v
    port map (
            O => \N__16663\,
            I => \N__16647\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__16656\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__16653\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__16650\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__2695\ : Odrv12
    port map (
            O => \N__16647\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__16638\,
            I => \N__16635\
        );

    \I__2693\ : CascadeBuf
    port map (
            O => \N__16635\,
            I => \N__16632\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__16632\,
            I => \N__16629\
        );

    \I__2691\ : InMux
    port map (
            O => \N__16629\,
            I => \N__16626\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__16626\,
            I => \N__16622\
        );

    \I__2689\ : InMux
    port map (
            O => \N__16625\,
            I => \N__16619\
        );

    \I__2688\ : Span4Mux_h
    port map (
            O => \N__16622\,
            I => \N__16616\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__16619\,
            I => \N__16611\
        );

    \I__2686\ : Span4Mux_h
    port map (
            O => \N__16616\,
            I => \N__16607\
        );

    \I__2685\ : InMux
    port map (
            O => \N__16615\,
            I => \N__16602\
        );

    \I__2684\ : InMux
    port map (
            O => \N__16614\,
            I => \N__16602\
        );

    \I__2683\ : Span4Mux_v
    port map (
            O => \N__16611\,
            I => \N__16599\
        );

    \I__2682\ : InMux
    port map (
            O => \N__16610\,
            I => \N__16596\
        );

    \I__2681\ : Span4Mux_v
    port map (
            O => \N__16607\,
            I => \N__16593\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__16602\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__16599\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__16596\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__2677\ : Odrv4
    port map (
            O => \N__16593\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__2676\ : SRMux
    port map (
            O => \N__16584\,
            I => \N__16579\
        );

    \I__2675\ : SRMux
    port map (
            O => \N__16583\,
            I => \N__16576\
        );

    \I__2674\ : SRMux
    port map (
            O => \N__16582\,
            I => \N__16573\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__16579\,
            I => \N__16570\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__16576\,
            I => \N__16567\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__16573\,
            I => \N__16564\
        );

    \I__2670\ : Span4Mux_v
    port map (
            O => \N__16570\,
            I => \N__16561\
        );

    \I__2669\ : Span4Mux_v
    port map (
            O => \N__16567\,
            I => \N__16558\
        );

    \I__2668\ : Span4Mux_h
    port map (
            O => \N__16564\,
            I => \N__16555\
        );

    \I__2667\ : Odrv4
    port map (
            O => \N__16561\,
            I => \this_ppu.M_state_q_RNIELANCZ0Z_0\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__16558\,
            I => \this_ppu.M_state_q_RNIELANCZ0Z_0\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__16555\,
            I => \this_ppu.M_state_q_RNIELANCZ0Z_0\
        );

    \I__2664\ : IoInMux
    port map (
            O => \N__16548\,
            I => \N__16545\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__16545\,
            I => \N__16542\
        );

    \I__2662\ : Span12Mux_s5_h
    port map (
            O => \N__16542\,
            I => \N__16538\
        );

    \I__2661\ : InMux
    port map (
            O => \N__16541\,
            I => \N__16535\
        );

    \I__2660\ : Span12Mux_h
    port map (
            O => \N__16538\,
            I => \N__16532\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__16535\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI4KCU6Z0Z_9\
        );

    \I__2658\ : Odrv12
    port map (
            O => \N__16532\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI4KCU6Z0Z_9\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__16527\,
            I => \this_vga_signals.g1_2_0_0_cascade_\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__16524\,
            I => \M_this_state_q_ns_17_cascade_\
        );

    \I__2655\ : CEMux
    port map (
            O => \N__16521\,
            I => \N__16517\
        );

    \I__2654\ : CEMux
    port map (
            O => \N__16520\,
            I => \N__16513\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__16517\,
            I => \N__16509\
        );

    \I__2652\ : CEMux
    port map (
            O => \N__16516\,
            I => \N__16506\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__16513\,
            I => \N__16503\
        );

    \I__2650\ : CEMux
    port map (
            O => \N__16512\,
            I => \N__16500\
        );

    \I__2649\ : Span4Mux_v
    port map (
            O => \N__16509\,
            I => \N__16494\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__16506\,
            I => \N__16494\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__16503\,
            I => \N__16489\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__16500\,
            I => \N__16489\
        );

    \I__2645\ : CEMux
    port map (
            O => \N__16499\,
            I => \N__16486\
        );

    \I__2644\ : Span4Mux_h
    port map (
            O => \N__16494\,
            I => \N__16483\
        );

    \I__2643\ : Span4Mux_h
    port map (
            O => \N__16489\,
            I => \N__16480\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__16486\,
            I => \N__16477\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__16483\,
            I => \M_this_state_q_ns_0_17\
        );

    \I__2640\ : Odrv4
    port map (
            O => \N__16480\,
            I => \M_this_state_q_ns_0_17\
        );

    \I__2639\ : Odrv12
    port map (
            O => \N__16477\,
            I => \M_this_state_q_ns_0_17\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__16470\,
            I => \N__16467\
        );

    \I__2637\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16464\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__16464\,
            I => \N__16461\
        );

    \I__2635\ : Span4Mux_v
    port map (
            O => \N__16461\,
            I => \N__16458\
        );

    \I__2634\ : Sp12to4
    port map (
            O => \N__16458\,
            I => \N__16455\
        );

    \I__2633\ : Span12Mux_h
    port map (
            O => \N__16455\,
            I => \N__16452\
        );

    \I__2632\ : Odrv12
    port map (
            O => \N__16452\,
            I => \M_this_map_ram_read_data_6\
        );

    \I__2631\ : InMux
    port map (
            O => \N__16449\,
            I => \N__16445\
        );

    \I__2630\ : InMux
    port map (
            O => \N__16448\,
            I => \N__16442\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__16445\,
            I => \N__16437\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__16442\,
            I => \N__16437\
        );

    \I__2627\ : Span4Mux_h
    port map (
            O => \N__16437\,
            I => \N__16434\
        );

    \I__2626\ : Span4Mux_h
    port map (
            O => \N__16434\,
            I => \N__16431\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__16431\,
            I => \M_this_oam_ram_read_data_8\
        );

    \I__2624\ : InMux
    port map (
            O => \N__16428\,
            I => \N__16425\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__16425\,
            I => \this_ppu.M_this_oam_ram_read_data_iZ0Z_8\
        );

    \I__2622\ : InMux
    port map (
            O => \N__16422\,
            I => \N__16419\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__16419\,
            I => \M_this_oam_ram_read_data_i_9\
        );

    \I__2620\ : InMux
    port map (
            O => \N__16416\,
            I => \N__16413\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__16413\,
            I => \this_ppu.un10_sprites_addr_cry_0_c_RNIMJ5BZ0\
        );

    \I__2618\ : InMux
    port map (
            O => \N__16410\,
            I => \this_ppu.un10_sprites_addr_cry_0\
        );

    \I__2617\ : InMux
    port map (
            O => \N__16407\,
            I => \N__16404\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__16404\,
            I => \N__16401\
        );

    \I__2615\ : Span4Mux_h
    port map (
            O => \N__16401\,
            I => \N__16398\
        );

    \I__2614\ : Span4Mux_h
    port map (
            O => \N__16398\,
            I => \N__16395\
        );

    \I__2613\ : Odrv4
    port map (
            O => \N__16395\,
            I => \M_this_oam_ram_read_data_i_10\
        );

    \I__2612\ : InMux
    port map (
            O => \N__16392\,
            I => \this_ppu.un10_sprites_addr_cry_1\
        );

    \I__2611\ : InMux
    port map (
            O => \N__16389\,
            I => \N__16386\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__16386\,
            I => \N__16383\
        );

    \I__2609\ : Span4Mux_h
    port map (
            O => \N__16383\,
            I => \N__16380\
        );

    \I__2608\ : Span4Mux_h
    port map (
            O => \N__16380\,
            I => \N__16377\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__16377\,
            I => \M_this_oam_ram_read_data_i_11\
        );

    \I__2606\ : InMux
    port map (
            O => \N__16374\,
            I => \this_ppu.un10_sprites_addr_cry_2\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__16371\,
            I => \N__16368\
        );

    \I__2604\ : InMux
    port map (
            O => \N__16368\,
            I => \N__16365\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__16365\,
            I => \N__16362\
        );

    \I__2602\ : Span4Mux_h
    port map (
            O => \N__16362\,
            I => \N__16359\
        );

    \I__2601\ : Span4Mux_h
    port map (
            O => \N__16359\,
            I => \N__16356\
        );

    \I__2600\ : Odrv4
    port map (
            O => \N__16356\,
            I => \M_this_oam_ram_read_data_i_12\
        );

    \I__2599\ : InMux
    port map (
            O => \N__16353\,
            I => \N__16350\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__16350\,
            I => \this_ppu.un10_sprites_addr_cry_3_c_RNISS8BZ0\
        );

    \I__2597\ : InMux
    port map (
            O => \N__16347\,
            I => \this_ppu.un10_sprites_addr_cry_3\
        );

    \I__2596\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16341\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__16341\,
            I => \N__16338\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__16338\,
            I => \N__16335\
        );

    \I__2593\ : Span4Mux_h
    port map (
            O => \N__16335\,
            I => \N__16332\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__16332\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__2591\ : InMux
    port map (
            O => \N__16329\,
            I => \this_ppu.un10_sprites_addr_cry_4\
        );

    \I__2590\ : InMux
    port map (
            O => \N__16326\,
            I => \N__16323\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__16323\,
            I => \this_reset_cond.M_stage_qZ0Z_6\
        );

    \I__2588\ : InMux
    port map (
            O => \N__16320\,
            I => \N__16305\
        );

    \I__2587\ : InMux
    port map (
            O => \N__16319\,
            I => \N__16305\
        );

    \I__2586\ : InMux
    port map (
            O => \N__16318\,
            I => \N__16305\
        );

    \I__2585\ : InMux
    port map (
            O => \N__16317\,
            I => \N__16305\
        );

    \I__2584\ : InMux
    port map (
            O => \N__16316\,
            I => \N__16305\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__16305\,
            I => \N__16299\
        );

    \I__2582\ : InMux
    port map (
            O => \N__16304\,
            I => \N__16294\
        );

    \I__2581\ : InMux
    port map (
            O => \N__16303\,
            I => \N__16294\
        );

    \I__2580\ : InMux
    port map (
            O => \N__16302\,
            I => \N__16290\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__16299\,
            I => \N__16287\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__16294\,
            I => \N__16284\
        );

    \I__2577\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16281\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__16290\,
            I => \N__16277\
        );

    \I__2575\ : Span4Mux_v
    port map (
            O => \N__16287\,
            I => \N__16270\
        );

    \I__2574\ : Span4Mux_h
    port map (
            O => \N__16284\,
            I => \N__16270\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__16281\,
            I => \N__16270\
        );

    \I__2572\ : InMux
    port map (
            O => \N__16280\,
            I => \N__16267\
        );

    \I__2571\ : Span4Mux_h
    port map (
            O => \N__16277\,
            I => \N__16264\
        );

    \I__2570\ : Span4Mux_v
    port map (
            O => \N__16270\,
            I => \N__16261\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__16267\,
            I => \N__16258\
        );

    \I__2568\ : Span4Mux_v
    port map (
            O => \N__16264\,
            I => \N__16255\
        );

    \I__2567\ : Span4Mux_v
    port map (
            O => \N__16261\,
            I => \N__16252\
        );

    \I__2566\ : Span12Mux_h
    port map (
            O => \N__16258\,
            I => \N__16249\
        );

    \I__2565\ : Span4Mux_v
    port map (
            O => \N__16255\,
            I => \N__16246\
        );

    \I__2564\ : Span4Mux_v
    port map (
            O => \N__16252\,
            I => \N__16243\
        );

    \I__2563\ : Span12Mux_v
    port map (
            O => \N__16249\,
            I => \N__16240\
        );

    \I__2562\ : Span4Mux_v
    port map (
            O => \N__16246\,
            I => \N__16237\
        );

    \I__2561\ : IoSpan4Mux
    port map (
            O => \N__16243\,
            I => \N__16234\
        );

    \I__2560\ : Odrv12
    port map (
            O => \N__16240\,
            I => rst_n_c
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__16237\,
            I => rst_n_c
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__16234\,
            I => rst_n_c
        );

    \I__2557\ : InMux
    port map (
            O => \N__16227\,
            I => \N__16224\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__16224\,
            I => \this_reset_cond.M_stage_qZ0Z_7\
        );

    \I__2555\ : InMux
    port map (
            O => \N__16221\,
            I => \N__16218\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__16218\,
            I => \this_reset_cond.M_stage_qZ0Z_8\
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__16215\,
            I => \N__16212\
        );

    \I__2552\ : InMux
    port map (
            O => \N__16212\,
            I => \N__16209\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__16209\,
            I => \this_vga_signals.vaddress_ac0_9_0_a0_2\
        );

    \I__2550\ : InMux
    port map (
            O => \N__16206\,
            I => \N__16202\
        );

    \I__2549\ : InMux
    port map (
            O => \N__16205\,
            I => \N__16199\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__16202\,
            I => \N__16192\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__16199\,
            I => \N__16192\
        );

    \I__2546\ : InMux
    port map (
            O => \N__16198\,
            I => \N__16189\
        );

    \I__2545\ : InMux
    port map (
            O => \N__16197\,
            I => \N__16186\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__16192\,
            I => \N__16183\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__16189\,
            I => \this_ppu.M_vaddress_qZ0Z_6\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__16186\,
            I => \this_ppu.M_vaddress_qZ0Z_6\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__16183\,
            I => \this_ppu.M_vaddress_qZ0Z_6\
        );

    \I__2540\ : InMux
    port map (
            O => \N__16176\,
            I => \N__16172\
        );

    \I__2539\ : InMux
    port map (
            O => \N__16175\,
            I => \N__16169\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__16172\,
            I => \N__16166\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__16169\,
            I => \N__16163\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__16166\,
            I => \this_ppu.un1_M_vaddress_q_c5\
        );

    \I__2535\ : Odrv4
    port map (
            O => \N__16163\,
            I => \this_ppu.un1_M_vaddress_q_c5\
        );

    \I__2534\ : InMux
    port map (
            O => \N__16158\,
            I => \N__16154\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__16157\,
            I => \N__16151\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__16154\,
            I => \N__16148\
        );

    \I__2531\ : InMux
    port map (
            O => \N__16151\,
            I => \N__16145\
        );

    \I__2530\ : Span4Mux_v
    port map (
            O => \N__16148\,
            I => \N__16142\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__16145\,
            I => \this_ppu.M_vaddress_qZ0Z_7\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__16142\,
            I => \this_ppu.M_vaddress_qZ0Z_7\
        );

    \I__2527\ : IoInMux
    port map (
            O => \N__16137\,
            I => \N__16132\
        );

    \I__2526\ : IoInMux
    port map (
            O => \N__16136\,
            I => \N__16127\
        );

    \I__2525\ : IoInMux
    port map (
            O => \N__16135\,
            I => \N__16124\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__16132\,
            I => \N__16117\
        );

    \I__2523\ : IoInMux
    port map (
            O => \N__16131\,
            I => \N__16114\
        );

    \I__2522\ : IoInMux
    port map (
            O => \N__16130\,
            I => \N__16109\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__16127\,
            I => \N__16104\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__16124\,
            I => \N__16104\
        );

    \I__2519\ : IoInMux
    port map (
            O => \N__16123\,
            I => \N__16101\
        );

    \I__2518\ : IoInMux
    port map (
            O => \N__16122\,
            I => \N__16098\
        );

    \I__2517\ : IoInMux
    port map (
            O => \N__16121\,
            I => \N__16095\
        );

    \I__2516\ : IoInMux
    port map (
            O => \N__16120\,
            I => \N__16092\
        );

    \I__2515\ : IoSpan4Mux
    port map (
            O => \N__16117\,
            I => \N__16086\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__16114\,
            I => \N__16086\
        );

    \I__2513\ : IoInMux
    port map (
            O => \N__16113\,
            I => \N__16083\
        );

    \I__2512\ : IoInMux
    port map (
            O => \N__16112\,
            I => \N__16080\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__16109\,
            I => \N__16076\
        );

    \I__2510\ : IoSpan4Mux
    port map (
            O => \N__16104\,
            I => \N__16073\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__16101\,
            I => \N__16064\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__16098\,
            I => \N__16064\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__16095\,
            I => \N__16064\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__16092\,
            I => \N__16064\
        );

    \I__2505\ : IoInMux
    port map (
            O => \N__16091\,
            I => \N__16061\
        );

    \I__2504\ : IoSpan4Mux
    port map (
            O => \N__16086\,
            I => \N__16056\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__16083\,
            I => \N__16056\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__16080\,
            I => \N__16053\
        );

    \I__2501\ : IoInMux
    port map (
            O => \N__16079\,
            I => \N__16050\
        );

    \I__2500\ : IoSpan4Mux
    port map (
            O => \N__16076\,
            I => \N__16045\
        );

    \I__2499\ : IoSpan4Mux
    port map (
            O => \N__16073\,
            I => \N__16042\
        );

    \I__2498\ : IoSpan4Mux
    port map (
            O => \N__16064\,
            I => \N__16037\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__16061\,
            I => \N__16037\
        );

    \I__2496\ : IoSpan4Mux
    port map (
            O => \N__16056\,
            I => \N__16030\
        );

    \I__2495\ : IoSpan4Mux
    port map (
            O => \N__16053\,
            I => \N__16030\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__16050\,
            I => \N__16030\
        );

    \I__2493\ : IoInMux
    port map (
            O => \N__16049\,
            I => \N__16027\
        );

    \I__2492\ : IoInMux
    port map (
            O => \N__16048\,
            I => \N__16024\
        );

    \I__2491\ : IoSpan4Mux
    port map (
            O => \N__16045\,
            I => \N__16021\
        );

    \I__2490\ : IoSpan4Mux
    port map (
            O => \N__16042\,
            I => \N__16016\
        );

    \I__2489\ : IoSpan4Mux
    port map (
            O => \N__16037\,
            I => \N__16016\
        );

    \I__2488\ : IoSpan4Mux
    port map (
            O => \N__16030\,
            I => \N__16012\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__16027\,
            I => \N__16008\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__16024\,
            I => \N__16005\
        );

    \I__2485\ : Span4Mux_s2_h
    port map (
            O => \N__16021\,
            I => \N__16002\
        );

    \I__2484\ : Span4Mux_s1_h
    port map (
            O => \N__16016\,
            I => \N__15999\
        );

    \I__2483\ : IoInMux
    port map (
            O => \N__16015\,
            I => \N__15996\
        );

    \I__2482\ : Span4Mux_s2_v
    port map (
            O => \N__16012\,
            I => \N__15993\
        );

    \I__2481\ : IoInMux
    port map (
            O => \N__16011\,
            I => \N__15990\
        );

    \I__2480\ : Span12Mux_s6_h
    port map (
            O => \N__16008\,
            I => \N__15985\
        );

    \I__2479\ : Span12Mux_s4_v
    port map (
            O => \N__16005\,
            I => \N__15985\
        );

    \I__2478\ : Sp12to4
    port map (
            O => \N__16002\,
            I => \N__15982\
        );

    \I__2477\ : Sp12to4
    port map (
            O => \N__15999\,
            I => \N__15977\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__15996\,
            I => \N__15977\
        );

    \I__2475\ : Sp12to4
    port map (
            O => \N__15993\,
            I => \N__15972\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__15990\,
            I => \N__15972\
        );

    \I__2473\ : Span12Mux_v
    port map (
            O => \N__15985\,
            I => \N__15965\
        );

    \I__2472\ : Span12Mux_h
    port map (
            O => \N__15982\,
            I => \N__15965\
        );

    \I__2471\ : Span12Mux_s6_h
    port map (
            O => \N__15977\,
            I => \N__15965\
        );

    \I__2470\ : Span12Mux_s10_v
    port map (
            O => \N__15972\,
            I => \N__15962\
        );

    \I__2469\ : Odrv12
    port map (
            O => \N__15965\,
            I => dma_0_i
        );

    \I__2468\ : Odrv12
    port map (
            O => \N__15962\,
            I => dma_0_i
        );

    \I__2467\ : CEMux
    port map (
            O => \N__15957\,
            I => \N__15954\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__15954\,
            I => \N__15951\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__15951\,
            I => \N__15948\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__15948\,
            I => \N__15944\
        );

    \I__2463\ : CEMux
    port map (
            O => \N__15947\,
            I => \N__15941\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__15944\,
            I => \N_1430_0\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__15941\,
            I => \N_1430_0\
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__15936\,
            I => \this_vga_signals.N_1028_cascade_\
        );

    \I__2459\ : InMux
    port map (
            O => \N__15933\,
            I => \N__15929\
        );

    \I__2458\ : InMux
    port map (
            O => \N__15932\,
            I => \N__15926\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__15929\,
            I => \this_vga_signals.N_999\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__15926\,
            I => \this_vga_signals.N_999\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__15921\,
            I => \this_vga_signals.N_1004_cascade_\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__15918\,
            I => \N__15915\
        );

    \I__2453\ : InMux
    port map (
            O => \N__15915\,
            I => \N__15912\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__15912\,
            I => \this_vga_signals.N_1013\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__15909\,
            I => \this_vga_signals.N_1013_cascade_\
        );

    \I__2450\ : CascadeMux
    port map (
            O => \N__15906\,
            I => \this_vga_signals.N_105_mux_cascade_\
        );

    \I__2449\ : InMux
    port map (
            O => \N__15903\,
            I => \N__15899\
        );

    \I__2448\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15896\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__15899\,
            I => \this_vga_signals.N_113_mux\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__15896\,
            I => \this_vga_signals.N_113_mux\
        );

    \I__2445\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15888\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__15888\,
            I => \this_reset_cond.M_stage_qZ0Z_4\
        );

    \I__2443\ : InMux
    port map (
            O => \N__15885\,
            I => \N__15882\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__15882\,
            I => \this_reset_cond.M_stage_qZ0Z_5\
        );

    \I__2441\ : InMux
    port map (
            O => \N__15879\,
            I => \N__15876\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__15876\,
            I => \N__15873\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__15873\,
            I => \N__15869\
        );

    \I__2438\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15866\
        );

    \I__2437\ : Span4Mux_v
    port map (
            O => \N__15869\,
            I => \N__15862\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__15866\,
            I => \N__15859\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__15865\,
            I => \N__15856\
        );

    \I__2434\ : Span4Mux_v
    port map (
            O => \N__15862\,
            I => \N__15851\
        );

    \I__2433\ : Span4Mux_v
    port map (
            O => \N__15859\,
            I => \N__15851\
        );

    \I__2432\ : InMux
    port map (
            O => \N__15856\,
            I => \N__15847\
        );

    \I__2431\ : Sp12to4
    port map (
            O => \N__15851\,
            I => \N__15844\
        );

    \I__2430\ : InMux
    port map (
            O => \N__15850\,
            I => \N__15841\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__15847\,
            I => \N__15838\
        );

    \I__2428\ : Span12Mux_h
    port map (
            O => \N__15844\,
            I => \N__15835\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__15841\,
            I => \N__15832\
        );

    \I__2426\ : Span4Mux_v
    port map (
            O => \N__15838\,
            I => \N__15829\
        );

    \I__2425\ : Odrv12
    port map (
            O => \N__15835\,
            I => this_vga_signals_vvisibility
        );

    \I__2424\ : Odrv4
    port map (
            O => \N__15832\,
            I => this_vga_signals_vvisibility
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__15829\,
            I => this_vga_signals_vvisibility
        );

    \I__2422\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15818\
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__15821\,
            I => \N__15811\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__15818\,
            I => \N__15806\
        );

    \I__2419\ : InMux
    port map (
            O => \N__15817\,
            I => \N__15803\
        );

    \I__2418\ : InMux
    port map (
            O => \N__15816\,
            I => \N__15800\
        );

    \I__2417\ : InMux
    port map (
            O => \N__15815\,
            I => \N__15797\
        );

    \I__2416\ : InMux
    port map (
            O => \N__15814\,
            I => \N__15790\
        );

    \I__2415\ : InMux
    port map (
            O => \N__15811\,
            I => \N__15790\
        );

    \I__2414\ : InMux
    port map (
            O => \N__15810\,
            I => \N__15790\
        );

    \I__2413\ : IoInMux
    port map (
            O => \N__15809\,
            I => \N__15787\
        );

    \I__2412\ : Span4Mux_v
    port map (
            O => \N__15806\,
            I => \N__15782\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__15803\,
            I => \N__15782\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__15800\,
            I => \N__15779\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__15797\,
            I => \N__15774\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__15790\,
            I => \N__15774\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__15787\,
            I => \N__15768\
        );

    \I__2406\ : Span4Mux_h
    port map (
            O => \N__15782\,
            I => \N__15765\
        );

    \I__2405\ : Span4Mux_v
    port map (
            O => \N__15779\,
            I => \N__15760\
        );

    \I__2404\ : Span4Mux_v
    port map (
            O => \N__15774\,
            I => \N__15760\
        );

    \I__2403\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15757\
        );

    \I__2402\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15754\
        );

    \I__2401\ : InMux
    port map (
            O => \N__15771\,
            I => \N__15751\
        );

    \I__2400\ : Span4Mux_s3_v
    port map (
            O => \N__15768\,
            I => \N__15748\
        );

    \I__2399\ : Span4Mux_v
    port map (
            O => \N__15765\,
            I => \N__15745\
        );

    \I__2398\ : Span4Mux_h
    port map (
            O => \N__15760\,
            I => \N__15736\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__15757\,
            I => \N__15736\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__15754\,
            I => \N__15736\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__15751\,
            I => \N__15736\
        );

    \I__2394\ : Span4Mux_v
    port map (
            O => \N__15748\,
            I => \N__15733\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__15745\,
            I => \M_this_reset_cond_out_0\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__15736\,
            I => \M_this_reset_cond_out_0\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__15733\,
            I => \M_this_reset_cond_out_0\
        );

    \I__2390\ : InMux
    port map (
            O => \N__15726\,
            I => \N__15723\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__15723\,
            I => \N__15720\
        );

    \I__2388\ : Span4Mux_h
    port map (
            O => \N__15720\,
            I => \N__15717\
        );

    \I__2387\ : Odrv4
    port map (
            O => \N__15717\,
            I => \this_ppu.un3_sprites_addr_cry_2_c_RNIVRCZ0Z8\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__15714\,
            I => \N__15711\
        );

    \I__2385\ : CascadeBuf
    port map (
            O => \N__15711\,
            I => \N__15708\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__15708\,
            I => \N__15705\
        );

    \I__2383\ : CascadeBuf
    port map (
            O => \N__15705\,
            I => \N__15702\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__15702\,
            I => \N__15699\
        );

    \I__2381\ : CascadeBuf
    port map (
            O => \N__15699\,
            I => \N__15696\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__15696\,
            I => \N__15693\
        );

    \I__2379\ : CascadeBuf
    port map (
            O => \N__15693\,
            I => \N__15690\
        );

    \I__2378\ : CascadeMux
    port map (
            O => \N__15690\,
            I => \N__15687\
        );

    \I__2377\ : CascadeBuf
    port map (
            O => \N__15687\,
            I => \N__15684\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__15684\,
            I => \N__15681\
        );

    \I__2375\ : CascadeBuf
    port map (
            O => \N__15681\,
            I => \N__15678\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__15678\,
            I => \N__15675\
        );

    \I__2373\ : CascadeBuf
    port map (
            O => \N__15675\,
            I => \N__15672\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__15672\,
            I => \N__15669\
        );

    \I__2371\ : CascadeBuf
    port map (
            O => \N__15669\,
            I => \N__15666\
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__15666\,
            I => \N__15663\
        );

    \I__2369\ : CascadeBuf
    port map (
            O => \N__15663\,
            I => \N__15660\
        );

    \I__2368\ : CascadeMux
    port map (
            O => \N__15660\,
            I => \N__15657\
        );

    \I__2367\ : CascadeBuf
    port map (
            O => \N__15657\,
            I => \N__15654\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__15654\,
            I => \N__15651\
        );

    \I__2365\ : CascadeBuf
    port map (
            O => \N__15651\,
            I => \N__15648\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__15648\,
            I => \N__15645\
        );

    \I__2363\ : CascadeBuf
    port map (
            O => \N__15645\,
            I => \N__15642\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__15642\,
            I => \N__15639\
        );

    \I__2361\ : CascadeBuf
    port map (
            O => \N__15639\,
            I => \N__15636\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__15636\,
            I => \N__15633\
        );

    \I__2359\ : CascadeBuf
    port map (
            O => \N__15633\,
            I => \N__15630\
        );

    \I__2358\ : CascadeMux
    port map (
            O => \N__15630\,
            I => \N__15627\
        );

    \I__2357\ : CascadeBuf
    port map (
            O => \N__15627\,
            I => \N__15624\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__15624\,
            I => \N__15621\
        );

    \I__2355\ : InMux
    port map (
            O => \N__15621\,
            I => \N__15618\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__15618\,
            I => \N__15615\
        );

    \I__2353\ : Span12Mux_h
    port map (
            O => \N__15615\,
            I => \N__15612\
        );

    \I__2352\ : Span12Mux_v
    port map (
            O => \N__15612\,
            I => \N__15609\
        );

    \I__2351\ : Odrv12
    port map (
            O => \N__15609\,
            I => \M_this_ppu_sprites_addr_3\
        );

    \I__2350\ : InMux
    port map (
            O => \N__15606\,
            I => \N__15603\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__15603\,
            I => \N__15600\
        );

    \I__2348\ : Span4Mux_h
    port map (
            O => \N__15600\,
            I => \N__15597\
        );

    \I__2347\ : Span4Mux_h
    port map (
            O => \N__15597\,
            I => \N__15594\
        );

    \I__2346\ : Odrv4
    port map (
            O => \N__15594\,
            I => \this_oam_ram.M_this_oam_ram_read_data_9\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__15591\,
            I => \N__15588\
        );

    \I__2344\ : InMux
    port map (
            O => \N__15588\,
            I => \N__15585\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__15585\,
            I => \N__15582\
        );

    \I__2342\ : Span4Mux_v
    port map (
            O => \N__15582\,
            I => \N__15579\
        );

    \I__2341\ : Span4Mux_h
    port map (
            O => \N__15579\,
            I => \N__15576\
        );

    \I__2340\ : Span4Mux_h
    port map (
            O => \N__15576\,
            I => \N__15573\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__15573\,
            I => \M_this_map_ram_read_data_3\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__15570\,
            I => \N__15567\
        );

    \I__2337\ : CascadeBuf
    port map (
            O => \N__15567\,
            I => \N__15564\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__15564\,
            I => \N__15561\
        );

    \I__2335\ : CascadeBuf
    port map (
            O => \N__15561\,
            I => \N__15558\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__15558\,
            I => \N__15555\
        );

    \I__2333\ : CascadeBuf
    port map (
            O => \N__15555\,
            I => \N__15552\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__15552\,
            I => \N__15549\
        );

    \I__2331\ : CascadeBuf
    port map (
            O => \N__15549\,
            I => \N__15546\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__15546\,
            I => \N__15543\
        );

    \I__2329\ : CascadeBuf
    port map (
            O => \N__15543\,
            I => \N__15540\
        );

    \I__2328\ : CascadeMux
    port map (
            O => \N__15540\,
            I => \N__15537\
        );

    \I__2327\ : CascadeBuf
    port map (
            O => \N__15537\,
            I => \N__15534\
        );

    \I__2326\ : CascadeMux
    port map (
            O => \N__15534\,
            I => \N__15531\
        );

    \I__2325\ : CascadeBuf
    port map (
            O => \N__15531\,
            I => \N__15528\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__15528\,
            I => \N__15525\
        );

    \I__2323\ : CascadeBuf
    port map (
            O => \N__15525\,
            I => \N__15522\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__15522\,
            I => \N__15519\
        );

    \I__2321\ : CascadeBuf
    port map (
            O => \N__15519\,
            I => \N__15516\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__15516\,
            I => \N__15513\
        );

    \I__2319\ : CascadeBuf
    port map (
            O => \N__15513\,
            I => \N__15510\
        );

    \I__2318\ : CascadeMux
    port map (
            O => \N__15510\,
            I => \N__15507\
        );

    \I__2317\ : CascadeBuf
    port map (
            O => \N__15507\,
            I => \N__15504\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__15504\,
            I => \N__15501\
        );

    \I__2315\ : CascadeBuf
    port map (
            O => \N__15501\,
            I => \N__15498\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__15498\,
            I => \N__15495\
        );

    \I__2313\ : CascadeBuf
    port map (
            O => \N__15495\,
            I => \N__15492\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__15492\,
            I => \N__15489\
        );

    \I__2311\ : CascadeBuf
    port map (
            O => \N__15489\,
            I => \N__15486\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__15486\,
            I => \N__15483\
        );

    \I__2309\ : CascadeBuf
    port map (
            O => \N__15483\,
            I => \N__15480\
        );

    \I__2308\ : CascadeMux
    port map (
            O => \N__15480\,
            I => \N__15477\
        );

    \I__2307\ : InMux
    port map (
            O => \N__15477\,
            I => \N__15474\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__15474\,
            I => \N__15471\
        );

    \I__2305\ : Span4Mux_h
    port map (
            O => \N__15471\,
            I => \N__15468\
        );

    \I__2304\ : Sp12to4
    port map (
            O => \N__15468\,
            I => \N__15465\
        );

    \I__2303\ : Span12Mux_s6_v
    port map (
            O => \N__15465\,
            I => \N__15462\
        );

    \I__2302\ : Span12Mux_h
    port map (
            O => \N__15462\,
            I => \N__15459\
        );

    \I__2301\ : Odrv12
    port map (
            O => \N__15459\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__15456\,
            I => \N__15453\
        );

    \I__2299\ : InMux
    port map (
            O => \N__15453\,
            I => \N__15447\
        );

    \I__2298\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15447\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__15447\,
            I => \this_ppu.M_state_d_0_sqmuxa_1\
        );

    \I__2296\ : InMux
    port map (
            O => \N__15444\,
            I => \N__15441\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__15441\,
            I => \N__15438\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__15438\,
            I => \this_ppu.M_count_q_RNO_0Z0Z_7\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__15435\,
            I => \N__15431\
        );

    \I__2292\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15428\
        );

    \I__2291\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15425\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__15428\,
            I => \N__15420\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__15425\,
            I => \N__15420\
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__15420\,
            I => \this_ppu.M_count_qZ0Z_7\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__15417\,
            I => \N__15414\
        );

    \I__2286\ : InMux
    port map (
            O => \N__15414\,
            I => \N__15411\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__15411\,
            I => \this_vga_signals.N_129_mux\
        );

    \I__2284\ : InMux
    port map (
            O => \N__15408\,
            I => \N__15405\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__15405\,
            I => \this_vga_signals.N_1028\
        );

    \I__2282\ : InMux
    port map (
            O => \N__15402\,
            I => \N__15399\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__15399\,
            I => \M_this_data_tmp_qZ0Z_10\
        );

    \I__2280\ : InMux
    port map (
            O => \N__15396\,
            I => \N__15393\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__15393\,
            I => \N__15390\
        );

    \I__2278\ : Span4Mux_h
    port map (
            O => \N__15390\,
            I => \N__15387\
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__15387\,
            I => \M_this_data_tmp_qZ0Z_17\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__15384\,
            I => \N__15381\
        );

    \I__2275\ : InMux
    port map (
            O => \N__15381\,
            I => \N__15378\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__15378\,
            I => \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\
        );

    \I__2273\ : InMux
    port map (
            O => \N__15375\,
            I => \N__15370\
        );

    \I__2272\ : InMux
    port map (
            O => \N__15374\,
            I => \N__15367\
        );

    \I__2271\ : InMux
    port map (
            O => \N__15373\,
            I => \N__15364\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__15370\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__15367\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__15364\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__2267\ : InMux
    port map (
            O => \N__15357\,
            I => \N__15352\
        );

    \I__2266\ : InMux
    port map (
            O => \N__15356\,
            I => \N__15349\
        );

    \I__2265\ : InMux
    port map (
            O => \N__15355\,
            I => \N__15346\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__15352\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__15349\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__15346\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__15339\,
            I => \N__15336\
        );

    \I__2260\ : InMux
    port map (
            O => \N__15336\,
            I => \N__15333\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__15333\,
            I => \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__15330\,
            I => \N__15327\
        );

    \I__2257\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15322\
        );

    \I__2256\ : InMux
    port map (
            O => \N__15326\,
            I => \N__15317\
        );

    \I__2255\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15317\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__15322\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__15317\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__2252\ : InMux
    port map (
            O => \N__15312\,
            I => \N__15309\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__15309\,
            I => \N__15306\
        );

    \I__2250\ : Span4Mux_h
    port map (
            O => \N__15306\,
            I => \N__15303\
        );

    \I__2249\ : Span4Mux_v
    port map (
            O => \N__15303\,
            I => \N__15300\
        );

    \I__2248\ : Span4Mux_h
    port map (
            O => \N__15300\,
            I => \N__15297\
        );

    \I__2247\ : Odrv4
    port map (
            O => \N__15297\,
            I => \M_this_map_ram_read_data_2\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__15294\,
            I => \this_ppu.un10_sprites_addr_axb_0_cascade_\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__15291\,
            I => \N__15288\
        );

    \I__2244\ : CascadeBuf
    port map (
            O => \N__15288\,
            I => \N__15285\
        );

    \I__2243\ : CascadeMux
    port map (
            O => \N__15285\,
            I => \N__15282\
        );

    \I__2242\ : CascadeBuf
    port map (
            O => \N__15282\,
            I => \N__15279\
        );

    \I__2241\ : CascadeMux
    port map (
            O => \N__15279\,
            I => \N__15276\
        );

    \I__2240\ : CascadeBuf
    port map (
            O => \N__15276\,
            I => \N__15273\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__15273\,
            I => \N__15270\
        );

    \I__2238\ : CascadeBuf
    port map (
            O => \N__15270\,
            I => \N__15267\
        );

    \I__2237\ : CascadeMux
    port map (
            O => \N__15267\,
            I => \N__15264\
        );

    \I__2236\ : CascadeBuf
    port map (
            O => \N__15264\,
            I => \N__15261\
        );

    \I__2235\ : CascadeMux
    port map (
            O => \N__15261\,
            I => \N__15258\
        );

    \I__2234\ : CascadeBuf
    port map (
            O => \N__15258\,
            I => \N__15255\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__15255\,
            I => \N__15252\
        );

    \I__2232\ : CascadeBuf
    port map (
            O => \N__15252\,
            I => \N__15249\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__15249\,
            I => \N__15246\
        );

    \I__2230\ : CascadeBuf
    port map (
            O => \N__15246\,
            I => \N__15243\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__15243\,
            I => \N__15240\
        );

    \I__2228\ : CascadeBuf
    port map (
            O => \N__15240\,
            I => \N__15237\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__15237\,
            I => \N__15234\
        );

    \I__2226\ : CascadeBuf
    port map (
            O => \N__15234\,
            I => \N__15231\
        );

    \I__2225\ : CascadeMux
    port map (
            O => \N__15231\,
            I => \N__15228\
        );

    \I__2224\ : CascadeBuf
    port map (
            O => \N__15228\,
            I => \N__15225\
        );

    \I__2223\ : CascadeMux
    port map (
            O => \N__15225\,
            I => \N__15222\
        );

    \I__2222\ : CascadeBuf
    port map (
            O => \N__15222\,
            I => \N__15219\
        );

    \I__2221\ : CascadeMux
    port map (
            O => \N__15219\,
            I => \N__15216\
        );

    \I__2220\ : CascadeBuf
    port map (
            O => \N__15216\,
            I => \N__15213\
        );

    \I__2219\ : CascadeMux
    port map (
            O => \N__15213\,
            I => \N__15210\
        );

    \I__2218\ : CascadeBuf
    port map (
            O => \N__15210\,
            I => \N__15207\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__15207\,
            I => \N__15204\
        );

    \I__2216\ : CascadeBuf
    port map (
            O => \N__15204\,
            I => \N__15201\
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__15201\,
            I => \N__15198\
        );

    \I__2214\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15195\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__15195\,
            I => \N__15192\
        );

    \I__2212\ : Span4Mux_h
    port map (
            O => \N__15192\,
            I => \N__15189\
        );

    \I__2211\ : Span4Mux_h
    port map (
            O => \N__15189\,
            I => \N__15186\
        );

    \I__2210\ : Span4Mux_v
    port map (
            O => \N__15186\,
            I => \N__15183\
        );

    \I__2209\ : Span4Mux_v
    port map (
            O => \N__15183\,
            I => \N__15180\
        );

    \I__2208\ : Span4Mux_v
    port map (
            O => \N__15180\,
            I => \N__15177\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__15177\,
            I => \M_this_ppu_sprites_addr_8\
        );

    \I__2206\ : InMux
    port map (
            O => \N__15174\,
            I => \N__15166\
        );

    \I__2205\ : InMux
    port map (
            O => \N__15173\,
            I => \N__15166\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__15172\,
            I => \N__15162\
        );

    \I__2203\ : InMux
    port map (
            O => \N__15171\,
            I => \N__15157\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__15166\,
            I => \N__15154\
        );

    \I__2201\ : InMux
    port map (
            O => \N__15165\,
            I => \N__15151\
        );

    \I__2200\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15144\
        );

    \I__2199\ : InMux
    port map (
            O => \N__15161\,
            I => \N__15144\
        );

    \I__2198\ : InMux
    port map (
            O => \N__15160\,
            I => \N__15144\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__15157\,
            I => \N__15141\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__15154\,
            I => \this_ppu.un10_0\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__15151\,
            I => \this_ppu.un10_0\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__15144\,
            I => \this_ppu.un10_0\
        );

    \I__2193\ : Odrv12
    port map (
            O => \N__15141\,
            I => \this_ppu.un10_0\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__15132\,
            I => \N__15129\
        );

    \I__2191\ : InMux
    port map (
            O => \N__15129\,
            I => \N__15126\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__15126\,
            I => \N__15123\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__15123\,
            I => \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\
        );

    \I__2188\ : InMux
    port map (
            O => \N__15120\,
            I => \N__15112\
        );

    \I__2187\ : InMux
    port map (
            O => \N__15119\,
            I => \N__15107\
        );

    \I__2186\ : InMux
    port map (
            O => \N__15118\,
            I => \N__15107\
        );

    \I__2185\ : InMux
    port map (
            O => \N__15117\,
            I => \N__15104\
        );

    \I__2184\ : InMux
    port map (
            O => \N__15116\,
            I => \N__15099\
        );

    \I__2183\ : InMux
    port map (
            O => \N__15115\,
            I => \N__15099\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__15112\,
            I => \N__15096\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__15107\,
            I => \this_ppu.N_1456_0\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__15104\,
            I => \this_ppu.N_1456_0\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__15099\,
            I => \this_ppu.N_1456_0\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__15096\,
            I => \this_ppu.N_1456_0\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__15087\,
            I => \N__15082\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__15086\,
            I => \N__15079\
        );

    \I__2175\ : InMux
    port map (
            O => \N__15085\,
            I => \N__15076\
        );

    \I__2174\ : InMux
    port map (
            O => \N__15082\,
            I => \N__15073\
        );

    \I__2173\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15070\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__15076\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__15073\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__15070\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__2169\ : InMux
    port map (
            O => \N__15063\,
            I => \N__15060\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__15060\,
            I => \N__15057\
        );

    \I__2167\ : Odrv12
    port map (
            O => \N__15057\,
            I => \this_reset_cond.M_stage_qZ0Z_3\
        );

    \I__2166\ : InMux
    port map (
            O => \N__15054\,
            I => \N__15046\
        );

    \I__2165\ : InMux
    port map (
            O => \N__15053\,
            I => \N__15046\
        );

    \I__2164\ : InMux
    port map (
            O => \N__15052\,
            I => \N__15041\
        );

    \I__2163\ : InMux
    port map (
            O => \N__15051\,
            I => \N__15041\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__15046\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__15041\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__15036\,
            I => \this_vga_signals.i21_mux_cascade_\
        );

    \I__2159\ : InMux
    port map (
            O => \N__15033\,
            I => \N__15027\
        );

    \I__2158\ : InMux
    port map (
            O => \N__15032\,
            I => \N__15024\
        );

    \I__2157\ : InMux
    port map (
            O => \N__15031\,
            I => \N__15019\
        );

    \I__2156\ : InMux
    port map (
            O => \N__15030\,
            I => \N__15019\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__15027\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__15024\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__15019\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__2152\ : InMux
    port map (
            O => \N__15012\,
            I => \N__15009\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__15009\,
            I => \N__15006\
        );

    \I__2150\ : Span4Mux_h
    port map (
            O => \N__15006\,
            I => \N__15003\
        );

    \I__2149\ : Span4Mux_h
    port map (
            O => \N__15003\,
            I => \N__15000\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__15000\,
            I => \N_817_0\
        );

    \I__2147\ : InMux
    port map (
            O => \N__14997\,
            I => \N__14994\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__14994\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__2145\ : InMux
    port map (
            O => \N__14991\,
            I => \N__14988\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__14988\,
            I => \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__14985\,
            I => \N__14982\
        );

    \I__2142\ : InMux
    port map (
            O => \N__14982\,
            I => \N__14979\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__14979\,
            I => \N__14976\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__14976\,
            I => \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\
        );

    \I__2139\ : InMux
    port map (
            O => \N__14973\,
            I => \N__14968\
        );

    \I__2138\ : InMux
    port map (
            O => \N__14972\,
            I => \N__14965\
        );

    \I__2137\ : InMux
    port map (
            O => \N__14971\,
            I => \N__14962\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__14968\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__14965\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__14962\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__14955\,
            I => \N__14952\
        );

    \I__2132\ : InMux
    port map (
            O => \N__14952\,
            I => \N__14947\
        );

    \I__2131\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14942\
        );

    \I__2130\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14942\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__14947\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__14942\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__2127\ : InMux
    port map (
            O => \N__14937\,
            I => \N__14932\
        );

    \I__2126\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14927\
        );

    \I__2125\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14927\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__14932\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__14927\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__2122\ : SRMux
    port map (
            O => \N__14922\,
            I => \N__14919\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__14919\,
            I => \N__14915\
        );

    \I__2120\ : SRMux
    port map (
            O => \N__14918\,
            I => \N__14912\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__14915\,
            I => \N__14909\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__14912\,
            I => \N__14906\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__14909\,
            I => \this_ppu.M_state_q_RNIE20V4Z0Z_0\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__14906\,
            I => \this_ppu.M_state_q_RNIE20V4Z0Z_0\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__14901\,
            I => \M_this_vga_signals_line_clk_0_cascade_\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__14898\,
            I => \this_ppu.M_state_d_0_sqmuxa_cascade_\
        );

    \I__2113\ : CascadeMux
    port map (
            O => \N__14895\,
            I => \this_vga_signals.N_1000_cascade_\
        );

    \I__2112\ : InMux
    port map (
            O => \N__14892\,
            I => \this_ppu.un1_M_count_q_1_cry_1_s1\
        );

    \I__2111\ : InMux
    port map (
            O => \N__14889\,
            I => \this_ppu.un1_M_count_q_1_cry_2_s1\
        );

    \I__2110\ : InMux
    port map (
            O => \N__14886\,
            I => \this_ppu.un1_M_count_q_1_cry_3_s1\
        );

    \I__2109\ : InMux
    port map (
            O => \N__14883\,
            I => \this_ppu.un1_M_count_q_1_cry_4_s1\
        );

    \I__2108\ : InMux
    port map (
            O => \N__14880\,
            I => \this_ppu.un1_M_count_q_1_cry_5_s1\
        );

    \I__2107\ : InMux
    port map (
            O => \N__14877\,
            I => \this_ppu.un1_M_count_q_1_cry_6_s1\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__14874\,
            I => \this_ppu.M_state_d_0_sqmuxa_1_cascade_\
        );

    \I__2105\ : InMux
    port map (
            O => \N__14871\,
            I => \N__14868\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__14868\,
            I => \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__14865\,
            I => \this_ppu.N_1456_0_cascade_\
        );

    \I__2102\ : CEMux
    port map (
            O => \N__14862\,
            I => \N__14859\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__14859\,
            I => \N__14856\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__14856\,
            I => \this_vga_signals.N_1090_1\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__14853\,
            I => \N__14850\
        );

    \I__2098\ : InMux
    port map (
            O => \N__14850\,
            I => \N__14845\
        );

    \I__2097\ : InMux
    port map (
            O => \N__14849\,
            I => \N__14842\
        );

    \I__2096\ : InMux
    port map (
            O => \N__14848\,
            I => \N__14839\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__14845\,
            I => \N__14834\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__14842\,
            I => \N__14829\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__14839\,
            I => \N__14829\
        );

    \I__2092\ : InMux
    port map (
            O => \N__14838\,
            I => \N__14823\
        );

    \I__2091\ : InMux
    port map (
            O => \N__14837\,
            I => \N__14823\
        );

    \I__2090\ : Span4Mux_v
    port map (
            O => \N__14834\,
            I => \N__14818\
        );

    \I__2089\ : Span4Mux_v
    port map (
            O => \N__14829\,
            I => \N__14818\
        );

    \I__2088\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14815\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__14823\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__14818\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__14815\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__14808\,
            I => \N__14803\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__14807\,
            I => \N__14800\
        );

    \I__2082\ : InMux
    port map (
            O => \N__14806\,
            I => \N__14795\
        );

    \I__2081\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14792\
        );

    \I__2080\ : InMux
    port map (
            O => \N__14800\,
            I => \N__14789\
        );

    \I__2079\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14784\
        );

    \I__2078\ : InMux
    port map (
            O => \N__14798\,
            I => \N__14784\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__14795\,
            I => \N__14776\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__14792\,
            I => \N__14776\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__14789\,
            I => \N__14776\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__14784\,
            I => \N__14773\
        );

    \I__2073\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14769\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__14776\,
            I => \N__14766\
        );

    \I__2071\ : Span4Mux_h
    port map (
            O => \N__14773\,
            I => \N__14763\
        );

    \I__2070\ : InMux
    port map (
            O => \N__14772\,
            I => \N__14760\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__14769\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__14766\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__14763\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__14760\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2065\ : SRMux
    port map (
            O => \N__14751\,
            I => \N__14746\
        );

    \I__2064\ : SRMux
    port map (
            O => \N__14750\,
            I => \N__14743\
        );

    \I__2063\ : SRMux
    port map (
            O => \N__14749\,
            I => \N__14739\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__14746\,
            I => \N__14736\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__14743\,
            I => \N__14733\
        );

    \I__2060\ : InMux
    port map (
            O => \N__14742\,
            I => \N__14730\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__14739\,
            I => \G_464\
        );

    \I__2058\ : Odrv12
    port map (
            O => \N__14736\,
            I => \G_464\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__14733\,
            I => \G_464\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__14730\,
            I => \G_464\
        );

    \I__2055\ : InMux
    port map (
            O => \N__14721\,
            I => \N__14718\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__14718\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__2053\ : InMux
    port map (
            O => \N__14715\,
            I => \N__14712\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__14712\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__2051\ : InMux
    port map (
            O => \N__14709\,
            I => \N__14706\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__14706\,
            I => \N__14703\
        );

    \I__2049\ : Span4Mux_h
    port map (
            O => \N__14703\,
            I => \N__14700\
        );

    \I__2048\ : Odrv4
    port map (
            O => \N__14700\,
            I => \M_this_oam_ram_write_data_10\
        );

    \I__2047\ : InMux
    port map (
            O => \N__14697\,
            I => \this_ppu.un1_M_count_q_1_cry_0_s1\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__14694\,
            I => \N__14691\
        );

    \I__2045\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14688\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__14688\,
            I => \this_ppu.M_state_qc_1_3\
        );

    \I__2043\ : InMux
    port map (
            O => \N__14685\,
            I => \N__14682\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__14682\,
            I => \N__14679\
        );

    \I__2041\ : Span4Mux_h
    port map (
            O => \N__14679\,
            I => \N__14676\
        );

    \I__2040\ : Sp12to4
    port map (
            O => \N__14676\,
            I => \N__14673\
        );

    \I__2039\ : Span12Mux_v
    port map (
            O => \N__14673\,
            I => \N__14669\
        );

    \I__2038\ : InMux
    port map (
            O => \N__14672\,
            I => \N__14666\
        );

    \I__2037\ : Odrv12
    port map (
            O => \N__14669\,
            I => \M_this_ppu_vram_data_0\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__14666\,
            I => \M_this_ppu_vram_data_0\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__14661\,
            I => \this_ppu.M_state_qc_1_1_cascade_\
        );

    \I__2034\ : InMux
    port map (
            O => \N__14658\,
            I => \N__14652\
        );

    \I__2033\ : InMux
    port map (
            O => \N__14657\,
            I => \N__14652\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__14652\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__14649\,
            I => \N__14644\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__14648\,
            I => \N__14641\
        );

    \I__2029\ : InMux
    port map (
            O => \N__14647\,
            I => \N__14635\
        );

    \I__2028\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14635\
        );

    \I__2027\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14632\
        );

    \I__2026\ : InMux
    port map (
            O => \N__14640\,
            I => \N__14629\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__14635\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__14632\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__14629\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__14622\,
            I => \N__14619\
        );

    \I__2021\ : InMux
    port map (
            O => \N__14619\,
            I => \N__14614\
        );

    \I__2020\ : InMux
    port map (
            O => \N__14618\,
            I => \N__14608\
        );

    \I__2019\ : InMux
    port map (
            O => \N__14617\,
            I => \N__14604\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__14614\,
            I => \N__14601\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__14613\,
            I => \N__14596\
        );

    \I__2016\ : InMux
    port map (
            O => \N__14612\,
            I => \N__14593\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__14611\,
            I => \N__14590\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__14608\,
            I => \N__14587\
        );

    \I__2013\ : InMux
    port map (
            O => \N__14607\,
            I => \N__14584\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__14604\,
            I => \N__14579\
        );

    \I__2011\ : Span4Mux_v
    port map (
            O => \N__14601\,
            I => \N__14579\
        );

    \I__2010\ : InMux
    port map (
            O => \N__14600\,
            I => \N__14572\
        );

    \I__2009\ : InMux
    port map (
            O => \N__14599\,
            I => \N__14572\
        );

    \I__2008\ : InMux
    port map (
            O => \N__14596\,
            I => \N__14572\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__14593\,
            I => \N__14569\
        );

    \I__2006\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14566\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__14587\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__14584\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__14579\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__14572\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2001\ : Odrv4
    port map (
            O => \N__14569\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__14566\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1999\ : InMux
    port map (
            O => \N__14553\,
            I => \N__14542\
        );

    \I__1998\ : InMux
    port map (
            O => \N__14552\,
            I => \N__14542\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__14551\,
            I => \N__14539\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__14550\,
            I => \N__14536\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__14549\,
            I => \N__14532\
        );

    \I__1994\ : InMux
    port map (
            O => \N__14548\,
            I => \N__14529\
        );

    \I__1993\ : InMux
    port map (
            O => \N__14547\,
            I => \N__14525\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__14542\,
            I => \N__14522\
        );

    \I__1991\ : InMux
    port map (
            O => \N__14539\,
            I => \N__14512\
        );

    \I__1990\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14512\
        );

    \I__1989\ : InMux
    port map (
            O => \N__14535\,
            I => \N__14512\
        );

    \I__1988\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14512\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__14529\,
            I => \N__14509\
        );

    \I__1986\ : InMux
    port map (
            O => \N__14528\,
            I => \N__14506\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__14525\,
            I => \N__14503\
        );

    \I__1984\ : Span4Mux_h
    port map (
            O => \N__14522\,
            I => \N__14500\
        );

    \I__1983\ : InMux
    port map (
            O => \N__14521\,
            I => \N__14497\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__14512\,
            I => \N__14494\
        );

    \I__1981\ : Odrv4
    port map (
            O => \N__14509\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__14506\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__14503\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__14500\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__14497\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1976\ : Odrv4
    port map (
            O => \N__14494\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1975\ : InMux
    port map (
            O => \N__14481\,
            I => \N__14463\
        );

    \I__1974\ : InMux
    port map (
            O => \N__14480\,
            I => \N__14463\
        );

    \I__1973\ : InMux
    port map (
            O => \N__14479\,
            I => \N__14463\
        );

    \I__1972\ : InMux
    port map (
            O => \N__14478\,
            I => \N__14463\
        );

    \I__1971\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14458\
        );

    \I__1970\ : InMux
    port map (
            O => \N__14476\,
            I => \N__14458\
        );

    \I__1969\ : InMux
    port map (
            O => \N__14475\,
            I => \N__14455\
        );

    \I__1968\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14451\
        );

    \I__1967\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14448\
        );

    \I__1966\ : InMux
    port map (
            O => \N__14472\,
            I => \N__14445\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__14463\,
            I => \N__14442\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__14458\,
            I => \N__14437\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__14455\,
            I => \N__14437\
        );

    \I__1962\ : InMux
    port map (
            O => \N__14454\,
            I => \N__14434\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__14451\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__14448\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__14445\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__14442\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__14437\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__14434\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1955\ : InMux
    port map (
            O => \N__14421\,
            I => \N__14413\
        );

    \I__1954\ : InMux
    port map (
            O => \N__14420\,
            I => \N__14413\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__14419\,
            I => \N__14407\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__14418\,
            I => \N__14403\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__14413\,
            I => \N__14398\
        );

    \I__1950\ : InMux
    port map (
            O => \N__14412\,
            I => \N__14395\
        );

    \I__1949\ : InMux
    port map (
            O => \N__14411\,
            I => \N__14392\
        );

    \I__1948\ : InMux
    port map (
            O => \N__14410\,
            I => \N__14387\
        );

    \I__1947\ : InMux
    port map (
            O => \N__14407\,
            I => \N__14387\
        );

    \I__1946\ : InMux
    port map (
            O => \N__14406\,
            I => \N__14378\
        );

    \I__1945\ : InMux
    port map (
            O => \N__14403\,
            I => \N__14378\
        );

    \I__1944\ : InMux
    port map (
            O => \N__14402\,
            I => \N__14378\
        );

    \I__1943\ : InMux
    port map (
            O => \N__14401\,
            I => \N__14378\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__14398\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__14395\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__14392\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__14387\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__14378\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__14367\,
            I => \this_vga_signals.N_18_0_cascade_\
        );

    \I__1936\ : InMux
    port map (
            O => \N__14364\,
            I => \N__14360\
        );

    \I__1935\ : InMux
    port map (
            O => \N__14363\,
            I => \N__14356\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__14360\,
            I => \N__14353\
        );

    \I__1933\ : InMux
    port map (
            O => \N__14359\,
            I => \N__14343\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__14356\,
            I => \N__14338\
        );

    \I__1931\ : Span4Mux_v
    port map (
            O => \N__14353\,
            I => \N__14338\
        );

    \I__1930\ : InMux
    port map (
            O => \N__14352\,
            I => \N__14335\
        );

    \I__1929\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14332\
        );

    \I__1928\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14321\
        );

    \I__1927\ : InMux
    port map (
            O => \N__14349\,
            I => \N__14321\
        );

    \I__1926\ : InMux
    port map (
            O => \N__14348\,
            I => \N__14321\
        );

    \I__1925\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14321\
        );

    \I__1924\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14321\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__14343\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__14338\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__14335\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__14332\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__14321\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1918\ : CascadeMux
    port map (
            O => \N__14310\,
            I => \N__14306\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__14309\,
            I => \N__14302\
        );

    \I__1916\ : InMux
    port map (
            O => \N__14306\,
            I => \N__14299\
        );

    \I__1915\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14296\
        );

    \I__1914\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14293\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__14299\,
            I => \N__14287\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__14296\,
            I => \N__14282\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__14293\,
            I => \N__14282\
        );

    \I__1910\ : InMux
    port map (
            O => \N__14292\,
            I => \N__14279\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__14291\,
            I => \N__14275\
        );

    \I__1908\ : InMux
    port map (
            O => \N__14290\,
            I => \N__14271\
        );

    \I__1907\ : Sp12to4
    port map (
            O => \N__14287\,
            I => \N__14264\
        );

    \I__1906\ : Sp12to4
    port map (
            O => \N__14282\,
            I => \N__14264\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__14279\,
            I => \N__14264\
        );

    \I__1904\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14261\
        );

    \I__1903\ : InMux
    port map (
            O => \N__14275\,
            I => \N__14256\
        );

    \I__1902\ : InMux
    port map (
            O => \N__14274\,
            I => \N__14256\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__14271\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1900\ : Odrv12
    port map (
            O => \N__14264\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__14261\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__14256\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1897\ : InMux
    port map (
            O => \N__14247\,
            I => \N__14242\
        );

    \I__1896\ : InMux
    port map (
            O => \N__14246\,
            I => \N__14237\
        );

    \I__1895\ : InMux
    port map (
            O => \N__14245\,
            I => \N__14237\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__14242\,
            I => \N__14230\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__14237\,
            I => \N__14230\
        );

    \I__1892\ : InMux
    port map (
            O => \N__14236\,
            I => \N__14227\
        );

    \I__1891\ : InMux
    port map (
            O => \N__14235\,
            I => \N__14221\
        );

    \I__1890\ : Sp12to4
    port map (
            O => \N__14230\,
            I => \N__14216\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__14227\,
            I => \N__14216\
        );

    \I__1888\ : InMux
    port map (
            O => \N__14226\,
            I => \N__14213\
        );

    \I__1887\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14208\
        );

    \I__1886\ : InMux
    port map (
            O => \N__14224\,
            I => \N__14208\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__14221\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1884\ : Odrv12
    port map (
            O => \N__14216\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__14213\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__14208\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__14199\,
            I => \this_vga_signals.m23_1_cascade_\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__14196\,
            I => \N__14193\
        );

    \I__1879\ : InMux
    port map (
            O => \N__14193\,
            I => \N__14188\
        );

    \I__1878\ : InMux
    port map (
            O => \N__14192\,
            I => \N__14183\
        );

    \I__1877\ : InMux
    port map (
            O => \N__14191\,
            I => \N__14183\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__14188\,
            I => \N__14175\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__14183\,
            I => \N__14175\
        );

    \I__1874\ : InMux
    port map (
            O => \N__14182\,
            I => \N__14172\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__14181\,
            I => \N__14167\
        );

    \I__1872\ : InMux
    port map (
            O => \N__14180\,
            I => \N__14164\
        );

    \I__1871\ : Sp12to4
    port map (
            O => \N__14175\,
            I => \N__14159\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__14172\,
            I => \N__14159\
        );

    \I__1869\ : InMux
    port map (
            O => \N__14171\,
            I => \N__14156\
        );

    \I__1868\ : InMux
    port map (
            O => \N__14170\,
            I => \N__14151\
        );

    \I__1867\ : InMux
    port map (
            O => \N__14167\,
            I => \N__14151\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__14164\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1865\ : Odrv12
    port map (
            O => \N__14159\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__14156\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__14151\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1862\ : InMux
    port map (
            O => \N__14142\,
            I => \N__14139\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__14139\,
            I => \N__14136\
        );

    \I__1860\ : Span4Mux_v
    port map (
            O => \N__14136\,
            I => \N__14133\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__14133\,
            I => \M_this_data_tmp_qZ0Z_6\
        );

    \I__1858\ : InMux
    port map (
            O => \N__14130\,
            I => \N__14127\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__14127\,
            I => \N__14124\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__14124\,
            I => \this_ppu.un3_sprites_addr_cry_1_c_RNITOBZ0Z8\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__14121\,
            I => \N__14118\
        );

    \I__1854\ : CascadeBuf
    port map (
            O => \N__14118\,
            I => \N__14115\
        );

    \I__1853\ : CascadeMux
    port map (
            O => \N__14115\,
            I => \N__14112\
        );

    \I__1852\ : CascadeBuf
    port map (
            O => \N__14112\,
            I => \N__14109\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__14109\,
            I => \N__14106\
        );

    \I__1850\ : CascadeBuf
    port map (
            O => \N__14106\,
            I => \N__14103\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__14103\,
            I => \N__14100\
        );

    \I__1848\ : CascadeBuf
    port map (
            O => \N__14100\,
            I => \N__14097\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__14097\,
            I => \N__14094\
        );

    \I__1846\ : CascadeBuf
    port map (
            O => \N__14094\,
            I => \N__14091\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__14091\,
            I => \N__14088\
        );

    \I__1844\ : CascadeBuf
    port map (
            O => \N__14088\,
            I => \N__14085\
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__14085\,
            I => \N__14082\
        );

    \I__1842\ : CascadeBuf
    port map (
            O => \N__14082\,
            I => \N__14079\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__14079\,
            I => \N__14076\
        );

    \I__1840\ : CascadeBuf
    port map (
            O => \N__14076\,
            I => \N__14073\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__14073\,
            I => \N__14070\
        );

    \I__1838\ : CascadeBuf
    port map (
            O => \N__14070\,
            I => \N__14067\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__14067\,
            I => \N__14064\
        );

    \I__1836\ : CascadeBuf
    port map (
            O => \N__14064\,
            I => \N__14061\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__14061\,
            I => \N__14058\
        );

    \I__1834\ : CascadeBuf
    port map (
            O => \N__14058\,
            I => \N__14055\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__14055\,
            I => \N__14052\
        );

    \I__1832\ : CascadeBuf
    port map (
            O => \N__14052\,
            I => \N__14049\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__14049\,
            I => \N__14046\
        );

    \I__1830\ : CascadeBuf
    port map (
            O => \N__14046\,
            I => \N__14043\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__14043\,
            I => \N__14040\
        );

    \I__1828\ : CascadeBuf
    port map (
            O => \N__14040\,
            I => \N__14037\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__14037\,
            I => \N__14034\
        );

    \I__1826\ : CascadeBuf
    port map (
            O => \N__14034\,
            I => \N__14031\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__14031\,
            I => \N__14028\
        );

    \I__1824\ : InMux
    port map (
            O => \N__14028\,
            I => \N__14025\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__14025\,
            I => \N__14022\
        );

    \I__1822\ : Span12Mux_s5_v
    port map (
            O => \N__14022\,
            I => \N__14019\
        );

    \I__1821\ : Span12Mux_h
    port map (
            O => \N__14019\,
            I => \N__14016\
        );

    \I__1820\ : Odrv12
    port map (
            O => \N__14016\,
            I => \M_this_ppu_sprites_addr_2\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__14013\,
            I => \this_ppu.un1_M_haddress_q_c1_cascade_\
        );

    \I__1818\ : CEMux
    port map (
            O => \N__14010\,
            I => \N__14007\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__14007\,
            I => \N__14004\
        );

    \I__1816\ : Span4Mux_h
    port map (
            O => \N__14004\,
            I => \N__14001\
        );

    \I__1815\ : Span4Mux_v
    port map (
            O => \N__14001\,
            I => \N__13998\
        );

    \I__1814\ : Span4Mux_v
    port map (
            O => \N__13998\,
            I => \N__13992\
        );

    \I__1813\ : InMux
    port map (
            O => \N__13997\,
            I => \N__13987\
        );

    \I__1812\ : InMux
    port map (
            O => \N__13996\,
            I => \N__13987\
        );

    \I__1811\ : InMux
    port map (
            O => \N__13995\,
            I => \N__13984\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__13992\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__13987\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__13984\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__1807\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13972\
        );

    \I__1806\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13967\
        );

    \I__1805\ : InMux
    port map (
            O => \N__13975\,
            I => \N__13967\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__13972\,
            I => \this_ppu.N_134\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__13967\,
            I => \this_ppu.N_134\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__13962\,
            I => \N__13959\
        );

    \I__1801\ : CascadeBuf
    port map (
            O => \N__13959\,
            I => \N__13956\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__13956\,
            I => \N__13953\
        );

    \I__1799\ : InMux
    port map (
            O => \N__13953\,
            I => \N__13949\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__13952\,
            I => \N__13946\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__13949\,
            I => \N__13942\
        );

    \I__1796\ : InMux
    port map (
            O => \N__13946\,
            I => \N__13939\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__13945\,
            I => \N__13936\
        );

    \I__1794\ : Span4Mux_h
    port map (
            O => \N__13942\,
            I => \N__13933\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__13939\,
            I => \N__13930\
        );

    \I__1792\ : InMux
    port map (
            O => \N__13936\,
            I => \N__13924\
        );

    \I__1791\ : Span4Mux_h
    port map (
            O => \N__13933\,
            I => \N__13921\
        );

    \I__1790\ : Sp12to4
    port map (
            O => \N__13930\,
            I => \N__13918\
        );

    \I__1789\ : InMux
    port map (
            O => \N__13929\,
            I => \N__13915\
        );

    \I__1788\ : InMux
    port map (
            O => \N__13928\,
            I => \N__13912\
        );

    \I__1787\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13909\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__13924\,
            I => \N__13906\
        );

    \I__1785\ : Sp12to4
    port map (
            O => \N__13921\,
            I => \N__13901\
        );

    \I__1784\ : Span12Mux_h
    port map (
            O => \N__13918\,
            I => \N__13901\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__13915\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__13912\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__13909\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__1780\ : Odrv12
    port map (
            O => \N__13906\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__1779\ : Odrv12
    port map (
            O => \N__13901\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__13890\,
            I => \N__13887\
        );

    \I__1777\ : InMux
    port map (
            O => \N__13887\,
            I => \N__13884\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__13884\,
            I => \N__13881\
        );

    \I__1775\ : Span4Mux_v
    port map (
            O => \N__13881\,
            I => \N__13877\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__13880\,
            I => \N__13874\
        );

    \I__1773\ : Span4Mux_v
    port map (
            O => \N__13877\,
            I => \N__13870\
        );

    \I__1772\ : InMux
    port map (
            O => \N__13874\,
            I => \N__13867\
        );

    \I__1771\ : InMux
    port map (
            O => \N__13873\,
            I => \N__13860\
        );

    \I__1770\ : Span4Mux_v
    port map (
            O => \N__13870\,
            I => \N__13855\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__13867\,
            I => \N__13855\
        );

    \I__1768\ : InMux
    port map (
            O => \N__13866\,
            I => \N__13850\
        );

    \I__1767\ : InMux
    port map (
            O => \N__13865\,
            I => \N__13850\
        );

    \I__1766\ : InMux
    port map (
            O => \N__13864\,
            I => \N__13845\
        );

    \I__1765\ : InMux
    port map (
            O => \N__13863\,
            I => \N__13845\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__13860\,
            I => \N__13840\
        );

    \I__1763\ : Span4Mux_h
    port map (
            O => \N__13855\,
            I => \N__13840\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__13850\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__13845\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__13840\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__1759\ : InMux
    port map (
            O => \N__13833\,
            I => \N__13830\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__13830\,
            I => \this_ppu.un1_M_haddress_q_c2\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__13827\,
            I => \N__13824\
        );

    \I__1756\ : CascadeBuf
    port map (
            O => \N__13824\,
            I => \N__13821\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__13821\,
            I => \N__13817\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__13820\,
            I => \N__13814\
        );

    \I__1753\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13810\
        );

    \I__1752\ : InMux
    port map (
            O => \N__13814\,
            I => \N__13807\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__13813\,
            I => \N__13804\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__13810\,
            I => \N__13801\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__13807\,
            I => \N__13798\
        );

    \I__1748\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13793\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__13801\,
            I => \N__13788\
        );

    \I__1746\ : Span4Mux_v
    port map (
            O => \N__13798\,
            I => \N__13788\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__13797\,
            I => \N__13785\
        );

    \I__1744\ : InMux
    port map (
            O => \N__13796\,
            I => \N__13782\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__13793\,
            I => \N__13779\
        );

    \I__1742\ : Span4Mux_h
    port map (
            O => \N__13788\,
            I => \N__13776\
        );

    \I__1741\ : InMux
    port map (
            O => \N__13785\,
            I => \N__13773\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__13782\,
            I => \N__13768\
        );

    \I__1739\ : Span4Mux_h
    port map (
            O => \N__13779\,
            I => \N__13768\
        );

    \I__1738\ : Span4Mux_v
    port map (
            O => \N__13776\,
            I => \N__13765\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__13773\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__1736\ : Odrv4
    port map (
            O => \N__13768\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__1735\ : Odrv4
    port map (
            O => \N__13765\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__1734\ : InMux
    port map (
            O => \N__13758\,
            I => \N__13755\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__13755\,
            I => \this_ppu.N_128\
        );

    \I__1732\ : InMux
    port map (
            O => \N__13752\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__1731\ : InMux
    port map (
            O => \N__13749\,
            I => \bfn_12_22_0_\
        );

    \I__1730\ : InMux
    port map (
            O => \N__13746\,
            I => \N__13742\
        );

    \I__1729\ : InMux
    port map (
            O => \N__13745\,
            I => \N__13739\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__13742\,
            I => \this_vga_signals.M_pcounter_q_i_3_0\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__13739\,
            I => \this_vga_signals.M_pcounter_q_i_3_0\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__13734\,
            I => \N__13729\
        );

    \I__1725\ : InMux
    port map (
            O => \N__13733\,
            I => \N__13725\
        );

    \I__1724\ : InMux
    port map (
            O => \N__13732\,
            I => \N__13722\
        );

    \I__1723\ : InMux
    port map (
            O => \N__13729\,
            I => \N__13717\
        );

    \I__1722\ : InMux
    port map (
            O => \N__13728\,
            I => \N__13717\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__13725\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__13722\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__13717\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__13710\,
            I => \N__13705\
        );

    \I__1717\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13702\
        );

    \I__1716\ : InMux
    port map (
            O => \N__13708\,
            I => \N__13697\
        );

    \I__1715\ : InMux
    port map (
            O => \N__13705\,
            I => \N__13697\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__13702\,
            I => \N__13692\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__13697\,
            I => \N__13692\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__13692\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__1711\ : InMux
    port map (
            O => \N__13689\,
            I => \N__13686\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__13686\,
            I => \N__13683\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__13683\,
            I => \N__13680\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__13680\,
            I => \N_815_0\
        );

    \I__1707\ : InMux
    port map (
            O => \N__13677\,
            I => \N__13674\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__13674\,
            I => \N__13671\
        );

    \I__1705\ : Span4Mux_h
    port map (
            O => \N__13671\,
            I => \N__13668\
        );

    \I__1704\ : Span4Mux_h
    port map (
            O => \N__13668\,
            I => \N__13665\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__13665\,
            I => \N_814_0\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__13662\,
            I => \N__13659\
        );

    \I__1701\ : CascadeBuf
    port map (
            O => \N__13659\,
            I => \N__13656\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__13656\,
            I => \N__13653\
        );

    \I__1699\ : InMux
    port map (
            O => \N__13653\,
            I => \N__13650\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__13650\,
            I => \N__13647\
        );

    \I__1697\ : Odrv12
    port map (
            O => \N__13647\,
            I => \this_ppu_M_vaddress_q_i_6\
        );

    \I__1696\ : InMux
    port map (
            O => \N__13644\,
            I => \N__13641\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__13641\,
            I => \N__13638\
        );

    \I__1694\ : Odrv12
    port map (
            O => \N__13638\,
            I => \M_this_data_tmp_qZ0Z_1\
        );

    \I__1693\ : InMux
    port map (
            O => \N__13635\,
            I => \N__13632\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__13632\,
            I => \N__13629\
        );

    \I__1691\ : Span4Mux_h
    port map (
            O => \N__13629\,
            I => \N__13626\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__13626\,
            I => \M_this_data_tmp_qZ0Z_24\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__13623\,
            I => \N__13620\
        );

    \I__1688\ : InMux
    port map (
            O => \N__13620\,
            I => \N__13617\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__13617\,
            I => \N__13614\
        );

    \I__1686\ : Span4Mux_h
    port map (
            O => \N__13614\,
            I => \N__13611\
        );

    \I__1685\ : Span4Mux_v
    port map (
            O => \N__13611\,
            I => \N__13608\
        );

    \I__1684\ : Span4Mux_v
    port map (
            O => \N__13608\,
            I => \N__13601\
        );

    \I__1683\ : InMux
    port map (
            O => \N__13607\,
            I => \N__13596\
        );

    \I__1682\ : InMux
    port map (
            O => \N__13606\,
            I => \N__13596\
        );

    \I__1681\ : InMux
    port map (
            O => \N__13605\,
            I => \N__13591\
        );

    \I__1680\ : InMux
    port map (
            O => \N__13604\,
            I => \N__13591\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__13601\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__13596\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__13591\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__13584\,
            I => \N__13581\
        );

    \I__1675\ : CascadeBuf
    port map (
            O => \N__13581\,
            I => \N__13578\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__13578\,
            I => \N__13573\
        );

    \I__1673\ : CascadeMux
    port map (
            O => \N__13577\,
            I => \N__13570\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__13576\,
            I => \N__13567\
        );

    \I__1671\ : InMux
    port map (
            O => \N__13573\,
            I => \N__13564\
        );

    \I__1670\ : InMux
    port map (
            O => \N__13570\,
            I => \N__13561\
        );

    \I__1669\ : InMux
    port map (
            O => \N__13567\,
            I => \N__13555\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__13564\,
            I => \N__13550\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__13561\,
            I => \N__13550\
        );

    \I__1666\ : InMux
    port map (
            O => \N__13560\,
            I => \N__13545\
        );

    \I__1665\ : InMux
    port map (
            O => \N__13559\,
            I => \N__13545\
        );

    \I__1664\ : InMux
    port map (
            O => \N__13558\,
            I => \N__13542\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__13555\,
            I => \N__13537\
        );

    \I__1662\ : Span12Mux_v
    port map (
            O => \N__13550\,
            I => \N__13537\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__13545\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__13542\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__1659\ : Odrv12
    port map (
            O => \N__13537\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__13530\,
            I => \this_ppu.un1_M_haddress_q_c5_cascade_\
        );

    \I__1657\ : InMux
    port map (
            O => \N__13527\,
            I => \N__13523\
        );

    \I__1656\ : InMux
    port map (
            O => \N__13526\,
            I => \N__13520\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__13523\,
            I => \this_ppu.M_haddress_qZ0Z_7\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__13520\,
            I => \this_ppu.M_haddress_qZ0Z_7\
        );

    \I__1653\ : InMux
    port map (
            O => \N__13515\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__1652\ : InMux
    port map (
            O => \N__13512\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__1651\ : InMux
    port map (
            O => \N__13509\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__1650\ : InMux
    port map (
            O => \N__13506\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__1649\ : InMux
    port map (
            O => \N__13503\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__1648\ : InMux
    port map (
            O => \N__13500\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__1647\ : InMux
    port map (
            O => \N__13497\,
            I => \N__13494\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__13494\,
            I => \N__13491\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__13491\,
            I => \M_this_data_tmp_qZ0Z_13\
        );

    \I__1644\ : InMux
    port map (
            O => \N__13488\,
            I => \N__13485\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__13485\,
            I => \N__13482\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__13482\,
            I => \M_this_data_tmp_qZ0Z_9\
        );

    \I__1641\ : InMux
    port map (
            O => \N__13479\,
            I => \N__13476\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__13476\,
            I => \N__13473\
        );

    \I__1639\ : Span4Mux_h
    port map (
            O => \N__13473\,
            I => \N__13470\
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__13470\,
            I => \M_this_data_tmp_qZ0Z_0\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__13467\,
            I => \M_this_ppu_vram_data_0_cascade_\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__13464\,
            I => \this_ppu.N_134_cascade_\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__13461\,
            I => \this_ppu.un1_M_haddress_q_c2_cascade_\
        );

    \I__1634\ : InMux
    port map (
            O => \N__13458\,
            I => \N__13452\
        );

    \I__1633\ : InMux
    port map (
            O => \N__13457\,
            I => \N__13452\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__13452\,
            I => \this_ppu.un1_M_haddress_q_c5\
        );

    \I__1631\ : InMux
    port map (
            O => \N__13449\,
            I => \N__13446\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__13446\,
            I => \this_vga_signals.i5_mux\
        );

    \I__1629\ : IoInMux
    port map (
            O => \N__13443\,
            I => \N__13440\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__13440\,
            I => \N__13437\
        );

    \I__1627\ : Span12Mux_s7_v
    port map (
            O => \N__13437\,
            I => \N__13434\
        );

    \I__1626\ : Odrv12
    port map (
            O => \N__13434\,
            I => this_vga_signals_hsync_1_i
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__13431\,
            I => \N__13428\
        );

    \I__1624\ : CascadeBuf
    port map (
            O => \N__13428\,
            I => \N__13425\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__13425\,
            I => \N__13422\
        );

    \I__1622\ : InMux
    port map (
            O => \N__13422\,
            I => \N__13419\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__13419\,
            I => \N__13416\
        );

    \I__1620\ : Span4Mux_h
    port map (
            O => \N__13416\,
            I => \N__13413\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__13413\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__1618\ : InMux
    port map (
            O => \N__13410\,
            I => \N__13407\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__13407\,
            I => \N__13404\
        );

    \I__1616\ : Span4Mux_v
    port map (
            O => \N__13404\,
            I => \N__13401\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__13401\,
            I => \N_63_0\
        );

    \I__1614\ : InMux
    port map (
            O => \N__13398\,
            I => \N__13395\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__13395\,
            I => \N__13391\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__13394\,
            I => \N__13387\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__13391\,
            I => \N__13383\
        );

    \I__1610\ : InMux
    port map (
            O => \N__13390\,
            I => \N__13380\
        );

    \I__1609\ : InMux
    port map (
            O => \N__13387\,
            I => \N__13375\
        );

    \I__1608\ : InMux
    port map (
            O => \N__13386\,
            I => \N__13375\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__13383\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__13380\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__13375\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1604\ : InMux
    port map (
            O => \N__13368\,
            I => \N__13365\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__13365\,
            I => \N__13359\
        );

    \I__1602\ : InMux
    port map (
            O => \N__13364\,
            I => \N__13356\
        );

    \I__1601\ : InMux
    port map (
            O => \N__13363\,
            I => \N__13351\
        );

    \I__1600\ : InMux
    port map (
            O => \N__13362\,
            I => \N__13351\
        );

    \I__1599\ : Odrv12
    port map (
            O => \N__13359\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__13356\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__13351\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__13344\,
            I => \N__13341\
        );

    \I__1595\ : InMux
    port map (
            O => \N__13341\,
            I => \N__13338\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__13338\,
            I => \N__13335\
        );

    \I__1593\ : Span4Mux_h
    port map (
            O => \N__13335\,
            I => \N__13332\
        );

    \I__1592\ : Odrv4
    port map (
            O => \N__13332\,
            I => \M_this_vga_signals_address_3\
        );

    \I__1591\ : InMux
    port map (
            O => \N__13329\,
            I => \N__13326\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__13326\,
            I => \this_vga_signals.SUM_3_1\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__13323\,
            I => \N__13320\
        );

    \I__1588\ : InMux
    port map (
            O => \N__13320\,
            I => \N__13317\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__13317\,
            I => \N__13314\
        );

    \I__1586\ : Span4Mux_h
    port map (
            O => \N__13314\,
            I => \N__13311\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__13311\,
            I => \M_this_vga_signals_address_6\
        );

    \I__1584\ : InMux
    port map (
            O => \N__13308\,
            I => \N__13305\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__13305\,
            I => \N__13302\
        );

    \I__1582\ : Span4Mux_h
    port map (
            O => \N__13302\,
            I => \N__13299\
        );

    \I__1581\ : Odrv4
    port map (
            O => \N__13299\,
            I => \M_this_data_tmp_qZ0Z_29\
        );

    \I__1580\ : InMux
    port map (
            O => \N__13296\,
            I => \N__13293\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__13293\,
            I => \N__13290\
        );

    \I__1578\ : Odrv12
    port map (
            O => \N__13290\,
            I => \M_this_data_tmp_qZ0Z_5\
        );

    \I__1577\ : InMux
    port map (
            O => \N__13287\,
            I => \N__13284\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__13284\,
            I => \N__13281\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__13281\,
            I => \M_this_data_tmp_qZ0Z_12\
        );

    \I__1574\ : InMux
    port map (
            O => \N__13278\,
            I => \N__13272\
        );

    \I__1573\ : InMux
    port map (
            O => \N__13277\,
            I => \N__13265\
        );

    \I__1572\ : InMux
    port map (
            O => \N__13276\,
            I => \N__13265\
        );

    \I__1571\ : InMux
    port map (
            O => \N__13275\,
            I => \N__13265\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__13272\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__13265\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1568\ : InMux
    port map (
            O => \N__13260\,
            I => \N__13256\
        );

    \I__1567\ : InMux
    port map (
            O => \N__13259\,
            I => \N__13253\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__13256\,
            I => \N_3_0\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__13253\,
            I => \N_3_0\
        );

    \I__1564\ : InMux
    port map (
            O => \N__13248\,
            I => \N__13245\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__13245\,
            I => \this_vga_signals.M_pcounter_q_3_0\
        );

    \I__1562\ : InMux
    port map (
            O => \N__13242\,
            I => \N__13236\
        );

    \I__1561\ : InMux
    port map (
            O => \N__13241\,
            I => \N__13236\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__13236\,
            I => \this_vga_signals.N_17_0\
        );

    \I__1559\ : InMux
    port map (
            O => \N__13233\,
            I => \N__13230\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__13230\,
            I => \this_vga_signals.M_hcounter_q_RNI9JJM1Z0Z_0\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__13227\,
            I => \this_vga_signals.M_hcounter_q_RNIADGD1Z0Z_5_cascade_\
        );

    \I__1556\ : IoInMux
    port map (
            O => \N__13224\,
            I => \N__13221\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__13221\,
            I => \N__13218\
        );

    \I__1554\ : Span4Mux_s1_v
    port map (
            O => \N__13218\,
            I => \N__13215\
        );

    \I__1553\ : Sp12to4
    port map (
            O => \N__13215\,
            I => \N__13212\
        );

    \I__1552\ : Span12Mux_s10_h
    port map (
            O => \N__13212\,
            I => \N__13209\
        );

    \I__1551\ : Odrv12
    port map (
            O => \N__13209\,
            I => this_vga_signals_hvisibility_i
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__13206\,
            I => \this_vga_signals.mult1_un89_sum_axbxc3_2_cascade_\
        );

    \I__1549\ : InMux
    port map (
            O => \N__13203\,
            I => \N__13200\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__13200\,
            I => \this_vga_signals.mult1_un89_sum_c3_0\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__13197\,
            I => \N__13194\
        );

    \I__1546\ : InMux
    port map (
            O => \N__13194\,
            I => \N__13191\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__13191\,
            I => \N__13188\
        );

    \I__1544\ : Span4Mux_v
    port map (
            O => \N__13188\,
            I => \N__13185\
        );

    \I__1543\ : Span4Mux_v
    port map (
            O => \N__13185\,
            I => \N__13182\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__13182\,
            I => \M_this_vga_signals_address_0\
        );

    \I__1541\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13176\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__13176\,
            I => \N__13173\
        );

    \I__1539\ : Span4Mux_v
    port map (
            O => \N__13173\,
            I => \N__13169\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__13172\,
            I => \N__13166\
        );

    \I__1537\ : Span4Mux_v
    port map (
            O => \N__13169\,
            I => \N__13162\
        );

    \I__1536\ : InMux
    port map (
            O => \N__13166\,
            I => \N__13157\
        );

    \I__1535\ : InMux
    port map (
            O => \N__13165\,
            I => \N__13157\
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__13162\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__13157\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1532\ : InMux
    port map (
            O => \N__13152\,
            I => \N__13149\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__13149\,
            I => \this_vga_signals.mult1_un82_sum_axb1\
        );

    \I__1530\ : InMux
    port map (
            O => \N__13146\,
            I => \N__13143\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__13143\,
            I => \N__13139\
        );

    \I__1528\ : InMux
    port map (
            O => \N__13142\,
            I => \N__13136\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__13139\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_1\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__13136\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_1\
        );

    \I__1525\ : InMux
    port map (
            O => \N__13131\,
            I => \N__13128\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__13128\,
            I => \N__13125\
        );

    \I__1523\ : Span4Mux_v
    port map (
            O => \N__13125\,
            I => \N__13121\
        );

    \I__1522\ : InMux
    port map (
            O => \N__13124\,
            I => \N__13118\
        );

    \I__1521\ : Odrv4
    port map (
            O => \N__13121\,
            I => \this_vga_signals.mult1_un82_sum_c3\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__13118\,
            I => \this_vga_signals.mult1_un82_sum_c3\
        );

    \I__1519\ : InMux
    port map (
            O => \N__13113\,
            I => \N__13107\
        );

    \I__1518\ : InMux
    port map (
            O => \N__13112\,
            I => \N__13107\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__13107\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3\
        );

    \I__1516\ : InMux
    port map (
            O => \N__13104\,
            I => \N__13101\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__13101\,
            I => \N__13098\
        );

    \I__1514\ : Span4Mux_h
    port map (
            O => \N__13098\,
            I => \N__13095\
        );

    \I__1513\ : Span4Mux_v
    port map (
            O => \N__13095\,
            I => \N__13091\
        );

    \I__1512\ : InMux
    port map (
            O => \N__13094\,
            I => \N__13088\
        );

    \I__1511\ : Odrv4
    port map (
            O => \N__13091\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__13088\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__1509\ : InMux
    port map (
            O => \N__13083\,
            I => \N__13077\
        );

    \I__1508\ : InMux
    port map (
            O => \N__13082\,
            I => \N__13077\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__13077\,
            I => \this_vga_signals.mult1_un61_sum_axb1\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__13074\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9_cascade_\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__13071\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_1_cascade_\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__13068\,
            I => \N__13065\
        );

    \I__1503\ : InMux
    port map (
            O => \N__13065\,
            I => \N__13056\
        );

    \I__1502\ : InMux
    port map (
            O => \N__13064\,
            I => \N__13056\
        );

    \I__1501\ : InMux
    port map (
            O => \N__13063\,
            I => \N__13056\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__13056\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9\
        );

    \I__1499\ : InMux
    port map (
            O => \N__13053\,
            I => \N__13050\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__13050\,
            I => \N__13046\
        );

    \I__1497\ : InMux
    port map (
            O => \N__13049\,
            I => \N__13043\
        );

    \I__1496\ : Span12Mux_s10_v
    port map (
            O => \N__13046\,
            I => \N__13035\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__13043\,
            I => \N__13032\
        );

    \I__1494\ : InMux
    port map (
            O => \N__13042\,
            I => \N__13023\
        );

    \I__1493\ : InMux
    port map (
            O => \N__13041\,
            I => \N__13023\
        );

    \I__1492\ : InMux
    port map (
            O => \N__13040\,
            I => \N__13023\
        );

    \I__1491\ : InMux
    port map (
            O => \N__13039\,
            I => \N__13023\
        );

    \I__1490\ : InMux
    port map (
            O => \N__13038\,
            I => \N__13020\
        );

    \I__1489\ : Odrv12
    port map (
            O => \N__13035\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__13032\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__13023\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__13020\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__13011\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_cascade_\
        );

    \I__1484\ : InMux
    port map (
            O => \N__13008\,
            I => \N__13005\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__13005\,
            I => \this_vga_signals.mult1_un68_sum_axb1\
        );

    \I__1482\ : CascadeMux
    port map (
            O => \N__13002\,
            I => \this_vga_signals.if_i4_mux_0_cascade_\
        );

    \I__1481\ : InMux
    port map (
            O => \N__12999\,
            I => \N__12994\
        );

    \I__1480\ : InMux
    port map (
            O => \N__12998\,
            I => \N__12991\
        );

    \I__1479\ : InMux
    port map (
            O => \N__12997\,
            I => \N__12988\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__12994\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__12991\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__12988\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0\
        );

    \I__1475\ : InMux
    port map (
            O => \N__12981\,
            I => \N__12978\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__12978\,
            I => \this_vga_signals.M_hcounter_q_RNIUULS4Z0Z_3\
        );

    \I__1473\ : InMux
    port map (
            O => \N__12975\,
            I => \N__12971\
        );

    \I__1472\ : InMux
    port map (
            O => \N__12974\,
            I => \N__12968\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__12971\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__12968\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__12963\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__12960\,
            I => \N__12957\
        );

    \I__1467\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12954\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__12954\,
            I => \this_vga_signals.if_m2_2\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__12951\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3_1_cascade_\
        );

    \I__1464\ : InMux
    port map (
            O => \N__12948\,
            I => \N__12944\
        );

    \I__1463\ : InMux
    port map (
            O => \N__12947\,
            I => \N__12941\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__12944\,
            I => \this_vga_signals.d_N_3_0_i\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__12941\,
            I => \this_vga_signals.d_N_3_0_i\
        );

    \I__1460\ : InMux
    port map (
            O => \N__12936\,
            I => \N__12933\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__12933\,
            I => \this_vga_signals.mult1_un82_sum_c2_0\
        );

    \I__1458\ : InMux
    port map (
            O => \N__12930\,
            I => \N__12927\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__12927\,
            I => \N__12924\
        );

    \I__1456\ : Odrv4
    port map (
            O => \N__12924\,
            I => \M_this_data_tmp_qZ0Z_28\
        );

    \I__1455\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12918\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__12918\,
            I => \N__12915\
        );

    \I__1453\ : Span4Mux_h
    port map (
            O => \N__12915\,
            I => \N__12912\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__12912\,
            I => \N_833_0\
        );

    \I__1451\ : InMux
    port map (
            O => \N__12909\,
            I => \N__12906\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__12906\,
            I => \N__12903\
        );

    \I__1449\ : Span4Mux_h
    port map (
            O => \N__12903\,
            I => \N__12899\
        );

    \I__1448\ : InMux
    port map (
            O => \N__12902\,
            I => \N__12896\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__12899\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__12896\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__1445\ : CascadeMux
    port map (
            O => \N__12891\,
            I => \N__12888\
        );

    \I__1444\ : CascadeBuf
    port map (
            O => \N__12888\,
            I => \N__12885\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__12885\,
            I => \N__12882\
        );

    \I__1442\ : InMux
    port map (
            O => \N__12882\,
            I => \N__12879\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__12879\,
            I => \N__12875\
        );

    \I__1440\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12872\
        );

    \I__1439\ : Span4Mux_v
    port map (
            O => \N__12875\,
            I => \N__12869\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__12872\,
            I => \N__12864\
        );

    \I__1437\ : Span4Mux_v
    port map (
            O => \N__12869\,
            I => \N__12864\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__12864\,
            I => \M_this_ppu_vram_addr_i_6\
        );

    \I__1435\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12858\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__12858\,
            I => \M_this_data_tmp_qZ0Z_18\
        );

    \I__1433\ : InMux
    port map (
            O => \N__12855\,
            I => \N__12852\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__12852\,
            I => \N__12849\
        );

    \I__1431\ : Span4Mux_v
    port map (
            O => \N__12849\,
            I => \N__12846\
        );

    \I__1430\ : Span4Mux_h
    port map (
            O => \N__12846\,
            I => \N__12843\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__12843\,
            I => \M_this_oam_ram_write_data_18\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__12840\,
            I => \N__12837\
        );

    \I__1427\ : CascadeBuf
    port map (
            O => \N__12837\,
            I => \N__12834\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__12834\,
            I => \N__12831\
        );

    \I__1425\ : InMux
    port map (
            O => \N__12831\,
            I => \N__12828\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__12828\,
            I => \N__12824\
        );

    \I__1423\ : InMux
    port map (
            O => \N__12827\,
            I => \N__12821\
        );

    \I__1422\ : Span4Mux_v
    port map (
            O => \N__12824\,
            I => \N__12818\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__12821\,
            I => \N__12813\
        );

    \I__1420\ : Span4Mux_v
    port map (
            O => \N__12818\,
            I => \N__12813\
        );

    \I__1419\ : Odrv4
    port map (
            O => \N__12813\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__1418\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12807\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__12807\,
            I => \N__12804\
        );

    \I__1416\ : Odrv4
    port map (
            O => \N__12804\,
            I => \M_this_data_tmp_qZ0Z_30\
        );

    \I__1415\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12798\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__12798\,
            I => \N__12795\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__12795\,
            I => \N_830_0\
        );

    \I__1412\ : InMux
    port map (
            O => \N__12792\,
            I => \N__12789\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__12789\,
            I => \M_this_data_tmp_qZ0Z_16\
        );

    \I__1410\ : InMux
    port map (
            O => \N__12786\,
            I => \N__12783\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__12783\,
            I => \N__12780\
        );

    \I__1408\ : Span4Mux_h
    port map (
            O => \N__12780\,
            I => \N__12777\
        );

    \I__1407\ : Odrv4
    port map (
            O => \N__12777\,
            I => \M_this_oam_ram_write_data_16\
        );

    \I__1406\ : InMux
    port map (
            O => \N__12774\,
            I => \N__12771\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__12771\,
            I => \N__12768\
        );

    \I__1404\ : Odrv4
    port map (
            O => \N__12768\,
            I => \M_this_data_tmp_qZ0Z_14\
        );

    \I__1403\ : InMux
    port map (
            O => \N__12765\,
            I => \N__12762\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__12762\,
            I => \N__12759\
        );

    \I__1401\ : Span4Mux_h
    port map (
            O => \N__12759\,
            I => \N__12756\
        );

    \I__1400\ : Odrv4
    port map (
            O => \N__12756\,
            I => \M_this_data_tmp_qZ0Z_27\
        );

    \I__1399\ : InMux
    port map (
            O => \N__12753\,
            I => \N__12750\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__12750\,
            I => \M_this_data_tmp_qZ0Z_3\
        );

    \I__1397\ : InMux
    port map (
            O => \N__12747\,
            I => \N__12744\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__12744\,
            I => \N__12741\
        );

    \I__1395\ : Odrv12
    port map (
            O => \N__12741\,
            I => \M_this_data_tmp_qZ0Z_7\
        );

    \I__1394\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12735\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__12735\,
            I => \M_this_data_tmp_qZ0Z_2\
        );

    \I__1392\ : InMux
    port map (
            O => \N__12732\,
            I => \N__12729\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__12729\,
            I => \N__12726\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__12726\,
            I => \M_this_data_tmp_qZ0Z_4\
        );

    \I__1389\ : InMux
    port map (
            O => \N__12723\,
            I => \N__12720\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__12720\,
            I => \M_this_data_tmp_qZ0Z_25\
        );

    \I__1387\ : InMux
    port map (
            O => \N__12717\,
            I => \N__12714\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__12714\,
            I => \N__12711\
        );

    \I__1385\ : Odrv4
    port map (
            O => \N__12711\,
            I => \M_this_data_tmp_qZ0Z_31\
        );

    \I__1384\ : InMux
    port map (
            O => \N__12708\,
            I => \N__12705\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__12705\,
            I => \M_this_vga_signals_pixel_clk_0_0\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__12702\,
            I => \this_vga_ramdac.i2_mux_0_cascade_\
        );

    \I__1381\ : InMux
    port map (
            O => \N__12699\,
            I => \N__12696\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__12696\,
            I => \N__12692\
        );

    \I__1379\ : InMux
    port map (
            O => \N__12695\,
            I => \N__12689\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__12692\,
            I => \this_vga_ramdac.N_2615_reto\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__12689\,
            I => \this_vga_ramdac.N_2615_reto\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__12684\,
            I => \this_vga_ramdac.m16_cascade_\
        );

    \I__1375\ : InMux
    port map (
            O => \N__12681\,
            I => \N__12676\
        );

    \I__1374\ : InMux
    port map (
            O => \N__12680\,
            I => \N__12671\
        );

    \I__1373\ : InMux
    port map (
            O => \N__12679\,
            I => \N__12671\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__12676\,
            I => \N__12663\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__12671\,
            I => \N__12663\
        );

    \I__1370\ : InMux
    port map (
            O => \N__12670\,
            I => \N__12660\
        );

    \I__1369\ : InMux
    port map (
            O => \N__12669\,
            I => \N__12655\
        );

    \I__1368\ : InMux
    port map (
            O => \N__12668\,
            I => \N__12655\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__12663\,
            I => \G_480\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__12660\,
            I => \G_480\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__12655\,
            I => \G_480\
        );

    \I__1364\ : InMux
    port map (
            O => \N__12648\,
            I => \N__12645\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__12645\,
            I => \N__12641\
        );

    \I__1362\ : InMux
    port map (
            O => \N__12644\,
            I => \N__12638\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__12641\,
            I => \this_vga_ramdac.N_2613_reto\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__12638\,
            I => \this_vga_ramdac.N_2613_reto\
        );

    \I__1359\ : InMux
    port map (
            O => \N__12633\,
            I => \N__12630\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__12630\,
            I => \N__12627\
        );

    \I__1357\ : Span4Mux_h
    port map (
            O => \N__12627\,
            I => \N__12624\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__12624\,
            I => \N_73_0\
        );

    \I__1355\ : InMux
    port map (
            O => \N__12621\,
            I => \N__12618\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__12618\,
            I => \N__12615\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__12615\,
            I => \this_vga_ramdac.N_24_mux\
        );

    \I__1352\ : InMux
    port map (
            O => \N__12612\,
            I => \N__12609\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__12609\,
            I => \N__12606\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__12606\,
            I => \this_vga_ramdac.m19\
        );

    \I__1349\ : InMux
    port map (
            O => \N__12603\,
            I => \N__12594\
        );

    \I__1348\ : InMux
    port map (
            O => \N__12602\,
            I => \N__12594\
        );

    \I__1347\ : InMux
    port map (
            O => \N__12601\,
            I => \N__12594\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__12594\,
            I => \N__12589\
        );

    \I__1345\ : InMux
    port map (
            O => \N__12593\,
            I => \N__12584\
        );

    \I__1344\ : InMux
    port map (
            O => \N__12592\,
            I => \N__12584\
        );

    \I__1343\ : Span4Mux_v
    port map (
            O => \N__12589\,
            I => \N__12578\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__12584\,
            I => \N__12578\
        );

    \I__1341\ : InMux
    port map (
            O => \N__12583\,
            I => \N__12575\
        );

    \I__1340\ : Span4Mux_h
    port map (
            O => \N__12578\,
            I => \N__12572\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__12575\,
            I => \N__12569\
        );

    \I__1338\ : Span4Mux_v
    port map (
            O => \N__12572\,
            I => \N__12566\
        );

    \I__1337\ : Span4Mux_v
    port map (
            O => \N__12569\,
            I => \N__12563\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__12566\,
            I => \M_this_vram_read_data_0\
        );

    \I__1335\ : Odrv4
    port map (
            O => \N__12563\,
            I => \M_this_vram_read_data_0\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__12558\,
            I => \N__12553\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__12557\,
            I => \N__12547\
        );

    \I__1332\ : CascadeMux
    port map (
            O => \N__12556\,
            I => \N__12544\
        );

    \I__1331\ : InMux
    port map (
            O => \N__12553\,
            I => \N__12537\
        );

    \I__1330\ : InMux
    port map (
            O => \N__12552\,
            I => \N__12537\
        );

    \I__1329\ : InMux
    port map (
            O => \N__12551\,
            I => \N__12537\
        );

    \I__1328\ : InMux
    port map (
            O => \N__12550\,
            I => \N__12532\
        );

    \I__1327\ : InMux
    port map (
            O => \N__12547\,
            I => \N__12532\
        );

    \I__1326\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12529\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__12537\,
            I => \N__12526\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__12532\,
            I => \N__12521\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__12529\,
            I => \N__12521\
        );

    \I__1322\ : Span4Mux_h
    port map (
            O => \N__12526\,
            I => \N__12518\
        );

    \I__1321\ : Span4Mux_h
    port map (
            O => \N__12521\,
            I => \N__12515\
        );

    \I__1320\ : Span4Mux_v
    port map (
            O => \N__12518\,
            I => \N__12512\
        );

    \I__1319\ : Odrv4
    port map (
            O => \N__12515\,
            I => \M_this_vram_read_data_3\
        );

    \I__1318\ : Odrv4
    port map (
            O => \N__12512\,
            I => \M_this_vram_read_data_3\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__12507\,
            I => \N__12502\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__12506\,
            I => \N__12498\
        );

    \I__1315\ : InMux
    port map (
            O => \N__12505\,
            I => \N__12489\
        );

    \I__1314\ : InMux
    port map (
            O => \N__12502\,
            I => \N__12489\
        );

    \I__1313\ : InMux
    port map (
            O => \N__12501\,
            I => \N__12489\
        );

    \I__1312\ : InMux
    port map (
            O => \N__12498\,
            I => \N__12484\
        );

    \I__1311\ : InMux
    port map (
            O => \N__12497\,
            I => \N__12484\
        );

    \I__1310\ : InMux
    port map (
            O => \N__12496\,
            I => \N__12481\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__12489\,
            I => \N__12476\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__12484\,
            I => \N__12476\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__12481\,
            I => \N__12473\
        );

    \I__1306\ : Span12Mux_v
    port map (
            O => \N__12476\,
            I => \N__12470\
        );

    \I__1305\ : Span4Mux_v
    port map (
            O => \N__12473\,
            I => \N__12467\
        );

    \I__1304\ : Odrv12
    port map (
            O => \N__12470\,
            I => \M_this_vram_read_data_1\
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__12467\,
            I => \M_this_vram_read_data_1\
        );

    \I__1302\ : InMux
    port map (
            O => \N__12462\,
            I => \N__12456\
        );

    \I__1301\ : InMux
    port map (
            O => \N__12461\,
            I => \N__12456\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__12456\,
            I => \N__12450\
        );

    \I__1299\ : InMux
    port map (
            O => \N__12455\,
            I => \N__12445\
        );

    \I__1298\ : InMux
    port map (
            O => \N__12454\,
            I => \N__12445\
        );

    \I__1297\ : InMux
    port map (
            O => \N__12453\,
            I => \N__12442\
        );

    \I__1296\ : Span4Mux_h
    port map (
            O => \N__12450\,
            I => \N__12439\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__12445\,
            I => \N__12434\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__12442\,
            I => \N__12434\
        );

    \I__1293\ : Span4Mux_v
    port map (
            O => \N__12439\,
            I => \N__12431\
        );

    \I__1292\ : Span4Mux_h
    port map (
            O => \N__12434\,
            I => \N__12428\
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__12431\,
            I => \M_this_vram_read_data_2\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__12428\,
            I => \M_this_vram_read_data_2\
        );

    \I__1289\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12420\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__12420\,
            I => \N__12417\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__12417\,
            I => \this_vga_ramdac.m6\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__12414\,
            I => \this_vga_signals.mult1_un68_sum_axb1_cascade_\
        );

    \I__1285\ : InMux
    port map (
            O => \N__12411\,
            I => \N__12408\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__12408\,
            I => \this_vga_signals.if_m2_0\
        );

    \I__1283\ : InMux
    port map (
            O => \N__12405\,
            I => \N__12402\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__12402\,
            I => \N__12399\
        );

    \I__1281\ : Span4Mux_h
    port map (
            O => \N__12399\,
            I => \N__12396\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__12396\,
            I => \N__12393\
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__12393\,
            I => \N_58_0\
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__12390\,
            I => \N_3_0_cascade_\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__12387\,
            I => \G_480_cascade_\
        );

    \I__1276\ : InMux
    port map (
            O => \N__12384\,
            I => \N__12381\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__12381\,
            I => \N__12377\
        );

    \I__1274\ : InMux
    port map (
            O => \N__12380\,
            I => \N__12374\
        );

    \I__1273\ : Span4Mux_v
    port map (
            O => \N__12377\,
            I => \N__12371\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__12374\,
            I => \N__12368\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__12371\,
            I => \this_vga_ramdac.N_2614_reto\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__12368\,
            I => \this_vga_ramdac.N_2614_reto\
        );

    \I__1269\ : InMux
    port map (
            O => \N__12363\,
            I => \N__12359\
        );

    \I__1268\ : InMux
    port map (
            O => \N__12362\,
            I => \N__12356\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__12359\,
            I => \this_vga_ramdac.N_2611_reto\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__12356\,
            I => \this_vga_ramdac.N_2611_reto\
        );

    \I__1265\ : InMux
    port map (
            O => \N__12351\,
            I => \N__12348\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__12348\,
            I => \N__12344\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__12347\,
            I => \N__12341\
        );

    \I__1262\ : Span4Mux_h
    port map (
            O => \N__12344\,
            I => \N__12338\
        );

    \I__1261\ : InMux
    port map (
            O => \N__12341\,
            I => \N__12335\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__12338\,
            I => \this_vga_ramdac.N_2610_reto\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__12335\,
            I => \this_vga_ramdac.N_2610_reto\
        );

    \I__1258\ : InMux
    port map (
            O => \N__12330\,
            I => \N__12327\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__12327\,
            I => \N_2_0\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__12324\,
            I => \N_2_0_cascade_\
        );

    \I__1255\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12318\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__12318\,
            I => \N__12315\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__12315\,
            I => \M_this_data_tmp_qZ0Z_20\
        );

    \I__1252\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12309\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__12309\,
            I => \M_this_data_tmp_qZ0Z_21\
        );

    \I__1250\ : InMux
    port map (
            O => \N__12306\,
            I => \N__12303\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__12303\,
            I => \M_this_data_tmp_qZ0Z_22\
        );

    \I__1248\ : InMux
    port map (
            O => \N__12300\,
            I => \N__12297\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__12297\,
            I => \N__12294\
        );

    \I__1246\ : Span4Mux_h
    port map (
            O => \N__12294\,
            I => \N__12291\
        );

    \I__1245\ : Odrv4
    port map (
            O => \N__12291\,
            I => \M_this_data_tmp_qZ0Z_23\
        );

    \I__1244\ : InMux
    port map (
            O => \N__12288\,
            I => \N__12285\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__12285\,
            I => \N__12282\
        );

    \I__1242\ : Odrv4
    port map (
            O => \N__12282\,
            I => \this_oam_ram.M_this_oam_ram_read_data_22\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__12279\,
            I => \N__12276\
        );

    \I__1240\ : InMux
    port map (
            O => \N__12276\,
            I => \N__12273\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__12273\,
            I => \M_this_oam_ram_read_data_i_22\
        );

    \I__1238\ : InMux
    port map (
            O => \N__12270\,
            I => \N__12267\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__12267\,
            I => \N__12264\
        );

    \I__1236\ : Span4Mux_h
    port map (
            O => \N__12264\,
            I => \N__12261\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__12261\,
            I => \N_890_0\
        );

    \I__1234\ : InMux
    port map (
            O => \N__12258\,
            I => \N__12255\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__12255\,
            I => \N__12252\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__12252\,
            I => \M_this_oam_ram_write_data_12\
        );

    \I__1231\ : InMux
    port map (
            O => \N__12249\,
            I => \N__12246\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__12246\,
            I => \N__12243\
        );

    \I__1229\ : Span4Mux_h
    port map (
            O => \N__12243\,
            I => \N__12240\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__12240\,
            I => \N_831_0\
        );

    \I__1227\ : InMux
    port map (
            O => \N__12237\,
            I => \N__12234\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__12234\,
            I => \N__12231\
        );

    \I__1225\ : Span4Mux_h
    port map (
            O => \N__12231\,
            I => \N__12228\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__12228\,
            I => \M_this_oam_ram_write_data_24\
        );

    \I__1223\ : InMux
    port map (
            O => \N__12225\,
            I => \N__12222\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__12222\,
            I => \N__12219\
        );

    \I__1221\ : Span4Mux_h
    port map (
            O => \N__12219\,
            I => \N__12216\
        );

    \I__1220\ : Odrv4
    port map (
            O => \N__12216\,
            I => \N_832_0\
        );

    \I__1219\ : InMux
    port map (
            O => \N__12213\,
            I => \N__12210\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__12210\,
            I => \N__12207\
        );

    \I__1217\ : Span4Mux_h
    port map (
            O => \N__12207\,
            I => \N__12204\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__12204\,
            I => \N_893_0\
        );

    \I__1215\ : InMux
    port map (
            O => \N__12201\,
            I => \N__12198\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__12198\,
            I => \M_this_data_tmp_qZ0Z_19\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__12195\,
            I => \N__12192\
        );

    \I__1212\ : InMux
    port map (
            O => \N__12192\,
            I => \N__12189\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__12189\,
            I => \M_this_vga_signals_address_4\
        );

    \I__1210\ : InMux
    port map (
            O => \N__12186\,
            I => \N__12183\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__12183\,
            I => \N__12180\
        );

    \I__1208\ : Span4Mux_s3_v
    port map (
            O => \N__12180\,
            I => \N__12177\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__12177\,
            I => \M_this_map_ram_read_data_1\
        );

    \I__1206\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12171\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__12171\,
            I => \N__12168\
        );

    \I__1204\ : Span12Mux_s6_v
    port map (
            O => \N__12168\,
            I => \N__12165\
        );

    \I__1203\ : Odrv12
    port map (
            O => \N__12165\,
            I => \this_ppu.un3_sprites_addr_cry_6_c_RNIP5LZ0Z8\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__12162\,
            I => \N__12159\
        );

    \I__1201\ : CascadeBuf
    port map (
            O => \N__12159\,
            I => \N__12156\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__12156\,
            I => \N__12153\
        );

    \I__1199\ : CascadeBuf
    port map (
            O => \N__12153\,
            I => \N__12150\
        );

    \I__1198\ : CascadeMux
    port map (
            O => \N__12150\,
            I => \N__12147\
        );

    \I__1197\ : CascadeBuf
    port map (
            O => \N__12147\,
            I => \N__12144\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__12144\,
            I => \N__12141\
        );

    \I__1195\ : CascadeBuf
    port map (
            O => \N__12141\,
            I => \N__12138\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__12138\,
            I => \N__12135\
        );

    \I__1193\ : CascadeBuf
    port map (
            O => \N__12135\,
            I => \N__12132\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__12132\,
            I => \N__12129\
        );

    \I__1191\ : CascadeBuf
    port map (
            O => \N__12129\,
            I => \N__12126\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__12126\,
            I => \N__12123\
        );

    \I__1189\ : CascadeBuf
    port map (
            O => \N__12123\,
            I => \N__12120\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__12120\,
            I => \N__12117\
        );

    \I__1187\ : CascadeBuf
    port map (
            O => \N__12117\,
            I => \N__12114\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__12114\,
            I => \N__12111\
        );

    \I__1185\ : CascadeBuf
    port map (
            O => \N__12111\,
            I => \N__12108\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__12108\,
            I => \N__12105\
        );

    \I__1183\ : CascadeBuf
    port map (
            O => \N__12105\,
            I => \N__12102\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__12102\,
            I => \N__12099\
        );

    \I__1181\ : CascadeBuf
    port map (
            O => \N__12099\,
            I => \N__12096\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__12096\,
            I => \N__12093\
        );

    \I__1179\ : CascadeBuf
    port map (
            O => \N__12093\,
            I => \N__12090\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__12090\,
            I => \N__12087\
        );

    \I__1177\ : CascadeBuf
    port map (
            O => \N__12087\,
            I => \N__12084\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__12084\,
            I => \N__12081\
        );

    \I__1175\ : CascadeBuf
    port map (
            O => \N__12081\,
            I => \N__12078\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__12078\,
            I => \N__12075\
        );

    \I__1173\ : CascadeBuf
    port map (
            O => \N__12075\,
            I => \N__12072\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__12072\,
            I => \N__12069\
        );

    \I__1171\ : InMux
    port map (
            O => \N__12069\,
            I => \N__12066\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__12066\,
            I => \N__12063\
        );

    \I__1169\ : Span12Mux_h
    port map (
            O => \N__12063\,
            I => \N__12060\
        );

    \I__1168\ : Odrv12
    port map (
            O => \N__12060\,
            I => \M_this_ppu_sprites_addr_7\
        );

    \I__1167\ : InMux
    port map (
            O => \N__12057\,
            I => \N__12054\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__12054\,
            I => \M_this_data_tmp_qZ0Z_15\
        );

    \I__1165\ : InMux
    port map (
            O => \N__12051\,
            I => \N__12048\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__12048\,
            I => \M_this_data_tmp_qZ0Z_8\
        );

    \I__1163\ : InMux
    port map (
            O => \N__12045\,
            I => \N__12042\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__12042\,
            I => \M_this_data_tmp_qZ0Z_11\
        );

    \I__1161\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12036\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__12036\,
            I => \N__12033\
        );

    \I__1159\ : Odrv4
    port map (
            O => \N__12033\,
            I => \N_835_0\
        );

    \I__1158\ : InMux
    port map (
            O => \N__12030\,
            I => \N__12027\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__12027\,
            I => \N__12024\
        );

    \I__1156\ : Span4Mux_h
    port map (
            O => \N__12024\,
            I => \N__12021\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__12021\,
            I => \N_897_0\
        );

    \I__1154\ : InMux
    port map (
            O => \N__12018\,
            I => \N__12015\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__12015\,
            I => \N__12012\
        );

    \I__1152\ : Span4Mux_h
    port map (
            O => \N__12012\,
            I => \N__12009\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__12009\,
            I => \N_53_0\
        );

    \I__1150\ : InMux
    port map (
            O => \N__12006\,
            I => \N__12003\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__12003\,
            I => \N__12000\
        );

    \I__1148\ : Span4Mux_v
    port map (
            O => \N__12000\,
            I => \N__11997\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__11997\,
            I => \M_this_oam_ram_write_data_2\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__11994\,
            I => \N__11991\
        );

    \I__1145\ : CascadeBuf
    port map (
            O => \N__11991\,
            I => \N__11988\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__11988\,
            I => \N__11985\
        );

    \I__1143\ : InMux
    port map (
            O => \N__11985\,
            I => \N__11982\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__11982\,
            I => \N__11978\
        );

    \I__1141\ : InMux
    port map (
            O => \N__11981\,
            I => \N__11975\
        );

    \I__1140\ : Span4Mux_v
    port map (
            O => \N__11978\,
            I => \N__11972\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__11975\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__11972\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__1137\ : InMux
    port map (
            O => \N__11967\,
            I => \un1_M_this_map_address_q_cry_6\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__11964\,
            I => \N__11961\
        );

    \I__1135\ : CascadeBuf
    port map (
            O => \N__11961\,
            I => \N__11958\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__11958\,
            I => \N__11955\
        );

    \I__1133\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11952\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__11952\,
            I => \N__11948\
        );

    \I__1131\ : InMux
    port map (
            O => \N__11951\,
            I => \N__11945\
        );

    \I__1130\ : Span4Mux_v
    port map (
            O => \N__11948\,
            I => \N__11942\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__11945\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__11942\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__1127\ : InMux
    port map (
            O => \N__11937\,
            I => \bfn_9_25_0_\
        );

    \I__1126\ : InMux
    port map (
            O => \N__11934\,
            I => \un1_M_this_map_address_q_cry_8\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__11931\,
            I => \N__11928\
        );

    \I__1124\ : CascadeBuf
    port map (
            O => \N__11928\,
            I => \N__11925\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__11925\,
            I => \N__11922\
        );

    \I__1122\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11919\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__11919\,
            I => \N__11915\
        );

    \I__1120\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11912\
        );

    \I__1119\ : Span4Mux_v
    port map (
            O => \N__11915\,
            I => \N__11909\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__11912\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__11909\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__1116\ : InMux
    port map (
            O => \N__11904\,
            I => \N__11901\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__11901\,
            I => \N__11898\
        );

    \I__1114\ : Odrv4
    port map (
            O => \N__11898\,
            I => \this_vga_ramdac.i2_mux\
        );

    \I__1113\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11892\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__11892\,
            I => \N__11888\
        );

    \I__1111\ : InMux
    port map (
            O => \N__11891\,
            I => \N__11885\
        );

    \I__1110\ : Span4Mux_v
    port map (
            O => \N__11888\,
            I => \N__11878\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__11885\,
            I => \N__11878\
        );

    \I__1108\ : InMux
    port map (
            O => \N__11884\,
            I => \N__11875\
        );

    \I__1107\ : InMux
    port map (
            O => \N__11883\,
            I => \N__11870\
        );

    \I__1106\ : Span4Mux_h
    port map (
            O => \N__11878\,
            I => \N__11865\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__11875\,
            I => \N__11865\
        );

    \I__1104\ : InMux
    port map (
            O => \N__11874\,
            I => \N__11862\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__11873\,
            I => \N__11858\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__11870\,
            I => \N__11855\
        );

    \I__1101\ : Span4Mux_v
    port map (
            O => \N__11865\,
            I => \N__11850\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__11862\,
            I => \N__11850\
        );

    \I__1099\ : InMux
    port map (
            O => \N__11861\,
            I => \N__11847\
        );

    \I__1098\ : InMux
    port map (
            O => \N__11858\,
            I => \N__11844\
        );

    \I__1097\ : Odrv12
    port map (
            O => \N__11855\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__1096\ : Odrv4
    port map (
            O => \N__11850\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__11847\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__11844\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__1093\ : IoInMux
    port map (
            O => \N__11835\,
            I => \N__11832\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__11832\,
            I => \N__11829\
        );

    \I__1091\ : Odrv12
    port map (
            O => \N__11829\,
            I => rgb_c_5
        );

    \I__1090\ : InMux
    port map (
            O => \N__11826\,
            I => \N__11823\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__11823\,
            I => \N_60_0\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__11820\,
            I => \N__11817\
        );

    \I__1087\ : InMux
    port map (
            O => \N__11817\,
            I => \N__11814\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__11814\,
            I => \N__11811\
        );

    \I__1085\ : Span4Mux_h
    port map (
            O => \N__11811\,
            I => \N__11808\
        );

    \I__1084\ : Odrv4
    port map (
            O => \N__11808\,
            I => \M_this_vga_signals_address_5\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__11805\,
            I => \N__11802\
        );

    \I__1082\ : InMux
    port map (
            O => \N__11802\,
            I => \N__11799\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__11799\,
            I => \M_this_vga_signals_address_2\
        );

    \I__1080\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11793\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__11793\,
            I => \N__11790\
        );

    \I__1078\ : Odrv4
    port map (
            O => \N__11790\,
            I => \N_816_0\
        );

    \I__1077\ : InMux
    port map (
            O => \N__11787\,
            I => \N__11784\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__11784\,
            I => \N__11780\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__11783\,
            I => \N__11777\
        );

    \I__1074\ : Span4Mux_v
    port map (
            O => \N__11780\,
            I => \N__11774\
        );

    \I__1073\ : InMux
    port map (
            O => \N__11777\,
            I => \N__11771\
        );

    \I__1072\ : Odrv4
    port map (
            O => \N__11774\,
            I => \this_vga_ramdac.N_2612_reto\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__11771\,
            I => \this_vga_ramdac.N_2612_reto\
        );

    \I__1070\ : CascadeMux
    port map (
            O => \N__11766\,
            I => \N__11763\
        );

    \I__1069\ : CascadeBuf
    port map (
            O => \N__11763\,
            I => \N__11760\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__11760\,
            I => \N__11757\
        );

    \I__1067\ : InMux
    port map (
            O => \N__11757\,
            I => \N__11754\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__11754\,
            I => \N__11750\
        );

    \I__1065\ : InMux
    port map (
            O => \N__11753\,
            I => \N__11747\
        );

    \I__1064\ : Span4Mux_v
    port map (
            O => \N__11750\,
            I => \N__11744\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__11747\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__11744\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__11739\,
            I => \N__11736\
        );

    \I__1060\ : CascadeBuf
    port map (
            O => \N__11736\,
            I => \N__11733\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__11733\,
            I => \N__11730\
        );

    \I__1058\ : InMux
    port map (
            O => \N__11730\,
            I => \N__11727\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__11727\,
            I => \N__11723\
        );

    \I__1056\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11720\
        );

    \I__1055\ : Span4Mux_v
    port map (
            O => \N__11723\,
            I => \N__11717\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__11720\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__1053\ : Odrv4
    port map (
            O => \N__11717\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__1052\ : InMux
    port map (
            O => \N__11712\,
            I => \un1_M_this_map_address_q_cry_0\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__11709\,
            I => \N__11706\
        );

    \I__1050\ : CascadeBuf
    port map (
            O => \N__11706\,
            I => \N__11703\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__11703\,
            I => \N__11700\
        );

    \I__1048\ : InMux
    port map (
            O => \N__11700\,
            I => \N__11696\
        );

    \I__1047\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11693\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__11696\,
            I => \N__11690\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__11693\,
            I => \N__11685\
        );

    \I__1044\ : Span4Mux_v
    port map (
            O => \N__11690\,
            I => \N__11685\
        );

    \I__1043\ : Odrv4
    port map (
            O => \N__11685\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__1042\ : InMux
    port map (
            O => \N__11682\,
            I => \un1_M_this_map_address_q_cry_1\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__11679\,
            I => \N__11676\
        );

    \I__1040\ : CascadeBuf
    port map (
            O => \N__11676\,
            I => \N__11673\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__11673\,
            I => \N__11670\
        );

    \I__1038\ : InMux
    port map (
            O => \N__11670\,
            I => \N__11666\
        );

    \I__1037\ : InMux
    port map (
            O => \N__11669\,
            I => \N__11663\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__11666\,
            I => \N__11660\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__11663\,
            I => \N__11655\
        );

    \I__1034\ : Span4Mux_v
    port map (
            O => \N__11660\,
            I => \N__11655\
        );

    \I__1033\ : Odrv4
    port map (
            O => \N__11655\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__1032\ : InMux
    port map (
            O => \N__11652\,
            I => \un1_M_this_map_address_q_cry_2\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__11649\,
            I => \N__11646\
        );

    \I__1030\ : CascadeBuf
    port map (
            O => \N__11646\,
            I => \N__11643\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__11643\,
            I => \N__11640\
        );

    \I__1028\ : InMux
    port map (
            O => \N__11640\,
            I => \N__11637\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__11637\,
            I => \N__11633\
        );

    \I__1026\ : InMux
    port map (
            O => \N__11636\,
            I => \N__11630\
        );

    \I__1025\ : Span4Mux_v
    port map (
            O => \N__11633\,
            I => \N__11627\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__11630\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__1023\ : Odrv4
    port map (
            O => \N__11627\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__1022\ : InMux
    port map (
            O => \N__11622\,
            I => \un1_M_this_map_address_q_cry_3\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__11619\,
            I => \N__11616\
        );

    \I__1020\ : CascadeBuf
    port map (
            O => \N__11616\,
            I => \N__11613\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__11613\,
            I => \N__11610\
        );

    \I__1018\ : InMux
    port map (
            O => \N__11610\,
            I => \N__11607\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__11607\,
            I => \N__11603\
        );

    \I__1016\ : InMux
    port map (
            O => \N__11606\,
            I => \N__11600\
        );

    \I__1015\ : Span4Mux_v
    port map (
            O => \N__11603\,
            I => \N__11597\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__11600\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__1013\ : Odrv4
    port map (
            O => \N__11597\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__1012\ : InMux
    port map (
            O => \N__11592\,
            I => \un1_M_this_map_address_q_cry_4\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__11589\,
            I => \N__11586\
        );

    \I__1010\ : CascadeBuf
    port map (
            O => \N__11586\,
            I => \N__11583\
        );

    \I__1009\ : CascadeMux
    port map (
            O => \N__11583\,
            I => \N__11580\
        );

    \I__1008\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11577\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__11577\,
            I => \N__11573\
        );

    \I__1006\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11570\
        );

    \I__1005\ : Span4Mux_v
    port map (
            O => \N__11573\,
            I => \N__11567\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__11570\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__11567\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__1002\ : InMux
    port map (
            O => \N__11562\,
            I => \un1_M_this_map_address_q_cry_5\
        );

    \I__1001\ : InMux
    port map (
            O => \N__11559\,
            I => \N__11556\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__11556\,
            I => \N__11553\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__11553\,
            I => \M_this_oam_ram_write_data_0\
        );

    \I__998\ : InMux
    port map (
            O => \N__11550\,
            I => \N__11547\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__11547\,
            I => \N__11544\
        );

    \I__996\ : Span4Mux_h
    port map (
            O => \N__11544\,
            I => \N__11541\
        );

    \I__995\ : Odrv4
    port map (
            O => \N__11541\,
            I => \this_oam_ram.M_this_oam_ram_read_data_12\
        );

    \I__994\ : InMux
    port map (
            O => \N__11538\,
            I => \N__11535\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__11535\,
            I => \this_oam_ram.M_this_oam_ram_read_data_17\
        );

    \I__992\ : InMux
    port map (
            O => \N__11532\,
            I => \N__11529\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__11529\,
            I => \M_this_oam_ram_read_data_i_17\
        );

    \I__990\ : InMux
    port map (
            O => \N__11526\,
            I => \N__11523\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__11523\,
            I => \this_oam_ram.M_this_oam_ram_read_data_18\
        );

    \I__988\ : InMux
    port map (
            O => \N__11520\,
            I => \N__11517\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__11517\,
            I => \M_this_oam_ram_read_data_i_18\
        );

    \I__986\ : InMux
    port map (
            O => \N__11514\,
            I => \N__11511\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__11511\,
            I => \this_oam_ram.M_this_oam_ram_read_data_20\
        );

    \I__984\ : InMux
    port map (
            O => \N__11508\,
            I => \N__11505\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__11505\,
            I => \M_this_oam_ram_read_data_i_20\
        );

    \I__982\ : InMux
    port map (
            O => \N__11502\,
            I => \N__11496\
        );

    \I__981\ : InMux
    port map (
            O => \N__11501\,
            I => \N__11496\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__11496\,
            I => \this_pixel_clk_M_counter_q_i_1\
        );

    \I__979\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11486\
        );

    \I__978\ : InMux
    port map (
            O => \N__11492\,
            I => \N__11486\
        );

    \I__977\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11483\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__11486\,
            I => \N__11480\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__11483\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__974\ : Odrv4
    port map (
            O => \N__11480\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__973\ : IoInMux
    port map (
            O => \N__11475\,
            I => \N__11472\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__11472\,
            I => \N__11469\
        );

    \I__971\ : Span12Mux_s8_h
    port map (
            O => \N__11469\,
            I => \N__11466\
        );

    \I__970\ : Odrv12
    port map (
            O => \N__11466\,
            I => rgb_c_1
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__11463\,
            I => \N__11460\
        );

    \I__968\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11457\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__11457\,
            I => \N__11454\
        );

    \I__966\ : Span4Mux_v
    port map (
            O => \N__11454\,
            I => \N__11451\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__11451\,
            I => \M_this_vga_signals_address_1\
        );

    \I__964\ : InMux
    port map (
            O => \N__11448\,
            I => \this_ppu.un3_sprites_addr_cry_0\
        );

    \I__963\ : InMux
    port map (
            O => \N__11445\,
            I => \this_ppu.un3_sprites_addr_cry_1\
        );

    \I__962\ : InMux
    port map (
            O => \N__11442\,
            I => \N__11439\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__11439\,
            I => \N__11436\
        );

    \I__960\ : Odrv4
    port map (
            O => \N__11436\,
            I => \M_this_oam_ram_read_data_i_19\
        );

    \I__959\ : InMux
    port map (
            O => \N__11433\,
            I => \this_ppu.un3_sprites_addr_cry_2\
        );

    \I__958\ : InMux
    port map (
            O => \N__11430\,
            I => \this_ppu.un3_sprites_addr_cry_3\
        );

    \I__957\ : InMux
    port map (
            O => \N__11427\,
            I => \this_ppu.un3_sprites_addr_cry_4\
        );

    \I__956\ : InMux
    port map (
            O => \N__11424\,
            I => \this_ppu.un3_sprites_addr_cry_5\
        );

    \I__955\ : CascadeMux
    port map (
            O => \N__11421\,
            I => \N__11418\
        );

    \I__954\ : InMux
    port map (
            O => \N__11418\,
            I => \N__11415\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__11415\,
            I => \N__11412\
        );

    \I__952\ : Odrv4
    port map (
            O => \N__11412\,
            I => \M_this_oam_ram_read_data_23\
        );

    \I__951\ : InMux
    port map (
            O => \N__11409\,
            I => \this_ppu.un3_sprites_addr_cry_6\
        );

    \I__950\ : InMux
    port map (
            O => \N__11406\,
            I => \N__11403\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__11403\,
            I => \this_oam_ram.M_this_oam_ram_read_data_21\
        );

    \I__948\ : InMux
    port map (
            O => \N__11400\,
            I => \N__11397\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__11397\,
            I => \M_this_oam_ram_read_data_i_21\
        );

    \I__946\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11391\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__11391\,
            I => \N__11388\
        );

    \I__944\ : Odrv4
    port map (
            O => \N__11388\,
            I => \M_this_oam_ram_write_data_4\
        );

    \I__943\ : InMux
    port map (
            O => \N__11385\,
            I => \N__11382\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__11382\,
            I => \N__11379\
        );

    \I__941\ : Odrv4
    port map (
            O => \N__11379\,
            I => \N_895_0\
        );

    \I__940\ : InMux
    port map (
            O => \N__11376\,
            I => \N__11373\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__11373\,
            I => \N__11370\
        );

    \I__938\ : Odrv4
    port map (
            O => \N__11370\,
            I => \N_891_0\
        );

    \I__937\ : InMux
    port map (
            O => \N__11367\,
            I => \N__11364\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__11364\,
            I => \this_oam_ram.M_this_oam_ram_read_data_10\
        );

    \I__935\ : InMux
    port map (
            O => \N__11361\,
            I => \N__11358\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__11358\,
            I => \this_oam_ram.M_this_oam_ram_read_data_11\
        );

    \I__933\ : InMux
    port map (
            O => \N__11355\,
            I => \N__11352\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__11352\,
            I => \M_this_oam_ram_write_data_28\
        );

    \I__931\ : InMux
    port map (
            O => \N__11349\,
            I => \N__11346\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__11346\,
            I => \N__11343\
        );

    \I__929\ : Odrv4
    port map (
            O => \N__11343\,
            I => \N_894_0\
        );

    \I__928\ : InMux
    port map (
            O => \N__11340\,
            I => \N__11337\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__11337\,
            I => \N_889_0\
        );

    \I__926\ : InMux
    port map (
            O => \N__11334\,
            I => \N__11331\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__11331\,
            I => \this_ppu.M_this_oam_ram_read_data_i_16\
        );

    \I__924\ : IoInMux
    port map (
            O => \N__11328\,
            I => \N__11325\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__11325\,
            I => \N__11322\
        );

    \I__922\ : Span12Mux_s2_h
    port map (
            O => \N__11322\,
            I => \N__11319\
        );

    \I__921\ : Odrv12
    port map (
            O => \N__11319\,
            I => rgb_c_3
        );

    \I__920\ : IoInMux
    port map (
            O => \N__11316\,
            I => \N__11313\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__11313\,
            I => \N__11310\
        );

    \I__918\ : Span4Mux_s3_h
    port map (
            O => \N__11310\,
            I => \N__11307\
        );

    \I__917\ : Span4Mux_v
    port map (
            O => \N__11307\,
            I => \N__11304\
        );

    \I__916\ : Odrv4
    port map (
            O => \N__11304\,
            I => rgb_c_4
        );

    \I__915\ : InMux
    port map (
            O => \N__11301\,
            I => \N__11298\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__11298\,
            I => \N__11295\
        );

    \I__913\ : Span4Mux_h
    port map (
            O => \N__11295\,
            I => \N__11292\
        );

    \I__912\ : Odrv4
    port map (
            O => \N__11292\,
            I => \N_834_0\
        );

    \I__911\ : InMux
    port map (
            O => \N__11289\,
            I => \N__11286\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__11286\,
            I => \N__11283\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__11283\,
            I => \N_818_0\
        );

    \I__908\ : InMux
    port map (
            O => \N__11280\,
            I => \N__11277\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__11277\,
            I => \N__11274\
        );

    \I__906\ : Span4Mux_v
    port map (
            O => \N__11274\,
            I => \N__11271\
        );

    \I__905\ : Odrv4
    port map (
            O => \N__11271\,
            I => \N_837_0\
        );

    \I__904\ : InMux
    port map (
            O => \N__11268\,
            I => \N__11265\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__11265\,
            I => \N__11262\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__11262\,
            I => \M_this_oam_ram_write_data_5\
        );

    \I__901\ : InMux
    port map (
            O => \N__11259\,
            I => \N__11256\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__11256\,
            I => \M_this_oam_ram_write_data_8\
        );

    \I__899\ : InMux
    port map (
            O => \N__11253\,
            I => \N__11250\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__11250\,
            I => \N_836_0\
        );

    \I__897\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11244\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__11244\,
            I => \N_896_0\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__11241\,
            I => \N__11238\
        );

    \I__894\ : CascadeBuf
    port map (
            O => \N__11238\,
            I => \N__11235\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__11235\,
            I => \N__11232\
        );

    \I__892\ : InMux
    port map (
            O => \N__11232\,
            I => \N__11228\
        );

    \I__891\ : InMux
    port map (
            O => \N__11231\,
            I => \N__11225\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__11228\,
            I => \N__11222\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__11225\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__888\ : Odrv4
    port map (
            O => \N__11222\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__887\ : InMux
    port map (
            O => \N__11217\,
            I => \un1_M_this_oam_address_q_cry_3\
        );

    \I__886\ : InMux
    port map (
            O => \N__11214\,
            I => \un1_M_this_oam_address_q_cry_4\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__11211\,
            I => \N__11208\
        );

    \I__884\ : CascadeBuf
    port map (
            O => \N__11208\,
            I => \N__11205\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__11205\,
            I => \N__11202\
        );

    \I__882\ : InMux
    port map (
            O => \N__11202\,
            I => \N__11199\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__11199\,
            I => \N__11195\
        );

    \I__880\ : InMux
    port map (
            O => \N__11198\,
            I => \N__11192\
        );

    \I__879\ : Span4Mux_h
    port map (
            O => \N__11195\,
            I => \N__11189\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__11192\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__877\ : Odrv4
    port map (
            O => \N__11189\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__876\ : InMux
    port map (
            O => \N__11184\,
            I => \N__11181\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__11181\,
            I => \this_oam_ram.M_this_oam_ram_read_data_19\
        );

    \I__874\ : InMux
    port map (
            O => \N__11178\,
            I => \N__11175\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__11175\,
            I => \M_this_data_tmp_qZ0Z_26\
        );

    \I__872\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11169\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__11169\,
            I => \M_this_oam_ram_write_data_26\
        );

    \I__870\ : InMux
    port map (
            O => \N__11166\,
            I => \N__11163\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__11163\,
            I => \M_this_oam_ram_write_data_20\
        );

    \I__868\ : InMux
    port map (
            O => \N__11160\,
            I => \N__11157\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__11157\,
            I => \N_892_0\
        );

    \I__866\ : IoInMux
    port map (
            O => \N__11154\,
            I => \N__11151\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__11151\,
            I => \N__11148\
        );

    \I__864\ : Span12Mux_s6_h
    port map (
            O => \N__11148\,
            I => \N__11145\
        );

    \I__863\ : Span12Mux_v
    port map (
            O => \N__11145\,
            I => \N__11142\
        );

    \I__862\ : Odrv12
    port map (
            O => \N__11142\,
            I => rgb_c_0
        );

    \I__861\ : IoInMux
    port map (
            O => \N__11139\,
            I => \N__11136\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__11136\,
            I => \N__11133\
        );

    \I__859\ : Odrv12
    port map (
            O => \N__11133\,
            I => this_vga_signals_vvisibility_i
        );

    \I__858\ : InMux
    port map (
            O => \N__11130\,
            I => \N__11127\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__11127\,
            I => \this_delay_clk.M_pipe_qZ0Z_1\
        );

    \I__856\ : IoInMux
    port map (
            O => \N__11124\,
            I => \N__11121\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__11121\,
            I => \N__11118\
        );

    \I__854\ : Span4Mux_s1_h
    port map (
            O => \N__11118\,
            I => \N__11115\
        );

    \I__853\ : Span4Mux_h
    port map (
            O => \N__11115\,
            I => \N__11112\
        );

    \I__852\ : Odrv4
    port map (
            O => \N__11112\,
            I => rgb_c_2
        );

    \I__851\ : InMux
    port map (
            O => \N__11109\,
            I => \N__11106\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__11106\,
            I => \N__11103\
        );

    \I__849\ : Odrv12
    port map (
            O => \N__11103\,
            I => port_clk_c
        );

    \I__848\ : InMux
    port map (
            O => \N__11100\,
            I => \N__11097\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__11097\,
            I => \this_delay_clk.M_pipe_qZ0Z_0\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__11094\,
            I => \N__11091\
        );

    \I__845\ : CascadeBuf
    port map (
            O => \N__11091\,
            I => \N__11088\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__11088\,
            I => \N__11085\
        );

    \I__843\ : InMux
    port map (
            O => \N__11085\,
            I => \N__11082\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__11082\,
            I => \N__11078\
        );

    \I__841\ : InMux
    port map (
            O => \N__11081\,
            I => \N__11075\
        );

    \I__840\ : Span4Mux_v
    port map (
            O => \N__11078\,
            I => \N__11072\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__11075\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__11072\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__11067\,
            I => \N__11064\
        );

    \I__836\ : CascadeBuf
    port map (
            O => \N__11064\,
            I => \N__11061\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__11061\,
            I => \N__11058\
        );

    \I__834\ : InMux
    port map (
            O => \N__11058\,
            I => \N__11055\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__11055\,
            I => \N__11051\
        );

    \I__832\ : InMux
    port map (
            O => \N__11054\,
            I => \N__11048\
        );

    \I__831\ : Span4Mux_v
    port map (
            O => \N__11051\,
            I => \N__11045\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__11048\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__829\ : Odrv4
    port map (
            O => \N__11045\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__828\ : InMux
    port map (
            O => \N__11040\,
            I => \un1_M_this_oam_address_q_cry_0\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__11037\,
            I => \N__11034\
        );

    \I__826\ : CascadeBuf
    port map (
            O => \N__11034\,
            I => \N__11031\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__11031\,
            I => \N__11028\
        );

    \I__824\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11024\
        );

    \I__823\ : InMux
    port map (
            O => \N__11027\,
            I => \N__11021\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__11024\,
            I => \N__11018\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__11021\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__11018\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__819\ : InMux
    port map (
            O => \N__11013\,
            I => \un1_M_this_oam_address_q_cry_1\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__11010\,
            I => \N__11007\
        );

    \I__817\ : CascadeBuf
    port map (
            O => \N__11007\,
            I => \N__11004\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__11004\,
            I => \N__11001\
        );

    \I__815\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10998\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__10998\,
            I => \N__10994\
        );

    \I__813\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10991\
        );

    \I__812\ : Span4Mux_h
    port map (
            O => \N__10994\,
            I => \N__10988\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__10991\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__810\ : Odrv4
    port map (
            O => \N__10988\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__809\ : InMux
    port map (
            O => \N__10983\,
            I => \un1_M_this_oam_address_q_cry_2\
        );

    \I__808\ : IoInMux
    port map (
            O => \N__10980\,
            I => \N__10977\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__10977\,
            I => \N__10974\
        );

    \I__806\ : Span4Mux_s3_h
    port map (
            O => \N__10974\,
            I => \N__10971\
        );

    \I__805\ : Span4Mux_v
    port map (
            O => \N__10971\,
            I => \N__10968\
        );

    \I__804\ : Odrv4
    port map (
            O => \N__10968\,
            I => port_nmib_0_i
        );

    \IN_MUX_bfv_23_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_17_0_\
        );

    \IN_MUX_bfv_23_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_sprites_address_q_cry_7\,
            carryinitout => \bfn_23_18_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_12_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_12_22_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_24_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_21_0_\
        );

    \IN_MUX_bfv_24_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \M_this_data_count_q_cry_7\,
            carryinitout => \bfn_24_22_0_\
        );

    \IN_MUX_bfv_21_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_20_0_\
        );

    \IN_MUX_bfv_21_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            carryinitout => \bfn_21_21_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_17_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_map_address_q_cry_7\,
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_26_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_26_23_0_\
        );

    \IN_MUX_bfv_26_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \M_this_external_address_q_cry_7\,
            carryinitout => \bfn_26_24_0_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI4KCU6_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__16548\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_1358_g\
        );

    \this_reset_cond.M_stage_q_RNIC5C7_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__15809\,
            GLOBALBUFFEROUTPUT => \M_this_reset_cond_out_g_0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI0JAO7_9_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17735\,
            in2 => \_gnd_net_\,
            in3 => \N__15879\,
            lcout => port_nmib_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_0_9_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15872\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => this_vga_signals_vvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_1_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11100\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32633\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_2_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11130\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32633\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11787\,
            in2 => \_gnd_net_\,
            in3 => \N__11895\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_0_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11109\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32636\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_0_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26788\,
            in1 => \N__11081\,
            in2 => \N__18624\,
            in3 => \N__18619\,
            lcout => \M_this_oam_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => \un1_M_this_oam_address_q_cry_0\,
            clk => \N__32616\,
            ce => 'H',
            sr => \N__26071\
        );

    \M_this_oam_address_q_1_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26792\,
            in1 => \N__11054\,
            in2 => \_gnd_net_\,
            in3 => \N__11040\,
            lcout => \M_this_oam_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_oam_address_q_cry_0\,
            carryout => \un1_M_this_oam_address_q_cry_1\,
            clk => \N__32616\,
            ce => 'H',
            sr => \N__26071\
        );

    \M_this_oam_address_q_2_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26789\,
            in1 => \N__11027\,
            in2 => \_gnd_net_\,
            in3 => \N__11013\,
            lcout => \M_this_oam_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_oam_address_q_cry_1\,
            carryout => \un1_M_this_oam_address_q_cry_2\,
            clk => \N__32616\,
            ce => 'H',
            sr => \N__26071\
        );

    \M_this_oam_address_q_3_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26793\,
            in1 => \N__10997\,
            in2 => \_gnd_net_\,
            in3 => \N__10983\,
            lcout => \M_this_oam_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_oam_address_q_cry_2\,
            carryout => \un1_M_this_oam_address_q_cry_3\,
            clk => \N__32616\,
            ce => 'H',
            sr => \N__26071\
        );

    \M_this_oam_address_q_4_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26790\,
            in1 => \N__11231\,
            in2 => \_gnd_net_\,
            in3 => \N__11217\,
            lcout => \M_this_oam_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_oam_address_q_cry_3\,
            carryout => \un1_M_this_oam_address_q_cry_4\,
            clk => \N__32616\,
            ce => 'H',
            sr => \N__26071\
        );

    \M_this_oam_address_q_5_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__11198\,
            in1 => \N__26791\,
            in2 => \_gnd_net_\,
            in3 => \N__11214\,
            lcout => \M_this_oam_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32616\,
            ce => 'H',
            sr => \N__26071\
        );

    \M_this_data_tmp_q_esr_26_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32919\,
            lcout => \M_this_data_tmp_qZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32620\,
            ce => \N__17664\,
            sr => \N__26070\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11184\,
            lcout => \M_this_oam_ram_read_data_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_26_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11178\,
            in2 => \_gnd_net_\,
            in3 => \N__18618\,
            lcout => \M_this_oam_ram_write_data_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_20_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12321\,
            in2 => \_gnd_net_\,
            in3 => \N__18617\,
            lcout => \M_this_oam_ram_write_data_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_23_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12300\,
            lcout => \N_892_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_0_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11491\,
            lcout => \this_pixel_clk_M_counter_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32637\,
            ce => 'H',
            sr => \N__26064\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11891\,
            in2 => \_gnd_net_\,
            in3 => \N__12351\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11884\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12648\,
            lcout => rgb_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11874\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12384\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_15_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18576\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12057\,
            lcout => \N_834_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_14_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12774\,
            in2 => \_gnd_net_\,
            in3 => \N__18575\,
            lcout => \N_818_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_1_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13644\,
            in2 => \_gnd_net_\,
            in3 => \N__18592\,
            lcout => \N_837_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_5_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13296\,
            in2 => \_gnd_net_\,
            in3 => \N__18591\,
            lcout => \M_this_oam_ram_write_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_8_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12051\,
            in2 => \_gnd_net_\,
            in3 => \N__18597\,
            lcout => \M_this_oam_ram_write_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_7_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__18601\,
            in1 => \N__12747\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_836_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_11_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12045\,
            in2 => \_gnd_net_\,
            in3 => \N__18598\,
            lcout => \N_896_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_4_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12732\,
            in2 => \_gnd_net_\,
            in3 => \N__18596\,
            lcout => \M_this_oam_ram_write_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_13_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18599\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13497\,
            lcout => \N_895_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_27_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12765\,
            in2 => \_gnd_net_\,
            in3 => \N__18600\,
            lcout => \N_891_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11367\,
            lcout => \M_this_oam_ram_read_data_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_0_RNISG75_1_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11361\,
            lcout => \M_this_oam_ram_read_data_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_28_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12930\,
            in2 => \_gnd_net_\,
            in3 => \N__18608\,
            lcout => \M_this_oam_ram_write_data_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_19_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18609\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12201\,
            lcout => \N_894_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_31_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12717\,
            in2 => \_gnd_net_\,
            in3 => \N__18610\,
            lcout => \N_889_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un3_sprites_addr_cry_0_c_inv_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11334\,
            in2 => \N__19318\,
            in3 => \N__12902\,
            lcout => \this_ppu.M_this_oam_ram_read_data_i_16\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \this_ppu.un3_sprites_addr_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un3_sprites_addr_cry_0_c_RNIRLA8_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11532\,
            in2 => \N__20926\,
            in3 => \N__11448\,
            lcout => \this_ppu.un3_sprites_addr_cry_0_c_RNIRLAZ0Z8\,
            ltout => OPEN,
            carryin => \this_ppu.un3_sprites_addr_cry_0\,
            carryout => \this_ppu.un3_sprites_addr_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un3_sprites_addr_cry_1_c_RNITOB8_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11520\,
            in2 => \N__13880\,
            in3 => \N__11445\,
            lcout => \this_ppu.un3_sprites_addr_cry_1_c_RNITOBZ0Z8\,
            ltout => OPEN,
            carryin => \this_ppu.un3_sprites_addr_cry_1\,
            carryout => \this_ppu.un3_sprites_addr_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un3_sprites_addr_cry_2_c_RNIVRC8_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11442\,
            in2 => \N__13945\,
            in3 => \N__11433\,
            lcout => \this_ppu.un3_sprites_addr_cry_2_c_RNIVRCZ0Z8\,
            ltout => OPEN,
            carryin => \this_ppu.un3_sprites_addr_cry_2\,
            carryout => \this_ppu.un3_sprites_addr_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un3_sprites_addr_cry_3_c_RNI1VD8_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11508\,
            in2 => \N__13813\,
            in3 => \N__11430\,
            lcout => \this_ppu.un3_sprites_addr_cry_3_c_RNI1VDZ0Z8\,
            ltout => OPEN,
            carryin => \this_ppu.un3_sprites_addr_cry_3\,
            carryout => \this_ppu.un3_sprites_addr_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un3_sprites_addr_cry_4_c_RNI32F8_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11400\,
            in2 => \N__13576\,
            in3 => \N__11427\,
            lcout => \this_ppu.un3_sprites_addr_cry_4_c_RNI32FZ0Z8\,
            ltout => OPEN,
            carryin => \this_ppu.un3_sprites_addr_cry_4\,
            carryout => \this_ppu.un3_sprites_addr_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un3_sprites_addr_cry_5_c_RNI55G8_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12878\,
            in2 => \N__12279\,
            in3 => \N__11424\,
            lcout => \this_ppu.un3_sprites_addr_cry_5_c_RNI55GZ0Z8\,
            ltout => OPEN,
            carryin => \this_ppu.un3_sprites_addr_cry_5\,
            carryout => \this_ppu.un3_sprites_addr_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un3_sprites_addr_cry_6_c_RNIP5L8_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__12827\,
            in1 => \_gnd_net_\,
            in2 => \N__11421\,
            in3 => \N__11409\,
            lcout => \this_ppu.un3_sprites_addr_cry_6_c_RNIP5LZ0Z8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m2_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22928\,
            in2 => \_gnd_net_\,
            in3 => \N__21578\,
            lcout => \this_vga_signals.if_m2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_3_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11406\,
            lcout => \M_this_oam_ram_read_data_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_0_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13479\,
            in2 => \_gnd_net_\,
            in3 => \N__18623\,
            lcout => \M_this_oam_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_0_RNISG75_2_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11550\,
            lcout => \M_this_oam_ram_read_data_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11538\,
            lcout => \M_this_oam_ram_read_data_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11526\,
            lcout => \M_this_oam_ram_read_data_i_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11514\,
            lcout => \M_this_oam_ram_read_data_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_1_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__11502\,
            in1 => \N__11493\,
            in2 => \_gnd_net_\,
            in3 => \N__26181\,
            lcout => \this_pixel_clk_M_counter_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32630\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.G_442_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__11501\,
            in1 => \N__11492\,
            in2 => \_gnd_net_\,
            in3 => \N__26180\,
            lcout => \G_442\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12363\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11883\,
            lcout => rgb_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI946123_9_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__13146\,
            in1 => \N__17129\,
            in2 => \_gnd_net_\,
            in3 => \N__13131\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI6B7F1_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32896\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19891\,
            lcout => \N_816_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__11904\,
            in1 => \N__15822\,
            in2 => \N__11783\,
            in3 => \N__12670\,
            lcout => \this_vga_ramdac.N_2612_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32638\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_0_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24041\,
            in1 => \N__11753\,
            in2 => \N__19896\,
            in3 => \N__19887\,
            lcout => \M_this_map_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \un1_M_this_map_address_q_cry_0\,
            clk => \N__32643\,
            ce => 'H',
            sr => \N__26050\
        );

    \M_this_map_address_q_1_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24046\,
            in1 => \N__11726\,
            in2 => \_gnd_net_\,
            in3 => \N__11712\,
            lcout => \M_this_map_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_0\,
            carryout => \un1_M_this_map_address_q_cry_1\,
            clk => \N__32643\,
            ce => 'H',
            sr => \N__26050\
        );

    \M_this_map_address_q_2_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24042\,
            in1 => \N__11699\,
            in2 => \_gnd_net_\,
            in3 => \N__11682\,
            lcout => \M_this_map_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_1\,
            carryout => \un1_M_this_map_address_q_cry_2\,
            clk => \N__32643\,
            ce => 'H',
            sr => \N__26050\
        );

    \M_this_map_address_q_3_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24047\,
            in1 => \N__11669\,
            in2 => \_gnd_net_\,
            in3 => \N__11652\,
            lcout => \M_this_map_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_2\,
            carryout => \un1_M_this_map_address_q_cry_3\,
            clk => \N__32643\,
            ce => 'H',
            sr => \N__26050\
        );

    \M_this_map_address_q_4_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24043\,
            in1 => \N__11636\,
            in2 => \_gnd_net_\,
            in3 => \N__11622\,
            lcout => \M_this_map_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_3\,
            carryout => \un1_M_this_map_address_q_cry_4\,
            clk => \N__32643\,
            ce => 'H',
            sr => \N__26050\
        );

    \M_this_map_address_q_5_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24048\,
            in1 => \N__11606\,
            in2 => \_gnd_net_\,
            in3 => \N__11592\,
            lcout => \M_this_map_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_4\,
            carryout => \un1_M_this_map_address_q_cry_5\,
            clk => \N__32643\,
            ce => 'H',
            sr => \N__26050\
        );

    \M_this_map_address_q_6_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24044\,
            in1 => \N__11576\,
            in2 => \_gnd_net_\,
            in3 => \N__11562\,
            lcout => \M_this_map_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_5\,
            carryout => \un1_M_this_map_address_q_cry_6\,
            clk => \N__32643\,
            ce => 'H',
            sr => \N__26050\
        );

    \M_this_map_address_q_7_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24045\,
            in1 => \N__11981\,
            in2 => \_gnd_net_\,
            in3 => \N__11967\,
            lcout => \M_this_map_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_6\,
            carryout => \un1_M_this_map_address_q_cry_7\,
            clk => \N__32643\,
            ce => 'H',
            sr => \N__26050\
        );

    \M_this_map_address_q_8_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24038\,
            in1 => \N__11951\,
            in2 => \_gnd_net_\,
            in3 => \N__11937\,
            lcout => \M_this_map_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_25_0_\,
            carryout => \un1_M_this_map_address_q_cry_8\,
            clk => \N__32647\,
            ce => 'H',
            sr => \N__26047\
        );

    \M_this_map_address_q_9_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__11918\,
            in1 => \N__24039\,
            in2 => \_gnd_net_\,
            in3 => \N__11934\,
            lcout => \M_this_map_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32647\,
            ce => 'H',
            sr => \N__26047\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111101"
        )
    port map (
            in0 => \N__12453\,
            in1 => \N__12496\,
            in2 => \N__12556\,
            in3 => \N__12583\,
            lcout => \this_vga_ramdac.i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_q_ret_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__15817\,
            in1 => \N__17128\,
            in2 => \N__11873\,
            in3 => \N__12681\,
            lcout => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32651\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12699\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11861\,
            lcout => rgb_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIAF7F1_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28191\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19897\,
            lcout => \N_60_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIT1827_9_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17119\,
            in2 => \_gnd_net_\,
            in3 => \N__13104\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI0MGR61_9_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17118\,
            in2 => \_gnd_net_\,
            in3 => \N__13179\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI7CFM8_9_LC_9_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17121\,
            in2 => \_gnd_net_\,
            in3 => \N__13053\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIPFB21_2_LC_9_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__12186\,
            in1 => \N__32119\,
            in2 => \N__31971\,
            in3 => \N__12174\,
            lcout => \M_this_ppu_sprites_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_15_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27907\,
            lcout => \M_this_data_tmp_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32560\,
            ce => \N__17357\,
            sr => \N__26069\
        );

    \M_this_data_tmp_q_esr_8_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28469\,
            lcout => \M_this_data_tmp_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32569\,
            ce => \N__17353\,
            sr => \N__26067\
        );

    \M_this_data_tmp_q_esr_11_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31356\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32569\,
            ce => \N__17353\,
            sr => \N__26067\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_9_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13488\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18582\,
            lcout => \N_835_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_3_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12753\,
            in2 => \_gnd_net_\,
            in3 => \N__18580\,
            lcout => \N_897_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_6_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18581\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14142\,
            lcout => \N_53_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_2_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12738\,
            in2 => \_gnd_net_\,
            in3 => \N__18578\,
            lcout => \M_this_oam_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_29_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18579\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13308\,
            lcout => \N_890_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_12_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13287\,
            in2 => \_gnd_net_\,
            in3 => \N__18577\,
            lcout => \M_this_oam_ram_write_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_25_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18590\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12723\,
            lcout => \N_831_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_24_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18587\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13635\,
            lcout => \M_this_oam_ram_write_data_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_22_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12306\,
            in2 => \_gnd_net_\,
            in3 => \N__18589\,
            lcout => \N_832_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_21_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18588\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12312\,
            lcout => \N_893_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_16_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28468\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32597\,
            ce => \N__15957\,
            sr => \N__26058\
        );

    \M_this_data_tmp_q_esr_18_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32908\,
            lcout => \M_this_data_tmp_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32597\,
            ce => \N__15957\,
            sr => \N__26058\
        );

    \M_this_data_tmp_q_esr_19_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31357\,
            lcout => \M_this_data_tmp_qZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32597\,
            ce => \N__15957\,
            sr => \N__26058\
        );

    \M_this_data_tmp_q_esr_20_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28266\,
            lcout => \M_this_data_tmp_qZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32597\,
            ce => \N__15957\,
            sr => \N__26058\
        );

    \M_this_data_tmp_q_esr_21_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24463\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32597\,
            ce => \N__15957\,
            sr => \N__26058\
        );

    \M_this_data_tmp_q_esr_22_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28190\,
            lcout => \M_this_data_tmp_qZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32597\,
            ce => \N__15957\,
            sr => \N__26058\
        );

    \M_this_data_tmp_q_esr_23_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27911\,
            lcout => \M_this_data_tmp_qZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32597\,
            ce => \N__15957\,
            sr => \N__26058\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_2_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011010010101"
        )
    port map (
            in0 => \N__12998\,
            in1 => \N__12411\,
            in2 => \N__14622\,
            in3 => \N__12974\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_4_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12288\,
            lcout => \M_this_oam_ram_read_data_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIUULS4_3_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__14480\,
            in1 => \_gnd_net_\,
            in2 => \N__14550\,
            in3 => \N__13041\,
            lcout => \this_vga_signals.M_hcounter_q_RNIUULS4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001111001001"
        )
    port map (
            in0 => \N__14481\,
            in1 => \N__13083\,
            in2 => \N__14551\,
            in3 => \N__13042\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101110001001"
        )
    port map (
            in0 => \N__14478\,
            in1 => \N__13082\,
            in2 => \N__14549\,
            in3 => \N__13039\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__13040\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14479\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1\,
            ltout => \this_vga_signals.mult1_un68_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m2_0_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__14535\,
            in1 => \N__13390\,
            in2 => \N__12414\,
            in3 => \N__13364\,
            lcout => \this_vga_signals.if_m2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIBG7F1_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27912\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19868\,
            lcout => \N_58_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNIR5V44_0_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21497\,
            in1 => \N__13708\,
            in2 => \_gnd_net_\,
            in3 => \N__13248\,
            lcout => \N_3_0\,
            ltout => \N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.G_480_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12708\,
            in2 => \N__12390\,
            in3 => \N__12330\,
            lcout => \G_480\,
            ltout => \G_480_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__12380\,
            in1 => \N__12612\,
            in2 => \N__12387\,
            in3 => \N__15814\,
            lcout => \this_vga_ramdac.N_2614_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001001110"
        )
    port map (
            in0 => \N__12669\,
            in1 => \N__12362\,
            in2 => \N__15821\,
            in3 => \N__12423\,
            lcout => \this_vga_ramdac.N_2611_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__12621\,
            in1 => \N__15810\,
            in2 => \N__12347\,
            in3 => \N__12668\,
            lcout => \this_vga_ramdac.N_2610_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_RNIIQFU3_1_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000010101010"
        )
    port map (
            in0 => \N__13732\,
            in1 => \N__21663\,
            in2 => \N__13710\,
            in3 => \N__21496\,
            lcout => \N_2_0\,
            ltout => \N_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_2_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12324\,
            in3 => \N__13260\,
            lcout => \M_this_vga_signals_pixel_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100100101"
        )
    port map (
            in0 => \N__12462\,
            in1 => \N__12505\,
            in2 => \N__12558\,
            in3 => \N__12603\,
            lcout => OPEN,
            ltout => \this_vga_ramdac.i2_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100000010"
        )
    port map (
            in0 => \N__12680\,
            in1 => \N__15816\,
            in2 => \N__12702\,
            in3 => \N__12695\,
            lcout => \this_vga_ramdac.N_2615_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32639\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101100010111"
        )
    port map (
            in0 => \N__12602\,
            in1 => \N__12552\,
            in2 => \N__12507\,
            in3 => \N__12461\,
            lcout => OPEN,
            ltout => \this_vga_ramdac.m16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__12644\,
            in1 => \N__15815\,
            in2 => \N__12684\,
            in3 => \N__12679\,
            lcout => \this_vga_ramdac.N_2613_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32639\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI497F1_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28395\,
            in2 => \_gnd_net_\,
            in3 => \N__19883\,
            lcout => \N_73_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100010"
        )
    port map (
            in0 => \N__12551\,
            in1 => \N__12501\,
            in2 => \_gnd_net_\,
            in3 => \N__12601\,
            lcout => \this_vga_ramdac.N_24_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010100101011"
        )
    port map (
            in0 => \N__12454\,
            in1 => \N__12497\,
            in2 => \N__12557\,
            in3 => \N__12592\,
            lcout => \this_vga_ramdac.m19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111101111"
        )
    port map (
            in0 => \N__12593\,
            in1 => \N__12550\,
            in2 => \N__12506\,
            in3 => \N__12455\,
            lcout => \this_vga_ramdac.m6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_14_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28179\,
            lcout => \M_this_data_tmp_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32549\,
            ce => \N__17361\,
            sr => \N__26068\
        );

    \M_this_data_tmp_q_esr_27_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31359\,
            lcout => \M_this_data_tmp_qZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32561\,
            ce => \N__17645\,
            sr => \N__26065\
        );

    \M_this_data_tmp_q_esr_30_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28189\,
            lcout => \M_this_data_tmp_qZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32561\,
            ce => \N__17645\,
            sr => \N__26065\
        );

    \M_this_data_tmp_q_esr_3_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31358\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32570\,
            ce => \N__16521\,
            sr => \N__26062\
        );

    \M_this_data_tmp_q_esr_7_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27945\,
            lcout => \M_this_data_tmp_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32570\,
            ce => \N__16521\,
            sr => \N__26062\
        );

    \M_this_data_tmp_q_esr_2_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32915\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32570\,
            ce => \N__16521\,
            sr => \N__26062\
        );

    \M_this_data_tmp_q_esr_4_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32570\,
            ce => \N__16521\,
            sr => \N__26062\
        );

    \M_this_data_tmp_q_esr_25_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30928\,
            lcout => \M_this_data_tmp_qZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32580\,
            ce => \N__17659\,
            sr => \N__26059\
        );

    \M_this_data_tmp_q_esr_31_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27937\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32580\,
            ce => \N__17659\,
            sr => \N__26059\
        );

    \M_this_data_tmp_q_esr_28_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28326\,
            lcout => \M_this_data_tmp_qZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32580\,
            ce => \N__17659\,
            sr => \N__26059\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_17_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18585\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15396\,
            lcout => \N_833_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI98B5_0_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19311\,
            in2 => \_gnd_net_\,
            in3 => \N__12909\,
            lcout => \this_ppu.un3_sprites_addr_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNIIT3_6_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13604\,
            lcout => \M_this_ppu_vram_addr_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_18_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18584\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12861\,
            lcout => \M_this_oam_ram_write_data_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI5S7_7_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13605\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13526\,
            lcout => \M_this_ppu_map_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_i_30_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__18586\,
            in1 => \N__12810\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_830_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_16_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12792\,
            in2 => \_gnd_net_\,
            in3 => \N__18583\,
            lcout => \M_this_oam_ram_write_data_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIB0ACH_2_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13363\,
            in1 => \N__14612\,
            in2 => \N__13394\,
            in3 => \N__14552\,
            lcout => \this_vga_signals.d_N_3_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13386\,
            in2 => \_gnd_net_\,
            in3 => \N__13362\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m4_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001100000"
        )
    port map (
            in0 => \N__14599\,
            in1 => \N__14798\,
            in2 => \N__13011\,
            in3 => \N__14553\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_i4_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__12997\,
            in1 => \N__13008\,
            in2 => \N__13002\,
            in3 => \N__12947\,
            lcout => \this_vga_signals.mult1_un82_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100110100110"
        )
    port map (
            in0 => \N__12999\,
            in1 => \N__12981\,
            in2 => \N__12960\,
            in3 => \N__12975\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c2_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100000101"
        )
    port map (
            in0 => \N__14799\,
            in1 => \_gnd_net_\,
            in2 => \N__12963\,
            in3 => \N__14600\,
            lcout => \this_vga_signals.mult1_un82_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m2_2_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001001000"
        )
    port map (
            in0 => \N__14547\,
            in1 => \N__14473\,
            in2 => \N__14613\,
            in3 => \N__13049\,
            lcout => \this_vga_signals.if_m2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_1_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13278\,
            in1 => \N__14351\,
            in2 => \N__14419\,
            in3 => \N__13038\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110101001011"
        )
    port map (
            in0 => \N__13094\,
            in1 => \N__14475\,
            in2 => \N__12951\,
            in3 => \N__14410\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_ac0_3_0_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001111000001"
        )
    port map (
            in0 => \N__14848\,
            in1 => \N__13152\,
            in2 => \N__14807\,
            in3 => \N__13112\,
            lcout => \this_vga_signals.mult1_un89_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13113\,
            in1 => \N__12948\,
            in2 => \N__13172\,
            in3 => \N__12936\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un89_sum_axbxc3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI6DOUP9_9_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__17120\,
            in1 => \_gnd_net_\,
            in2 => \N__13206\,
            in3 => \N__13203\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axb1_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14607\,
            in2 => \_gnd_net_\,
            in3 => \N__13165\,
            lcout => \this_vga_signals.mult1_un82_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13142\,
            in2 => \_gnd_net_\,
            in3 => \N__13124\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111010001100"
        )
    port map (
            in0 => \N__13276\,
            in1 => \N__13064\,
            in2 => \N__14418\,
            in3 => \N__14349\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000110000011"
        )
    port map (
            in0 => \N__14350\,
            in1 => \N__14406\,
            in2 => \N__13068\,
            in3 => \N__13277\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010111101"
        )
    port map (
            in0 => \N__14225\,
            in1 => \N__14170\,
            in2 => \N__14291\,
            in3 => \N__14346\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9\,
            ltout => \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_1_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101110"
        )
    port map (
            in0 => \N__14348\,
            in1 => \N__14401\,
            in2 => \N__13074\,
            in3 => \N__13275\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101000011010"
        )
    port map (
            in0 => \N__14402\,
            in1 => \N__14454\,
            in2 => \N__13071\,
            in3 => \N__13063\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000101111111"
        )
    port map (
            in0 => \N__14347\,
            in1 => \N__14274\,
            in2 => \N__14181\,
            in3 => \N__14224\,
            lcout => \this_vga_signals.SUM_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13259\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_pcounter_q_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32623\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_RNIC95C3_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__13745\,
            in1 => \N__13728\,
            in2 => \_gnd_net_\,
            in3 => \N__21661\,
            lcout => \this_vga_signals.M_pcounter_q_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI3O9R_1_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14806\,
            in1 => \N__14618\,
            in2 => \_gnd_net_\,
            in3 => \N__14548\,
            lcout => \this_vga_signals.N_17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_1_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010011110000"
        )
    port map (
            in0 => \N__21662\,
            in1 => \N__13709\,
            in2 => \N__13734\,
            in3 => \N__21525\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32623\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI9JJM1_0_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__13241\,
            in1 => \N__14476\,
            in2 => \N__14853\,
            in3 => \N__14420\,
            lcout => \this_vga_signals.M_hcounter_q_RNI9JJM1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIADGD1_5_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__13242\,
            in1 => \N__14477\,
            in2 => \_gnd_net_\,
            in3 => \N__14421\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_hcounter_q_RNIADGD1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIOC7D3_6_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__14363\,
            in1 => \N__13233\,
            in2 => \N__13227\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.i5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000101"
        )
    port map (
            in0 => \N__14247\,
            in1 => \_gnd_net_\,
            in2 => \N__14196\,
            in3 => \N__14305\,
            lcout => this_vga_signals_hvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111010111"
        )
    port map (
            in0 => \N__14245\,
            in1 => \N__14191\,
            in2 => \N__14309\,
            in3 => \N__14364\,
            lcout => \this_vga_signals.SUM_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIML464_9_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__14192\,
            in1 => \N__13449\,
            in2 => \N__14310\,
            in3 => \N__14246\,
            lcout => this_vga_signals_hsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNI1DAA_7_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16158\,
            in2 => \_gnd_net_\,
            in3 => \N__16205\,
            lcout => \M_this_ppu_map_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI9E7F1_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24507\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19892\,
            lcout => \N_63_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIMF36L_9_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17079\,
            in1 => \N__13398\,
            in2 => \_gnd_net_\,
            in3 => \N__13368\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIHL0E5_9_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13329\,
            in2 => \_gnd_net_\,
            in3 => \N__17078\,
            lcout => \M_this_vga_signals_address_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_29_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24502\,
            lcout => \M_this_data_tmp_qZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32541\,
            ce => \N__17663\,
            sr => \N__26066\
        );

    \M_this_data_tmp_q_esr_5_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24490\,
            lcout => \M_this_data_tmp_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32550\,
            ce => \N__16520\,
            sr => \N__26063\
        );

    \M_this_data_tmp_q_esr_12_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28324\,
            lcout => \M_this_data_tmp_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32562\,
            ce => \N__17352\,
            sr => \N__26060\
        );

    \M_this_data_tmp_q_esr_13_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24489\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32562\,
            ce => \N__17352\,
            sr => \N__26060\
        );

    \M_this_data_tmp_q_esr_9_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30929\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32562\,
            ce => \N__17352\,
            sr => \N__26060\
        );

    \M_this_data_tmp_q_esr_0_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28447\,
            lcout => \M_this_data_tmp_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32571\,
            ce => \N__16512\,
            sr => \N__26056\
        );

    \this_ppu.M_haddress_q_5_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13558\,
            in2 => \_gnd_net_\,
            in3 => \N__13457\,
            lcout => \M_this_ppu_map_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32581\,
            ce => 'H',
            sr => \N__14922\
        );

    \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__28527\,
            in1 => \N__26991\,
            in2 => \N__28677\,
            in3 => \N__28626\,
            lcout => \M_this_ppu_vram_data_0\,
            ltout => \M_this_ppu_vram_data_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.vram_en_i_a2_0_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28783\,
            in1 => \N__17182\,
            in2 => \N__13467\,
            in3 => \N__21160\,
            lcout => \this_ppu.N_134\,
            ltout => \this_ppu.N_134_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIUTM1G_5_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14640\,
            in2 => \N__13464\,
            in3 => \N__32123\,
            lcout => \M_this_ppu_vram_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_6_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__13559\,
            in1 => \N__13606\,
            in2 => \_gnd_net_\,
            in3 => \N__13458\,
            lcout => \M_this_ppu_vram_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32581\,
            ce => 'H',
            sr => \N__14922\
        );

    \this_ppu.M_haddress_q_RNINDU1G_1_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20910\,
            in1 => \N__19285\,
            in2 => \_gnd_net_\,
            in3 => \N__13995\,
            lcout => \this_ppu.un1_M_haddress_q_c2\,
            ltout => \this_ppu.un1_M_haddress_q_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI4T92G_4_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13796\,
            in1 => \N__13927\,
            in2 => \N__13461\,
            in3 => \N__13873\,
            lcout => \this_ppu.un1_M_haddress_q_c5\,
            ltout => \this_ppu.un1_M_haddress_q_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_7_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__13607\,
            in1 => \N__13560\,
            in2 => \N__13530\,
            in3 => \N__13527\,
            lcout => \this_ppu.M_haddress_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32581\,
            ce => 'H',
            sr => \N__14922\
        );

    \this_ppu.M_state_q_1_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__32140\,
            in1 => \N__13977\,
            in2 => \N__14694\,
            in3 => \N__13758\,
            lcout => \this_ppu.M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32590\,
            ce => 'H',
            sr => \N__26051\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14849\,
            in2 => \N__14808\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_21_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21491\,
            in1 => \N__14617\,
            in2 => \_gnd_net_\,
            in3 => \N__13515\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__32598\,
            ce => 'H',
            sr => \N__14750\
        );

    \this_vga_signals.M_hcounter_q_3_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21488\,
            in1 => \N__14528\,
            in2 => \_gnd_net_\,
            in3 => \N__13512\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__32598\,
            ce => 'H',
            sr => \N__14750\
        );

    \this_vga_signals.M_hcounter_q_4_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21492\,
            in1 => \N__14474\,
            in2 => \_gnd_net_\,
            in3 => \N__13509\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__32598\,
            ce => 'H',
            sr => \N__14750\
        );

    \this_vga_signals.M_hcounter_q_5_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21489\,
            in1 => \N__14412\,
            in2 => \_gnd_net_\,
            in3 => \N__13506\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \N__32598\,
            ce => 'H',
            sr => \N__14750\
        );

    \this_vga_signals.M_hcounter_q_6_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21493\,
            in1 => \N__14359\,
            in2 => \_gnd_net_\,
            in3 => \N__13503\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \N__32598\,
            ce => 'H',
            sr => \N__14750\
        );

    \this_vga_signals.M_hcounter_q_7_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21490\,
            in1 => \N__14180\,
            in2 => \_gnd_net_\,
            in3 => \N__13500\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \N__32598\,
            ce => 'H',
            sr => \N__14750\
        );

    \this_vga_signals.M_hcounter_q_8_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21494\,
            in1 => \N__14235\,
            in2 => \_gnd_net_\,
            in3 => \N__13752\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \N__32598\,
            ce => 'H',
            sr => \N__14750\
        );

    \this_vga_signals.M_hcounter_q_esr_9_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14290\,
            in2 => \_gnd_net_\,
            in3 => \N__13749\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32607\,
            ce => \N__14862\,
            sr => \N__14749\
        );

    \this_vga_signals.M_pcounter_q_0_e_0_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__13746\,
            in1 => \N__13733\,
            in2 => \_gnd_net_\,
            in3 => \N__21638\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32617\,
            ce => \N__21524\,
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI7C7F1_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31330\,
            in2 => \_gnd_net_\,
            in3 => \N__19876\,
            lcout => \N_815_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIE00C4_9_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__14292\,
            in1 => \N__14236\,
            in2 => \N__15865\,
            in3 => \N__14182\,
            lcout => \M_this_vga_ramdac_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI8D7F1_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28245\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19823\,
            lcout => \N_814_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNI0655_6_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16206\,
            lcout => \this_ppu_M_vaddress_q_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_1_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30846\,
            lcout => \M_this_data_tmp_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32542\,
            ce => \N__16516\,
            sr => \N__26061\
        );

    \M_this_data_tmp_q_esr_24_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28454\,
            lcout => \M_this_data_tmp_qZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32551\,
            ce => \N__17649\,
            sr => \N__26057\
        );

    \M_this_data_tmp_q_esr_6_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28148\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32563\,
            ce => \N__16499\,
            sr => \N__26054\
        );

    \this_ppu.M_haddress_q_RNIEV7R_2_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__32134\,
            in1 => \N__13863\,
            in2 => \N__31935\,
            in3 => \N__14130\,
            lcout => \M_this_ppu_sprites_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_2_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__13997\,
            in1 => \N__13865\,
            in2 => \N__19307\,
            in3 => \N__20912\,
            lcout => \M_this_ppu_vram_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32572\,
            ce => 'H',
            sr => \N__14918\
        );

    \this_ppu.M_haddress_q_RNO_0_3_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__32133\,
            in1 => \N__19286\,
            in2 => \N__14649\,
            in3 => \N__13975\,
            lcout => OPEN,
            ltout => \this_ppu.un1_M_haddress_q_c1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_3_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__13928\,
            in1 => \N__13866\,
            in2 => \N__14013\,
            in3 => \N__20913\,
            lcout => \M_this_ppu_map_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32572\,
            ce => 'H',
            sr => \N__14918\
        );

    \this_ppu.M_haddress_q_1_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__20911\,
            in1 => \N__19290\,
            in2 => \_gnd_net_\,
            in3 => \N__13996\,
            lcout => \M_this_ppu_vram_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32572\,
            ce => 'H',
            sr => \N__14918\
        );

    \this_ppu.M_haddress_q_0_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010110100111100"
        )
    port map (
            in0 => \N__13976\,
            in1 => \N__14647\,
            in2 => \N__19306\,
            in3 => \N__32135\,
            lcout => \M_this_ppu_vram_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32572\,
            ce => 'H',
            sr => \N__14918\
        );

    \this_ppu.M_haddress_q_4_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__13929\,
            in1 => \N__13864\,
            in2 => \N__13797\,
            in3 => \N__13833\,
            lcout => \M_this_ppu_map_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32572\,
            ce => 'H',
            sr => \N__14918\
        );

    \this_ppu.M_state_q_RNO_1_1_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__16982\,
            in1 => \N__32132\,
            in2 => \N__14648\,
            in3 => \N__16917\,
            lcout => \this_ppu.N_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_1_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__14657\,
            in1 => \N__31883\,
            in2 => \_gnd_net_\,
            in3 => \N__17459\,
            lcout => \this_ppu.M_state_qc_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_4_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14672\,
            in2 => \_gnd_net_\,
            in3 => \N__28791\,
            lcout => OPEN,
            ltout => \this_ppu.M_state_qc_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_4_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32136\,
            in1 => \N__17189\,
            in2 => \N__14661\,
            in3 => \N__21161\,
            lcout => \this_ppu.M_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32582\,
            ce => 'H',
            sr => \N__26048\
        );

    \this_ppu.M_state_q_5_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14658\,
            lcout => \this_ppu.M_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32582\,
            ce => 'H',
            sr => \N__26048\
        );

    \this_start_data_delay.G_464_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21478\,
            in2 => \_gnd_net_\,
            in3 => \N__21637\,
            lcout => \G_464\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111111111111"
        )
    port map (
            in0 => \N__14772\,
            in1 => \N__14828\,
            in2 => \N__14611\,
            in3 => \N__14521\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_18_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIEVMV1_5_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__14472\,
            in1 => \N__14411\,
            in2 => \N__14367\,
            in3 => \N__14352\,
            lcout => OPEN,
            ltout => \this_vga_signals.m23_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000001000"
        )
    port map (
            in0 => \N__14278\,
            in1 => \N__14226\,
            in2 => \N__14199\,
            in3 => \N__14171\,
            lcout => \this_vga_signals_M_hcounter_d7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21521\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14742\,
            lcout => \this_vga_signals.N_1090_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_0_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21522\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14838\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32608\,
            ce => 'H',
            sr => \N__14751\
        );

    \this_vga_signals.M_hcounter_q_1_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__14837\,
            in1 => \N__21523\,
            in2 => \_gnd_net_\,
            in3 => \N__14783\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32608\,
            ce => 'H',
            sr => \N__14751\
        );

    \this_reset_cond.M_stage_q_1_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16303\,
            in2 => \_gnd_net_\,
            in3 => \N__14997\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16304\,
            in2 => \_gnd_net_\,
            in3 => \N__14721\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__16302\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14715\,
            lcout => \this_reset_cond.M_stage_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_0_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__15357\,
            in1 => \N__15171\,
            in2 => \_gnd_net_\,
            in3 => \N__15120\,
            lcout => \this_ppu.M_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_oam_ram_write_data_10_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15402\,
            in2 => \_gnd_net_\,
            in3 => \N__18527\,
            lcout => \M_this_oam_ram_write_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15356\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \this_ppu.un1_M_count_q_1_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14937\,
            in2 => \N__29676\,
            in3 => \N__14697\,
            lcout => \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_0_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29569\,
            in2 => \N__15330\,
            in3 => \N__14892\,
            lcout => \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_1_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15374\,
            in2 => \N__29677\,
            in3 => \N__14889\,
            lcout => \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_2_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29573\,
            in2 => \N__14955\,
            in3 => \N__14886\,
            lcout => \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_3_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14972\,
            in2 => \N__29678\,
            in3 => \N__14883\,
            lcout => \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_4_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29577\,
            in2 => \N__15087\,
            in3 => \N__14880\,
            lcout => \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_5_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_7_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110110"
        )
    port map (
            in0 => \N__17467\,
            in1 => \N__15434\,
            in2 => \N__16887\,
            in3 => \N__14877\,
            lcout => \this_ppu.M_count_q_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIKRC91_1_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17466\,
            in1 => \N__17420\,
            in2 => \_gnd_net_\,
            in3 => \N__17402\,
            lcout => \this_ppu.M_state_d_0_sqmuxa_1\,
            ltout => \this_ppu.M_state_d_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI2UC86_1_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15773\,
            in2 => \N__14874\,
            in3 => \N__16876\,
            lcout => \this_ppu.N_1456_0\,
            ltout => \this_ppu.N_1456_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_4_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000010000"
        )
    port map (
            in0 => \N__15161\,
            in1 => \N__14871\,
            in2 => \N__14865\,
            in3 => \N__14951\,
            lcout => \this_ppu.M_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_5_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000000010"
        )
    port map (
            in0 => \N__15116\,
            in1 => \N__14991\,
            in2 => \N__15172\,
            in3 => \N__14973\,
            lcout => \this_ppu.M_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_1_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100100000000"
        )
    port map (
            in0 => \N__14936\,
            in1 => \N__15160\,
            in2 => \N__14985\,
            in3 => \N__15115\,
            lcout => \this_ppu.M_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32564\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNICD0G_1_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14971\,
            in1 => \N__14950\,
            in2 => \N__15086\,
            in3 => \N__14935\,
            lcout => \this_ppu.M_state_q_srsts_i_a3_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIE20V4_0_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__16974\,
            in1 => \N__15772\,
            in2 => \N__16922\,
            in3 => \N__16944\,
            lcout => \this_ppu.M_state_q_RNIE20V4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNIAUKV3_0_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__15030\,
            in1 => \N__15051\,
            in2 => \_gnd_net_\,
            in3 => \N__15902\,
            lcout => \M_this_vga_signals_line_clk_0\,
            ltout => \M_this_vga_signals_line_clk_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI2TJN4_0_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__16972\,
            in1 => \_gnd_net_\,
            in2 => \N__14901\,
            in3 => \N__16943\,
            lcout => \this_ppu.M_state_d_0_sqmuxa\,
            ltout => \this_ppu.M_state_d_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIJV275_2_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30281\,
            in1 => \N__16833\,
            in2 => \N__14898\,
            in3 => \N__32177\,
            lcout => \this_ppu.un1_M_vaddress_q_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNO_0_0_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15031\,
            in2 => \_gnd_net_\,
            in3 => \N__15932\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_1000_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_0_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010011001100"
        )
    port map (
            in0 => \N__21660\,
            in1 => \N__15052\,
            in2 => \N__14895\,
            in3 => \N__21536\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32573\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI22015_0_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__16973\,
            in1 => \N__16945\,
            in2 => \N__17468\,
            in3 => \N__16916\,
            lcout => \this_ppu.un10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_4_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16280\,
            in2 => \_gnd_net_\,
            in3 => \N__15063\,
            lcout => \this_reset_cond.M_stage_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__15054\,
            in1 => \N__15032\,
            in2 => \_gnd_net_\,
            in3 => \N__15903\,
            lcout => \this_ppu.M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIE6DH5_4_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16625\,
            in1 => \N__16691\,
            in2 => \_gnd_net_\,
            in3 => \N__16712\,
            lcout => \this_ppu.un1_M_vaddress_q_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNO_0_1_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15053\,
            in2 => \_gnd_net_\,
            in3 => \N__15933\,
            lcout => OPEN,
            ltout => \this_vga_signals.i21_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_1_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110001011101010"
        )
    port map (
            in0 => \N__15033\,
            in1 => \N__21495\,
            in2 => \N__15036\,
            in3 => \N__21639\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32583\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIGB2A6_6_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__21622\,
            in1 => \N__15408\,
            in2 => \_gnd_net_\,
            in3 => \N__22400\,
            lcout => \this_vga_signals.N_129_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_6_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__16197\,
            in1 => \N__16775\,
            in2 => \_gnd_net_\,
            in3 => \N__16175\,
            lcout => \this_ppu.M_vaddress_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32609\,
            ce => 'H',
            sr => \N__16584\
        );

    \this_start_data_delay.M_last_q_RNI5A7F1_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30863\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19872\,
            lcout => \N_817_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16293\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_10_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32826\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32535\,
            ce => \N__17339\,
            sr => \N__26055\
        );

    \M_this_data_tmp_q_esr_17_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30913\,
            lcout => \M_this_data_tmp_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32538\,
            ce => \N__15947\,
            sr => \N__26052\
        );

    \this_ppu.M_count_q_3_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100100000000"
        )
    port map (
            in0 => \N__15375\,
            in1 => \N__15174\,
            in2 => \N__15384\,
            in3 => \N__15119\,
            lcout => \this_ppu.M_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNI890G_7_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15373\,
            in1 => \N__15325\,
            in2 => \N__15435\,
            in3 => \N__15355\,
            lcout => \this_ppu.M_state_q_srsts_i_a3_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_2_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100100000000"
        )
    port map (
            in0 => \N__15326\,
            in1 => \N__15173\,
            in2 => \N__15339\,
            in3 => \N__15118\,
            lcout => \this_ppu.M_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIMGCA_0_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16820\,
            in2 => \_gnd_net_\,
            in3 => \N__16449\,
            lcout => OPEN,
            ltout => \this_ppu.un10_sprites_addr_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIMQ241_2_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101001110"
        )
    port map (
            in0 => \N__31884\,
            in1 => \N__15312\,
            in2 => \N__15294\,
            in3 => \N__32076\,
            lcout => \M_this_ppu_sprites_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_6_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100100000000"
        )
    port map (
            in0 => \N__15085\,
            in1 => \N__15165\,
            in2 => \N__15132\,
            in3 => \N__15117\,
            lcout => \this_ppu.M_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIS8A01_0_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__16821\,
            in1 => \N__32078\,
            in2 => \N__31912\,
            in3 => \N__15726\,
            lcout => \M_this_ppu_sprites_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_0_RNISG75_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15606\,
            lcout => \M_this_oam_ram_read_data_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIMTR41_2_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32077\,
            in1 => \N__31885\,
            in2 => \N__15591\,
            in3 => \N__16416\,
            lcout => \M_this_ppu_sprites_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.dmalto4_0_o2_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110100010"
        )
    port map (
            in0 => \N__17775\,
            in1 => \N__19046\,
            in2 => \N__24318\,
            in3 => \N__22178\,
            lcout => \this_start_data_delay.N_43_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIELANC_0_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110101010"
        )
    port map (
            in0 => \N__15771\,
            in1 => \N__15850\,
            in2 => \N__17724\,
            in3 => \N__16871\,
            lcout => \this_ppu.M_state_q_RNIELANCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_0_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111100011111100"
        )
    port map (
            in0 => \N__16978\,
            in1 => \N__16946\,
            in2 => \N__15456\,
            in3 => \N__16921\,
            lcout => \this_ppu.M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32565\,
            ce => 'H',
            sr => \N__26045\
        );

    \this_ppu.M_count_q_7_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__15452\,
            in1 => \N__15444\,
            in2 => \_gnd_net_\,
            in3 => \N__16872\,
            lcout => \this_ppu.M_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32565\,
            ce => 'H',
            sr => \N__26045\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI4KCU6_9_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__22580\,
            in1 => \_gnd_net_\,
            in2 => \N__15417\,
            in3 => \N__21476\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNI4KCU6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI8O063_8_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21990\,
            in1 => \N__23091\,
            in2 => \N__15918\,
            in3 => \N__21893\,
            lcout => \this_vga_signals.N_1028\,
            ltout => \this_vga_signals.N_1028_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIFPFL6_9_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011001100"
        )
    port map (
            in0 => \N__22403\,
            in1 => \N__21670\,
            in2 => \N__15936\,
            in3 => \N__22581\,
            lcout => \this_vga_signals.N_999\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22929\,
            in2 => \_gnd_net_\,
            in3 => \N__21579\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_1004_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIILO32_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__22859\,
            in1 => \N__22704\,
            in2 => \N__15921\,
            in3 => \N__20518\,
            lcout => \this_vga_signals.N_1013\,
            ltout => \this_vga_signals.N_1013_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI9AJQ2_5_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010001"
        )
    port map (
            in0 => \N__22401\,
            in1 => \N__23090\,
            in2 => \N__15909\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_105_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI3HRS3_8_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100111"
        )
    port map (
            in0 => \N__21892\,
            in1 => \N__21989\,
            in2 => \N__15906\,
            in3 => \N__22579\,
            lcout => \this_vga_signals.N_113_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_6_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16317\,
            in2 => \_gnd_net_\,
            in3 => \N__15885\,
            lcout => \this_reset_cond.M_stage_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_5_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__16316\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15891\,
            lcout => \this_reset_cond.M_stage_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIGN2J3_9_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__17025\,
            in1 => \N__20255\,
            in2 => \N__16215\,
            in3 => \N__22584\,
            lcout => this_vga_signals_vvisibility,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_9_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__16320\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16221\,
            lcout => \M_this_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_7_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16318\,
            in2 => \_gnd_net_\,
            in3 => \N__16326\,
            lcout => \this_reset_cond.M_stage_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_8_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__16319\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16227\,
            lcout => \this_reset_cond.M_stage_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_8_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21902\,
            in1 => \N__22000\,
            in2 => \N__22402\,
            in3 => \N__22583\,
            lcout => \this_vga_signals.vaddress_ac0_9_0_a0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_7_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__16198\,
            in1 => \N__16771\,
            in2 => \N__16157\,
            in3 => \N__16176\,
            lcout => \this_ppu.M_vaddress_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32599\,
            ce => 'H',
            sr => \N__16583\
        );

    \this_ppu.M_state_q_3_LC_15_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31965\,
            lcout => \this_ppu.M_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32640\,
            ce => 'H',
            sr => \N__26044\
        );

    \M_this_state_q_17_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19404\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24243\,
            lcout => led23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32530\,
            ce => 'H',
            sr => \N__26053\
        );

    \dma_0_sbtinv_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17734\,
            lcout => dma_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI8G791_14_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__26204\,
            in1 => \N__19119\,
            in2 => \_gnd_net_\,
            in3 => \N__24235\,
            lcout => \N_1430_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.port_data_rw_0_a2_1_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__31649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23913\,
            lcout => \this_start_data_delay.port_data_rw_0_a2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIUCR11_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19403\,
            in2 => \_gnd_net_\,
            in3 => \N__24242\,
            lcout => OPEN,
            ltout => \M_this_state_q_ns_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_RNIAI791_9_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16524\,
            in3 => \N__26203\,
            lcout => \M_this_state_q_ns_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_12_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31856\,
            in1 => \N__32142\,
            in2 => \N__16470\,
            in3 => \N__16353\,
            lcout => \this_sprites_ram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un10_sprites_addr_cry_0_c_inv_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16428\,
            in2 => \N__16832\,
            in3 => \N__16448\,
            lcout => \this_ppu.M_this_oam_ram_read_data_iZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \this_ppu.un10_sprites_addr_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un10_sprites_addr_cry_0_c_RNIMJ5B_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16422\,
            in2 => \N__32176\,
            in3 => \N__16410\,
            lcout => \this_ppu.un10_sprites_addr_cry_0_c_RNIMJ5BZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un10_sprites_addr_cry_0\,
            carryout => \this_ppu.un10_sprites_addr_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un10_sprites_addr_cry_1_c_RNIOM6B_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16407\,
            in2 => \N__30280\,
            in3 => \N__16392\,
            lcout => \this_ppu.un10_sprites_addr_cry_1_c_RNIOM6BZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un10_sprites_addr_cry_1\,
            carryout => \this_ppu.un10_sprites_addr_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un10_sprites_addr_cry_2_c_RNIQP7B_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16389\,
            in2 => \N__16682\,
            in3 => \N__16374\,
            lcout => \this_ppu.un10_sprites_addr_cry_2_c_RNIQP7BZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un10_sprites_addr_cry_2\,
            carryout => \this_ppu.un10_sprites_addr_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un10_sprites_addr_cry_3_c_RNISS8B_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16610\,
            in2 => \N__16371\,
            in3 => \N__16347\,
            lcout => \this_ppu.un10_sprites_addr_cry_3_c_RNISS8BZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un10_sprites_addr_cry_3\,
            carryout => \this_ppu.un10_sprites_addr_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un10_sprites_addr_cry_4_c_RNIUV9B_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__16751\,
            in1 => \N__16344\,
            in2 => \_gnd_net_\,
            in3 => \N__16329\,
            lcout => \this_ppu.un10_sprites_addr_cry_4_c_RNIUV9BZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_0_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__16986\,
            in1 => \N__16947\,
            in2 => \N__16834\,
            in3 => \N__16923\,
            lcout => \M_this_ppu_vram_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32548\,
            ce => 'H',
            sr => \N__16582\
        );

    \this_ppu.M_vaddress_q_1_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__32174\,
            in1 => \N__16825\,
            in2 => \_gnd_net_\,
            in3 => \N__16886\,
            lcout => \this_ppu.M_vaddress_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32548\,
            ce => 'H',
            sr => \N__16582\
        );

    \this_ppu.M_vaddress_q_2_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__16885\,
            in1 => \N__32175\,
            in2 => \N__16835\,
            in3 => \N__30279\,
            lcout => \this_ppu.M_vaddress_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32548\,
            ce => 'H',
            sr => \N__16582\
        );

    \this_ppu.M_vaddress_q_5_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__16722\,
            in1 => \N__16755\,
            in2 => \N__16687\,
            in3 => \N__16615\,
            lcout => \M_this_ppu_map_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32548\,
            ce => 'H',
            sr => \N__16582\
        );

    \this_ppu.M_vaddress_q_3_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16672\,
            in2 => \_gnd_net_\,
            in3 => \N__16720\,
            lcout => \M_this_ppu_map_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32548\,
            ce => 'H',
            sr => \N__16582\
        );

    \this_ppu.M_vaddress_q_4_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__16721\,
            in1 => \_gnd_net_\,
            in2 => \N__16686\,
            in3 => \N__16614\,
            lcout => \M_this_ppu_map_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32548\,
            ce => 'H',
            sr => \N__16582\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIPE977_9_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21477\,
            in2 => \_gnd_net_\,
            in3 => \N__16541\,
            lcout => \this_vga_signals.N_1090_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101110010"
        )
    port map (
            in0 => \N__17019\,
            in1 => \N__17673\,
            in2 => \N__17580\,
            in3 => \N__17562\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__17373\,
            in1 => \N__22935\,
            in2 => \N__16527\,
            in3 => \N__17007\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_c3_0_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI3KH3P1_1_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__17130\,
            in1 => \N__17385\,
            in2 => \N__17049\,
            in3 => \N__17523\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICM2P1_5_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__23087\,
            in1 => \N__23248\,
            in2 => \N__22437\,
            in3 => \N__22386\,
            lcout => \this_vga_signals.un6_vvisibilitylt9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__16992\,
            in1 => \N__17967\,
            in2 => \N__18057\,
            in3 => \N__17571\,
            lcout => \this_vga_signals.g2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_8_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011100111"
        )
    port map (
            in0 => \N__21903\,
            in1 => \N__22001\,
            in2 => \N__20187\,
            in3 => \N__22582\,
            lcout => OPEN,
            ltout => \this_vga_signals.SUM_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_13_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010100101"
        )
    port map (
            in0 => \N__22002\,
            in1 => \N__22391\,
            in2 => \N__17013\,
            in3 => \N__20256\,
            lcout => \this_vga_signals.g3_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_2_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__22861\,
            in1 => \N__20286\,
            in2 => \N__23286\,
            in3 => \N__18260\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c2_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_8_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18261\,
            in1 => \N__18702\,
            in2 => \N__17010\,
            in3 => \N__17586\,
            lcout => \this_vga_signals.N_4_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_a3_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111101"
        )
    port map (
            in0 => \N__23278\,
            in1 => \N__22392\,
            in2 => \N__23100\,
            in3 => \N__20424\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g4_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011111100"
        )
    port map (
            in0 => \N__22393\,
            in1 => \N__17001\,
            in2 => \N__16995\,
            in3 => \N__18885\,
            lcout => \this_vga_signals.g4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI9H791_15_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__26205\,
            in1 => \N__19146\,
            in2 => \_gnd_net_\,
            in3 => \N__24241\,
            lcout => \N_1438_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.port_data_rw_0_i_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__23576\,
            in1 => \N__17304\,
            in2 => \N__18153\,
            in3 => \N__17766\,
            lcout => port_data_rw_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17274\,
            in1 => \N__17262\,
            in2 => \_gnd_net_\,
            in3 => \N__30108\,
            lcout => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_3_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17250\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30100\,
            in1 => \N__17232\,
            in2 => \_gnd_net_\,
            in3 => \N__17217\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__28719\,
            in1 => \N__28661\,
            in2 => \N__17202\,
            in3 => \N__28587\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__28662\,
            in1 => \N__17199\,
            in2 => \N__17193\,
            in3 => \N__17475\,
            lcout => \M_this_ppu_vram_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_11_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__17157\,
            in1 => \N__17151\,
            in2 => \N__31882\,
            in3 => \N__32124\,
            lcout => \this_sprites_ram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30101\,
            in1 => \N__17505\,
            in2 => \_gnd_net_\,
            in3 => \N__17490\,
            lcout => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_2_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__17469\,
            in1 => \N__17427\,
            in2 => \_gnd_net_\,
            in3 => \N__17409\,
            lcout => \this_ppu.M_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32566\,
            ce => 'H',
            sr => \N__26046\
        );

    \m1_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__17886\,
            in1 => \N__17929\,
            in2 => \_gnd_net_\,
            in3 => \N__18078\,
            lcout => OPEN,
            ltout => \N_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIRPN94A_2_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101100100100"
        )
    port map (
            in0 => \N__22840\,
            in1 => \N__22715\,
            in2 => \N__17391\,
            in3 => \N__17514\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI75QSCH1_2_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101101000111"
        )
    port map (
            in0 => \N__17367\,
            in1 => \N__17826\,
            in2 => \N__17388\,
            in3 => \N__17379\,
            lcout => \this_vga_signals.vaddress_N_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010001001011"
        )
    port map (
            in0 => \N__18080\,
            in1 => \N__17885\,
            in2 => \N__18009\,
            in3 => \N__17838\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_11_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17871\,
            in1 => \N__17547\,
            in2 => \N__17910\,
            in3 => \N__18007\,
            lcout => \this_vga_signals.mult1_un75_sum_axb1_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIDON0D8_3_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011011000011"
        )
    port map (
            in0 => \N__18079\,
            in1 => \N__22839\,
            in2 => \N__17934\,
            in3 => \N__17884\,
            lcout => \this_vga_signals.N_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_m2_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000001111"
        )
    port map (
            in0 => \N__22714\,
            in1 => \N__18324\,
            in2 => \N__22865\,
            in3 => \N__17597\,
            lcout => \this_vga_signals.mult1_un68_sum_c3\,
            ltout => \this_vga_signals.mult1_un68_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIKLMK17_2_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18027\,
            in1 => \N__17953\,
            in2 => \N__17553\,
            in3 => \N__17820\,
            lcout => \this_vga_signals.g0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_0_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001011001"
        )
    port map (
            in0 => \N__18297\,
            in1 => \N__18099\,
            in2 => \N__23277\,
            in3 => \N__19008\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__18230\,
            in1 => \_gnd_net_\,
            in2 => \N__17550\,
            in3 => \N__18767\,
            lcout => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100101011"
        )
    port map (
            in0 => \N__18766\,
            in1 => \N__23266\,
            in2 => \N__22868\,
            in3 => \N__18231\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m2_3_1_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18232\,
            in1 => \N__17546\,
            in2 => \N__17958\,
            in3 => \N__17928\,
            lcout => \this_vga_signals.if_m2_3_1\,
            ltout => \this_vga_signals.if_m2_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIBALLEF_2_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010001000001"
        )
    port map (
            in0 => \N__22706\,
            in1 => \N__18033\,
            in2 => \N__17535\,
            in3 => \N__18008\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIOP5EV51_1_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101111110100"
        )
    port map (
            in0 => \N__17985\,
            in1 => \N__22934\,
            in2 => \N__17532\,
            in3 => \N__17529\,
            lcout => \this_vga_signals.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m1_0_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18768\,
            in1 => \N__23267\,
            in2 => \_gnd_net_\,
            in3 => \N__18229\,
            lcout => \this_vga_signals.if_m1_0\,
            ltout => \this_vga_signals.if_m1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m1_9_0_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001110111100"
        )
    port map (
            in0 => \N__18323\,
            in1 => \N__22854\,
            in2 => \N__17517\,
            in3 => \N__22705\,
            lcout => \this_vga_signals.if_m1_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIVGRQM1_1_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__18249\,
            in1 => \N__22933\,
            in2 => \_gnd_net_\,
            in3 => \N__18120\,
            lcout => \this_vga_signals.N_129_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23259\,
            in2 => \_gnd_net_\,
            in3 => \N__18762\,
            lcout => \this_vga_signals.if_m1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000001111"
        )
    port map (
            in0 => \N__22707\,
            in1 => \N__18316\,
            in2 => \N__22869\,
            in3 => \N__17598\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_0_a3_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18114\,
            in1 => \N__18763\,
            in2 => \N__18108\,
            in3 => \N__18251\,
            lcout => \this_vga_signals.g0_3_0_a3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100101011"
        )
    port map (
            in0 => \N__18250\,
            in1 => \N__22857\,
            in2 => \N__23282\,
            in3 => \N__18781\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111111111001"
        )
    port map (
            in0 => \N__18782\,
            in1 => \N__18247\,
            in2 => \N__23099\,
            in3 => \N__20667\,
            lcout => \this_vga_signals.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_1_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100101011"
        )
    port map (
            in0 => \N__18248\,
            in1 => \N__22856\,
            in2 => \N__23283\,
            in3 => \N__18783\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c2_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_10_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22361\,
            in1 => \N__18126\,
            in2 => \N__17565\,
            in3 => \N__18138\,
            lcout => \this_vga_signals.g0_i_x4_7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_9_N_2L1_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23284\,
            in3 => \N__18772\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_9_N_2L1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_9_N_3L3_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100010000101"
        )
    port map (
            in0 => \N__22866\,
            in1 => \N__18636\,
            in2 => \N__17556\,
            in3 => \N__18242\,
            lcout => \this_vga_signals.g0_9_N_3L3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_1_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18924\,
            in1 => \N__18270\,
            in2 => \_gnd_net_\,
            in3 => \N__20372\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_i_x4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_3_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101110001"
        )
    port map (
            in0 => \N__22867\,
            in1 => \N__23272\,
            in2 => \N__17685\,
            in3 => \N__18243\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c2_0_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_9_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010001000001"
        )
    port map (
            in0 => \N__22708\,
            in1 => \N__18168\,
            in2 => \N__17682\,
            in3 => \N__17679\,
            lcout => \this_vga_signals.g0_i_a4_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_a0_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20580\,
            in2 => \_gnd_net_\,
            in3 => \N__20520\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_a1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI7F791_13_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__26206\,
            in1 => \N__19092\,
            in2 => \_gnd_net_\,
            in3 => \N__24227\,
            lcout => \N_1422_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_3_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__28965\,
            in1 => \N__29212\,
            in2 => \_gnd_net_\,
            in3 => \N__28979\,
            lcout => \M_this_data_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32546\,
            ce => \N__29108\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_14_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__29295\,
            in1 => \N__26963\,
            in2 => \N__28167\,
            in3 => \N__29188\,
            lcout => \M_this_data_count_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32554\,
            ce => \N__29103\,
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIICAO1_0_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__19628\,
            in1 => \N__18673\,
            in2 => \N__19705\,
            in3 => \N__18684\,
            lcout => \M_this_state_d_0_sqmuxa_2\,
            ltout => \M_this_state_d_0_sqmuxa_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_substate_q_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__18674\,
            in1 => \_gnd_net_\,
            in2 => \N__17601\,
            in3 => \N__18690\,
            lcout => \M_this_substate_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32567\,
            ce => 'H',
            sr => \N__26049\
        );

    \this_start_data_delay.M_last_q_RNILCRA6_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111001011111"
        )
    port map (
            in0 => \N__26967\,
            in1 => \N__26196\,
            in2 => \N__24462\,
            in3 => \N__24624\,
            lcout => \M_this_data_count_q_3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIK0EI1_3_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__19704\,
            in1 => \N__19627\,
            in2 => \N__19569\,
            in3 => \N__19490\,
            lcout => \this_start_data_delay.N_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.dmalto4_0_a2_0_1_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21262\,
            in2 => \_gnd_net_\,
            in3 => \N__23780\,
            lcout => \this_start_data_delay.N_76_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_1_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010100"
        )
    port map (
            in0 => \N__26207\,
            in1 => \N__21319\,
            in2 => \N__17787\,
            in3 => \N__24224\,
            lcout => \M_this_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIK0EI1_2_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__19703\,
            in1 => \N__19626\,
            in2 => \N__19568\,
            in3 => \N__19491\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_65_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_4_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110100"
        )
    port map (
            in0 => \N__24225\,
            in1 => \N__21263\,
            in2 => \N__17778\,
            in3 => \N__26208\,
            lcout => \M_this_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.dmalto4_0_o2_0_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011100000"
        )
    port map (
            in0 => \N__23781\,
            in1 => \N__21100\,
            in2 => \N__24313\,
            in3 => \N__21318\,
            lcout => \this_start_data_delay.N_42_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.dmalto4_0_a2_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__17762\,
            in1 => \N__23571\,
            in2 => \N__18399\,
            in3 => \N__19431\,
            lcout => dma_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_2_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22270\,
            in1 => \N__20245\,
            in2 => \N__20373\,
            in3 => \N__18884\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2\,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000110"
        )
    port map (
            in0 => \N__20371\,
            in1 => \N__22272\,
            in2 => \N__17688\,
            in3 => \N__17799\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000001110000"
        )
    port map (
            in0 => \N__18797\,
            in1 => \N__18785\,
            in2 => \N__17889\,
            in3 => \N__18257\,
            lcout => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3,
            ltout => \this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17874\,
            in3 => \N__18081\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un61_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m4_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__17865\,
            in1 => \N__17847\,
            in2 => \N__17841\,
            in3 => \N__17837\,
            lcout => \this_vga_signals.if_i4_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIKL00E1_2_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18258\,
            in1 => \N__22858\,
            in2 => \_gnd_net_\,
            in3 => \N__22713\,
            lcout => \this_vga_signals.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_1_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110101011"
        )
    port map (
            in0 => \N__22269\,
            in1 => \N__18883\,
            in2 => \N__17814\,
            in3 => \N__20423\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_0_2_1\,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_0_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_0_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20370\,
            in2 => \N__17793\,
            in3 => \N__22271\,
            lcout => \this_vga_signals.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__20660\,
            in1 => \N__23000\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc1\,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_0_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17790\,
            in3 => \N__18764\,
            lcout => \this_vga_signals.mult1_un61_sum_axb2_0\,
            ltout => \this_vga_signals.mult1_un61_sum_axb2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000100000"
        )
    port map (
            in0 => \N__22849\,
            in1 => \N__18233\,
            in2 => \N__18084\,
            in3 => \N__17975\,
            lcout => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d,
            ltout => \this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__18063\,
            in1 => \N__18047\,
            in2 => \N__18036\,
            in3 => \N__18132\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0_0\,
            ltout => \this_vga_signals.mult1_un61_sum_c3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17906\,
            in1 => \N__18026\,
            in2 => \N__18012\,
            in3 => \N__18003\,
            lcout => \this_vga_signals.mult1_un75_sum_axb1_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_19_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20661\,
            in2 => \N__23039\,
            in3 => \N__18765\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_4_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_12_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000010"
        )
    port map (
            in0 => \N__22850\,
            in1 => \N__18234\,
            in2 => \N__17979\,
            in3 => \N__17976\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_d_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_1_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18235\,
            in1 => \N__17957\,
            in2 => \N__22716\,
            in3 => \N__17933\,
            lcout => \this_vga_signals.mult1_un75_sum_axb1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_ns_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19023\,
            in1 => \N__20366\,
            in2 => \_gnd_net_\,
            in3 => \N__18930\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000001"
        )
    port map (
            in0 => \N__19014\,
            in1 => \N__19000\,
            in2 => \N__17895\,
            in3 => \N__18292\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_28_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23202\,
            in2 => \N__17892\,
            in3 => \N__18777\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_4_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_25_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101001111010"
        )
    port map (
            in0 => \N__22855\,
            in1 => \N__22702\,
            in2 => \N__18141\,
            in3 => \N__20610\,
            lcout => \this_vga_signals.N_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111001111101"
        )
    port map (
            in0 => \N__18776\,
            in1 => \N__20589\,
            in2 => \N__23092\,
            in3 => \N__18236\,
            lcout => \this_vga_signals.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_10_1_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__20656\,
            in1 => \N__23069\,
            in2 => \_gnd_net_\,
            in3 => \N__20691\,
            lcout => \this_vga_signals.g0_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20297\,
            in2 => \_gnd_net_\,
            in3 => \N__20655\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_0_8_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100101001101"
        )
    port map (
            in0 => \N__22578\,
            in1 => \N__21901\,
            in2 => \N__20183\,
            in3 => \N__21985\,
            lcout => \this_vga_signals.SUM_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNISDV89_4_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110110000111"
        )
    port map (
            in0 => \N__18984\,
            in1 => \N__18162\,
            in2 => \N__23203\,
            in3 => \N__20151\,
            lcout => \this_vga_signals.N_24_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_2_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100011010"
        )
    port map (
            in0 => \N__23268\,
            in1 => \N__18098\,
            in2 => \N__23097\,
            in3 => \N__20654\,
            lcout => \this_vga_signals.g1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_0_a3_3_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20653\,
            in1 => \N__18828\,
            in2 => \N__20274\,
            in3 => \N__22387\,
            lcout => \this_vga_signals.g0_3_0_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23077\,
            in1 => \N__23158\,
            in2 => \_gnd_net_\,
            in3 => \N__20652\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1\,
            ltout => \this_vga_signals.mult1_un54_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_x4_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110011010011"
        )
    port map (
            in0 => \N__23159\,
            in1 => \N__19004\,
            in2 => \N__18327\,
            in3 => \N__18293\,
            lcout => \this_vga_signals.if_N_9_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__18978\,
            in1 => \_gnd_net_\,
            in2 => \N__18882\,
            in3 => \N__20651\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_m2_LC_18_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111100001001"
        )
    port map (
            in0 => \N__18660\,
            in1 => \N__18276\,
            in2 => \N__18909\,
            in3 => \N__18920\,
            lcout => \this_vga_signals.mult1_un47_sum_c3_1_0\,
            ltout => \this_vga_signals.mult1_un47_sum_c3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_4_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18897\,
            in1 => \N__18784\,
            in2 => \N__18264\,
            in3 => \N__18259\,
            lcout => \this_vga_signals.g2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_7_LC_18_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001111101100"
        )
    port map (
            in0 => \N__23183\,
            in1 => \N__22362\,
            in2 => \N__23098\,
            in3 => \N__21999\,
            lcout => \this_vga_signals.m12_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_16_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__19394\,
            in1 => \N__19144\,
            in2 => \N__26226\,
            in3 => \N__24231\,
            lcout => \M_this_state_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32547\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_14_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__19115\,
            in1 => \N__19091\,
            in2 => \N__26225\,
            in3 => \N__24239\,
            lcout => \M_this_state_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un25_i_a2_3_a2_2_a3_3_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__23489\,
            in1 => \N__19764\,
            in2 => \N__20741\,
            in3 => \N__19427\,
            lcout => \this_start_data_delay.N_400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_12_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__18387\,
            in1 => \N__26214\,
            in2 => \N__26786\,
            in3 => \N__18483\,
            lcout => \M_this_state_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32555\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un25_i_a2_i_o2_4_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18482\,
            in2 => \_gnd_net_\,
            in3 => \N__19395\,
            lcout => \this_start_data_delay.N_55_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_ns_0_i_o2_0_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22167\,
            in1 => \N__21093\,
            in2 => \N__24317\,
            in3 => \N__21320\,
            lcout => \this_start_data_delay.N_112_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.dmalto4_0_a2_1_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23906\,
            in1 => \N__19755\,
            in2 => \N__23496\,
            in3 => \N__20730\,
            lcout => \this_start_data_delay.dmalto4_0_a2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_data_count_qlde_i_o2_1_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__20729\,
            in1 => \N__19754\,
            in2 => \_gnd_net_\,
            in3 => \N__23905\,
            lcout => \this_start_data_delay.N_90_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNICA9G3_0_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20731\,
            in2 => \_gnd_net_\,
            in3 => \N__23663\,
            lcout => \this_start_data_delay.N_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_3_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010100"
        )
    port map (
            in0 => \N__26211\,
            in1 => \N__22171\,
            in2 => \N__18381\,
            in3 => \N__24240\,
            lcout => \M_this_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI3MH61_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__18372\,
            in1 => \N__31596\,
            in2 => \N__18354\,
            in3 => \N__23733\,
            lcout => \this_start_data_delay.N_47_0\,
            ltout => \this_start_data_delay.N_47_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIVMHD1_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18333\,
            in3 => \N__19932\,
            lcout => \this_start_data_delay.N_48_0\,
            ltout => \this_start_data_delay.N_48_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIK0EI1_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001100000"
        )
    port map (
            in0 => \N__19687\,
            in1 => \N__19550\,
            in2 => \N__18330\,
            in3 => \N__19620\,
            lcout => \N_28_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI7R5F1_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__19933\,
            in1 => \N__19549\,
            in2 => \_gnd_net_\,
            in3 => \N__19967\,
            lcout => \this_start_data_delay.N_82\,
            ltout => \this_start_data_delay.N_82_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIICAO1_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__19619\,
            in1 => \N__19686\,
            in2 => \N__18678\,
            in3 => \N__18675\,
            lcout => \this_start_data_delay.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_x4_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000010011"
        )
    port map (
            in0 => \N__20504\,
            in1 => \N__22265\,
            in2 => \N__20579\,
            in3 => \N__21951\,
            lcout => \this_vga_signals.g0_0_x4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_6_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21715\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32585\,
            ce => \N__23407\,
            sr => \N__23313\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_0_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20130\,
            in3 => \N__20028\,
            lcout => \this_vga_signals.vaddress_c2\,
            ltout => \this_vga_signals.vaddress_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_24_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21949\,
            in1 => \N__20084\,
            in2 => \N__18648\,
            in3 => \N__22570\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_5_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_1_LC_19_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001011"
        )
    port map (
            in0 => \N__22571\,
            in1 => \N__21897\,
            in2 => \N__18645\,
            in3 => \N__21950\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_1_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__18804\,
            in1 => \N__19992\,
            in2 => \N__18642\,
            in3 => \N__19986\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_21_LC_19_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010110100"
        )
    port map (
            in0 => \N__23221\,
            in1 => \N__23065\,
            in2 => \N__18639\,
            in3 => \N__20666\,
            lcout => \this_vga_signals.N_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_0_LC_19_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__22264\,
            in1 => \N__20572\,
            in2 => \_gnd_net_\,
            in3 => \N__20503\,
            lcout => \this_vga_signals.g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_0_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__22703\,
            in1 => \N__18798\,
            in2 => \N__22860\,
            in3 => \N__18786\,
            lcout => \this_vga_signals.g0_5_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21385\,
            lcout => \this_vga_signals.M_vcounter_q_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32591\,
            ce => \N__23360\,
            sr => \N__23315\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__20552\,
            in1 => \N__20502\,
            in2 => \_gnd_net_\,
            in3 => \N__20073\,
            lcout => \this_vga_signals.vaddress_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21720\,
            lcout => \this_vga_signals.M_vcounter_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32591\,
            ce => \N__23360\,
            sr => \N__23315\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_a4_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21775\,
            in1 => \N__20072\,
            in2 => \N__20247\,
            in3 => \N__22545\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_0_a4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_1_LC_19_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111011"
        )
    port map (
            in0 => \N__22544\,
            in1 => \N__21819\,
            in2 => \N__20086\,
            in3 => \N__20233\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_19_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22994\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23201\,
            lcout => \this_vga_signals.vaddress_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_5_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21353\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32600\,
            ce => \N__23397\,
            sr => \N__23318\
        );

    \this_vga_signals.un5_vaddress_g2_1_0_LC_19_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22995\,
            in1 => \N__22843\,
            in2 => \_gnd_net_\,
            in3 => \N__22672\,
            lcout => \this_vga_signals.g2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_5_LC_19_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21354\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32600\,
            ce => \N__23397\,
            sr => \N__23318\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_ns_LC_19_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20126\,
            in2 => \N__20007\,
            in3 => \N__20262\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_602_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21352\,
            lcout => \this_vga_signals.M_vcounter_q_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32600\,
            ce => \N__23397\,
            sr => \N__23318\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_2_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__18839\,
            in1 => \N__21735\,
            in2 => \N__18855\,
            in3 => \N__18818\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_16_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__18819\,
            in1 => \N__18854\,
            in2 => \N__22020\,
            in3 => \N__18840\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_2_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110000110110"
        )
    port map (
            in0 => \N__18953\,
            in1 => \N__20334\,
            in2 => \N__20456\,
            in3 => \N__20414\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_3_ns_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20697\,
            in2 => \_gnd_net_\,
            in3 => \N__20246\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_19_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__20100\,
            in1 => \N__21734\,
            in2 => \N__18822\,
            in3 => \N__18817\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_x1_LC_19_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111010000000"
        )
    port map (
            in0 => \N__20450\,
            in1 => \N__18952\,
            in2 => \N__18807\,
            in3 => \N__18977\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_4_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_19_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000111011001"
        )
    port map (
            in0 => \N__18951\,
            in1 => \N__20333\,
            in2 => \N__20455\,
            in3 => \N__20413\,
            lcout => \this_vga_signals.mult1_un47_sum_c3\,
            ltout => \this_vga_signals.mult1_un47_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_19_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__20514\,
            in1 => \_gnd_net_\,
            in2 => \N__19017\,
            in3 => \N__20565\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_LC_19_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000110"
        )
    port map (
            in0 => \N__20351\,
            in1 => \N__18962\,
            in2 => \N__20457\,
            in3 => \N__20410\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI6FO86_LC_19_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110100000"
        )
    port map (
            in0 => \N__20412\,
            in1 => \_gnd_net_\,
            in2 => \N__18966\,
            in3 => \N__20454\,
            lcout => \this_vga_signals.i1_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_0_LC_19_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111101110"
        )
    port map (
            in0 => \N__20509\,
            in1 => \N__20569\,
            in2 => \_gnd_net_\,
            in3 => \N__20087\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc1_0\,
            ltout => \this_vga_signals.mult1_un47_sum_axbxc1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_x0_LC_19_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18961\,
            in2 => \N__18933\,
            in3 => \N__20409\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_4_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_6_LC_19_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011101110001"
        )
    port map (
            in0 => \N__20411\,
            in1 => \N__22334\,
            in2 => \N__20519\,
            in3 => \N__20570\,
            lcout => \this_vga_signals.g1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_19_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010100001111"
        )
    port map (
            in0 => \N__20571\,
            in1 => \_gnd_net_\,
            in2 => \N__22363\,
            in3 => \N__20513\,
            lcout => \this_vga_signals.vaddress_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_4_LC_19_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21390\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32624\,
            ce => \N__23409\,
            sr => \N__23319\
        );

    \this_ppu.M_haddress_q_RNIOC7O_0_LC_19_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101010100"
        )
    port map (
            in0 => \N__19353\,
            in1 => \N__32075\,
            in2 => \N__31939\,
            in3 => \N__19334\,
            lcout => \M_this_ppu_sprites_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNILR691_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__26187\,
            in1 => \N__21099\,
            in2 => \_gnd_net_\,
            in3 => \N__24158\,
            lcout => \this_start_data_delay.N_993\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_13_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100110000"
        )
    port map (
            in0 => \N__24159\,
            in1 => \N__26188\,
            in2 => \N__20709\,
            in3 => \N__19087\,
            lcout => \M_this_state_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32556\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_15_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__24160\,
            in1 => \N__26189\,
            in2 => \N__19145\,
            in3 => \N__19111\,
            lcout => \M_this_state_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32556\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_o2_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19137\,
            in1 => \N__19110\,
            in2 => \_gnd_net_\,
            in3 => \N__19086\,
            lcout => \this_start_data_delay.N_80_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIHQLO2_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__19068\,
            in1 => \N__26255\,
            in2 => \_gnd_net_\,
            in3 => \N__24157\,
            lcout => \this_start_data_delay.M_this_state_q_ns_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_o2_0_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__19455\,
            in1 => \N__19058\,
            in2 => \_gnd_net_\,
            in3 => \N__23955\,
            lcout => \this_start_data_delay.N_89_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_a2_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19390\,
            in2 => \_gnd_net_\,
            in3 => \N__19059\,
            lcout => OPEN,
            ltout => \this_start_data_delay.un1_M_this_state_q_1_i_a2_0_aZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_external_address_qlde_i_a3_0_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__23956\,
            in1 => \N__19456\,
            in2 => \N__19050\,
            in3 => \N__19047\,
            lcout => \this_start_data_delay.N_122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIA89G3_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__23727\,
            in1 => \N__19763\,
            in2 => \_gnd_net_\,
            in3 => \N__26877\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_127_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_11_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000110010"
        )
    port map (
            in0 => \N__19458\,
            in1 => \N__26218\,
            in2 => \N__19461\,
            in3 => \N__24217\,
            lcout => \M_this_state_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32568\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIP7R11_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19457\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24126\,
            lcout => \N_822_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un30_3_0_o2_1_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__23958\,
            in1 => \N__21089\,
            in2 => \_gnd_net_\,
            in3 => \N__21321\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_844_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIEFRT1_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000001"
        )
    port map (
            in0 => \N__23490\,
            in1 => \N__22163\,
            in2 => \N__19437\,
            in3 => \N__24125\,
            lcout => \this_start_data_delay.N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un1_M_this_substate_q4_2_i_0_303_i_a2_i_a2_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__19423\,
            in1 => \N__19723\,
            in2 => \_gnd_net_\,
            in3 => \N__23491\,
            lcout => \this_start_data_delay.N_151\,
            ltout => \this_start_data_delay.N_151_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un1_M_this_substate_q4_2_i_0_303_i_a2_i_i_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__26183\,
            in1 => \_gnd_net_\,
            in2 => \N__19434\,
            in3 => \N__26867\,
            lcout => \N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIOU691_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__24127\,
            in1 => \N__24309\,
            in2 => \_gnd_net_\,
            in3 => \N__26182\,
            lcout => \N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_o2_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19422\,
            in2 => \_gnd_net_\,
            in3 => \N__19399\,
            lcout => \this_start_data_delay.N_93_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIK0EI1_0_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__19624\,
            in1 => \N__19559\,
            in2 => \N__19706\,
            in3 => \N__19488\,
            lcout => \this_start_data_delay.N_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIOVDB1_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111000000000"
        )
    port map (
            in0 => \N__19625\,
            in1 => \N__19560\,
            in2 => \N__19707\,
            in3 => \N__19968\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_909_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_0_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100111011"
        )
    port map (
            in0 => \N__19934\,
            in1 => \N__19905\,
            in2 => \N__19956\,
            in3 => \N__26212\,
            lcout => led_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32586\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI3F19A_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__19727\,
            in1 => \N__19914\,
            in2 => \N__21117\,
            in3 => \N__26875\,
            lcout => \this_start_data_delay.M_this_state_q_ns_0_i_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIA89G3_0_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19756\,
            in2 => \_gnd_net_\,
            in3 => \N__23664\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_910_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_10_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__24040\,
            in1 => \N__19794\,
            in2 => \N__19767\,
            in3 => \N__26213\,
            lcout => \M_this_state_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32586\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIDHST1_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000001"
        )
    port map (
            in0 => \N__24308\,
            in1 => \N__23776\,
            in2 => \N__19731\,
            in3 => \N__24221\,
            lcout => \this_start_data_delay.M_this_data_count_qlde_i_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIK0EI1_1_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19696\,
            in1 => \N__19629\,
            in2 => \N__19567\,
            in3 => \N__19489\,
            lcout => \this_start_data_delay.N_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_2_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100110000"
        )
    port map (
            in0 => \N__24222\,
            in1 => \N__26209\,
            in2 => \N__19470\,
            in3 => \N__21088\,
            lcout => \M_this_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32592\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_6_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011100"
        )
    port map (
            in0 => \N__24223\,
            in1 => \N__19998\,
            in2 => \N__23795\,
            in3 => \N__26210\,
            lcout => \M_this_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32592\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_22_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111101"
        )
    port map (
            in0 => \N__21871\,
            in1 => \N__20237\,
            in2 => \N__22316\,
            in3 => \N__22533\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_23_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111011"
        )
    port map (
            in0 => \N__20238\,
            in1 => \N__21862\,
            in2 => \N__22327\,
            in3 => \N__21948\,
            lcout => \this_vga_signals.N_4558_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_7_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23429\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32601\,
            ce => \N__23401\,
            sr => \N__23314\
        );

    \this_vga_signals.un5_vaddress_g0_4_i_a3_1_0_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__22531\,
            in1 => \N__21860\,
            in2 => \N__20088\,
            in3 => \N__21946\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_4_i_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_i_1_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011111001111"
        )
    port map (
            in0 => \N__19974\,
            in1 => \N__20239\,
            in2 => \N__19980\,
            in3 => \N__20083\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_4_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_i_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111101001111"
        )
    port map (
            in0 => \N__22532\,
            in1 => \N__21861\,
            in2 => \N__19977\,
            in3 => \N__21947\,
            lcout => \this_vga_signals.N_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_i_o3_1_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__21776\,
            in1 => \N__21813\,
            in2 => \_gnd_net_\,
            in3 => \N__22530\,
            lcout => \this_vga_signals.N_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23428\,
            lcout => \this_vga_signals.M_vcounter_q_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32601\,
            ce => \N__23401\,
            sr => \N__23314\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_x0_LC_20_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21768\,
            in2 => \N__20085\,
            in3 => \N__21812\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_602_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_4_LC_20_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21389\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32610\,
            ce => \N__23408\,
            sr => \N__23316\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001101001"
        )
    port map (
            in0 => \N__21770\,
            in1 => \N__20248\,
            in2 => \N__20147\,
            in3 => \N__20071\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_4_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__20026\,
            in1 => \N__20124\,
            in2 => \_gnd_net_\,
            in3 => \N__21691\,
            lcout => \this_vga_signals.r_N_4_mux\,
            ltout => \this_vga_signals.r_N_4_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIEC471_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011100111"
        )
    port map (
            in0 => \N__21811\,
            in1 => \N__21774\,
            in2 => \N__20154\,
            in3 => \N__22501\,
            lcout => \this_vga_signals.SUM_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_x1_LC_20_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__20027\,
            in1 => \N__21810\,
            in2 => \N__22536\,
            in3 => \N__21692\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a1_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_ns_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__20125\,
            in1 => \_gnd_net_\,
            in2 => \N__20103\,
            in3 => \N__20094\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a1_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a1_x0_LC_20_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21690\,
            in2 => \N__22535\,
            in3 => \N__21806\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a1_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_602_x1_LC_20_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111101111"
        )
    port map (
            in0 => \N__21769\,
            in1 => \N__20070\,
            in2 => \N__21818\,
            in3 => \N__20025\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_602_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_3_x1_LC_20_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000001000"
        )
    port map (
            in0 => \N__22537\,
            in1 => \N__21693\,
            in2 => \N__22044\,
            in3 => \N__23415\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_0_3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_1_LC_20_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011010101001"
        )
    port map (
            in0 => \N__22352\,
            in1 => \N__22997\,
            in2 => \N__23250\,
            in3 => \N__20687\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_26_LC_20_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011010010"
        )
    port map (
            in0 => \N__22998\,
            in1 => \N__23213\,
            in2 => \N__20670\,
            in3 => \N__20662\,
            lcout => \this_vga_signals.N_4_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_5_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101010101"
        )
    port map (
            in0 => \N__22351\,
            in1 => \_gnd_net_\,
            in2 => \N__23249\,
            in3 => \N__22996\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001111001011"
        )
    port map (
            in0 => \N__20601\,
            in1 => \N__20341\,
            in2 => \N__20592\,
            in3 => \N__20418\,
            lcout => \this_vga_signals.mult1_un47_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20551\,
            in2 => \_gnd_net_\,
            in3 => \N__20508\,
            lcout => \this_vga_signals.vaddress_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_1_LC_20_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011011100111"
        )
    port map (
            in0 => \N__22999\,
            in1 => \N__23214\,
            in2 => \N__22404\,
            in3 => \N__20419\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_LC_20_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111010110001"
        )
    port map (
            in0 => \N__20342\,
            in1 => \N__20961\,
            in2 => \N__20301\,
            in3 => \N__20298\,
            lcout => \this_vga_signals.g0_i_x4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_0_a3_1_LC_20_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100101010110"
        )
    port map (
            in0 => \N__22841\,
            in1 => \N__23200\,
            in2 => \N__23093\,
            in3 => \N__22673\,
            lcout => \this_vga_signals.g0_3_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHT721_5_LC_20_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__23073\,
            in1 => \N__23199\,
            in2 => \_gnd_net_\,
            in3 => \N__22356\,
            lcout => \this_vga_signals.vaddress_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNIBR6R_1_LC_20_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__32102\,
            in1 => \N__20955\,
            in2 => \N__31934\,
            in3 => \N__20933\,
            lcout => \M_this_ppu_sprites_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_21_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30106\,
            in1 => \N__20775\,
            in2 => \_gnd_net_\,
            in3 => \N__20760\,
            lcout => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_4_LC_21_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110111010101"
        )
    port map (
            in0 => \N__21045\,
            in1 => \N__27517\,
            in2 => \N__24744\,
            in3 => \N__24708\,
            lcout => \M_this_sprites_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32557\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIK6R81_LC_21_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23472\,
            in1 => \N__23947\,
            in2 => \_gnd_net_\,
            in3 => \N__24164\,
            lcout => \M_this_sprites_ram_write_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNICA9G3_LC_21_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__23731\,
            in1 => \N__20742\,
            in2 => \_gnd_net_\,
            in3 => \N__26876\,
            lcout => \this_start_data_delay.N_125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIOCPV6_0_LC_21_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110111111"
        )
    port map (
            in0 => \N__23799\,
            in1 => \N__23532\,
            in2 => \N__23577\,
            in3 => \N__24609\,
            lcout => OPEN,
            ltout => \this_start_data_delay.un30_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNINS0N8_LC_21_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27822\,
            in2 => \N__20700\,
            in3 => \N__26199\,
            lcout => \this_start_data_delay.N_990\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIHV2L3_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__30573\,
            in1 => \N__28302\,
            in2 => \N__27658\,
            in3 => \N__27603\,
            lcout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__20979\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21009\,
            lcout => \this_start_data_delay.M_last_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32576\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIBJQQ_0_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__21010\,
            in1 => \N__21025\,
            in2 => \_gnd_net_\,
            in3 => \N__20978\,
            lcout => \N_554_0\,
            ltout => \N_554_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIIT6G1_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000100"
        )
    port map (
            in0 => \N__26185\,
            in1 => \N__21101\,
            in2 => \N__21108\,
            in3 => \N__21323\,
            lcout => \this_start_data_delay.N_992\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIIT6G1_0_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110010"
        )
    port map (
            in0 => \N__21324\,
            in1 => \N__26186\,
            in2 => \N__21105\,
            in3 => \N__24161\,
            lcout => \this_start_data_delay.N_109\,
            ltout => \this_start_data_delay.N_109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI433C3_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__28301\,
            in1 => \N__24745\,
            in2 => \N__21048\,
            in3 => \N__25330\,
            lcout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIBOQ11_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21272\,
            in2 => \_gnd_net_\,
            in3 => \N__24128\,
            lcout => \this_start_data_delay.N_86_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIBJQQ_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__21027\,
            in1 => \N__21011\,
            in2 => \_gnd_net_\,
            in3 => \N__20977\,
            lcout => \this_start_data_delay.N_555_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_4_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21036\,
            lcout => \M_this_delay_clk_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIDQQ11_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__21026\,
            in1 => \N__21012\,
            in2 => \N__23798\,
            in3 => \N__20976\,
            lcout => \this_start_data_delay.N_91_0\,
            ltout => \this_start_data_delay.N_91_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI12SC4_0_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28032\,
            in1 => \N__24474\,
            in2 => \N__21327\,
            in3 => \N__32874\,
            lcout => \N_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIKQ691_LC_21_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__24129\,
            in1 => \N__26184\,
            in2 => \_gnd_net_\,
            in3 => \N__21322\,
            lcout => \this_start_data_delay.N_110\,
            ltout => \this_start_data_delay.N_110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI653C3_0_LC_21_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__26308\,
            in1 => \N__32875\,
            in2 => \N__21279\,
            in3 => \N__27645\,
            lcout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI6UUI2_LC_21_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100010"
        )
    port map (
            in0 => \N__24130\,
            in1 => \N__24680\,
            in2 => \N__21276\,
            in3 => \N__23791\,
            lcout => \this_start_data_delay.N_121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21249\,
            in1 => \N__21237\,
            in2 => \_gnd_net_\,
            in3 => \N__30036\,
            lcout => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30035\,
            in1 => \N__21219\,
            in2 => \_gnd_net_\,
            in3 => \N__21204\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_21_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__28727\,
            in1 => \N__28668\,
            in2 => \N__21186\,
            in3 => \N__21183\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_21_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28669\,
            in1 => \N__23583\,
            in2 => \N__21171\,
            in3 => \N__21168\,
            lcout => \M_this_ppu_vram_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI12SC4_1_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000000"
        )
    port map (
            in0 => \N__32892\,
            in1 => \N__28036\,
            in2 => \N__24473\,
            in3 => \N__23827\,
            lcout => \this_start_data_delay.M_this_state_q_ns_0_i_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21537\,
            in1 => \N__21568\,
            in2 => \N__21675\,
            in3 => \N__21674\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_21_20_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            clk => \N__32602\,
            ce => 'H',
            sr => \N__23311\
        );

    \this_vga_signals.M_vcounter_q_1_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21539\,
            in1 => \N__22898\,
            in2 => \_gnd_net_\,
            in3 => \N__21546\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            clk => \N__32602\,
            ce => 'H',
            sr => \N__23311\
        );

    \this_vga_signals.M_vcounter_q_2_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21538\,
            in1 => \N__22648\,
            in2 => \_gnd_net_\,
            in3 => \N__21543\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            clk => \N__32602\,
            ce => 'H',
            sr => \N__23311\
        );

    \this_vga_signals.M_vcounter_q_3_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21540\,
            in1 => \N__22771\,
            in2 => \_gnd_net_\,
            in3 => \N__21393\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            clk => \N__32602\,
            ce => 'H',
            sr => \N__23311\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_21_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23285\,
            in2 => \_gnd_net_\,
            in3 => \N__21357\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23088\,
            in2 => \_gnd_net_\,
            in3 => \N__21336\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22320\,
            in2 => \_gnd_net_\,
            in3 => \N__21333\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_21_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21967\,
            in2 => \_gnd_net_\,
            in3 => \N__21330\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21882\,
            in2 => \_gnd_net_\,
            in3 => \N__22050\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\,
            ltout => OPEN,
            carryin => \bfn_21_21_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_9_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22534\,
            in2 => \_gnd_net_\,
            in3 => \N__22047\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32611\,
            ce => \N__23402\,
            sr => \N__23312\
        );

    \this_vga_signals.M_vcounter_q_esr_8_LC_21_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22031\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32611\,
            ce => \N__23402\,
            sr => \N__23312\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_8_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32611\,
            ce => \N__23402\,
            sr => \N__23312\
        );

    \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22030\,
            lcout => \this_vga_signals.M_vcounter_q_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32611\,
            ce => \N__23402\,
            sr => \N__23312\
        );

    \this_vga_signals.un5_vaddress_g0_17_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111011101"
        )
    port map (
            in0 => \N__21872\,
            in1 => \N__21962\,
            in2 => \_gnd_net_\,
            in3 => \N__22503\,
            lcout => \this_vga_signals.N_4557_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIROQM_8_LC_21_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21963\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21873\,
            lcout => \this_vga_signals.m58_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_601_LC_21_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21814\,
            in2 => \N__21777\,
            in3 => \N__22502\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_6_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21719\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32625\,
            ce => \N__23406\,
            sr => \N__23317\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_7_LC_21_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23433\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32625\,
            ce => \N__23406\,
            sr => \N__23317\
        );

    \this_start_data_delay.M_last_q_RNI75F36_LC_21_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011101"
        )
    port map (
            in0 => \N__26755\,
            in1 => \N__26271\,
            in2 => \N__28275\,
            in3 => \N__26194\,
            lcout => \M_this_external_address_q_3_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI97F36_LC_21_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__23999\,
            in1 => \N__26272\,
            in2 => \N__28166\,
            in3 => \N__26195\,
            lcout => \M_this_external_address_q_3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_21_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__23276\,
            in1 => \N__23089\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.m58_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNICVQL1_1_LC_21_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__22915\,
            in1 => \N__22842\,
            in2 => \N__22709\,
            in3 => \N__22569\,
            lcout => OPEN,
            ltout => \this_vga_signals.m58_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_21_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__22433\,
            in1 => \N__22413\,
            in2 => \N__22407\,
            in3 => \N__22360\,
            lcout => this_vga_signals_vsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI12SC4_2_LC_21_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__32800\,
            in1 => \N__24503\,
            in2 => \N__28044\,
            in3 => \N__23832\,
            lcout => \N_911\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIJARF1_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100110011"
        )
    port map (
            in0 => \N__22179\,
            in1 => \N__23954\,
            in2 => \N__23495\,
            in3 => \N__24204\,
            lcout => \this_start_data_delay.N_123\,
            ltout => \this_start_data_delay.N_123_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIUFEC3_LC_22_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__30935\,
            in1 => \N__24488\,
            in2 => \N__22137\,
            in3 => \N__27979\,
            lcout => \N_812_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_7_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110111010101"
        )
    port map (
            in0 => \N__23508\,
            in1 => \N__27518\,
            in2 => \N__25589\,
            in3 => \N__25554\,
            lcout => \M_this_sprites_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32577\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI213C3_0_LC_22_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__27646\,
            in1 => \N__28471\,
            in2 => \N__25588\,
            in3 => \N__27611\,
            lcout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI12SC4_3_LC_22_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__28014\,
            in1 => \N__32891\,
            in2 => \N__24487\,
            in3 => \N__23820\,
            lcout => \this_start_data_delay.N_938_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI0T8G3_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__23901\,
            in1 => \N__23726\,
            in2 => \_gnd_net_\,
            in3 => \N__26871\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_129_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_8_LC_22_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110100"
        )
    port map (
            in0 => \N__24163\,
            in1 => \N__23474\,
            in2 => \N__23502\,
            in3 => \N__26223\,
            lcout => \M_this_state_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIJ13L3_LC_22_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__27607\,
            in1 => \N__24458\,
            in2 => \N__30677\,
            in3 => \N__27657\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_12_LC_22_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111110001111"
        )
    port map (
            in0 => \N__27533\,
            in1 => \N__30657\,
            in2 => \N__23499\,
            in3 => \N__25395\,
            lcout => \M_this_sprites_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIFSQ11_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23473\,
            in2 => \_gnd_net_\,
            in3 => \N__24162\,
            lcout => \this_start_data_delay.N_821_0\,
            ltout => \this_start_data_delay.N_821_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_9_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23436\,
            in3 => \N__26224\,
            lcout => \M_this_state_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_11_LC_22_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110111010101"
        )
    port map (
            in0 => \N__23625\,
            in1 => \N__27532\,
            in2 => \N__30592\,
            in3 => \N__25404\,
            lcout => \M_this_sprites_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32588\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIFT2L3_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__27602\,
            in1 => \N__25435\,
            in2 => \N__31342\,
            in3 => \N__27653\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_10_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111110001111"
        )
    port map (
            in0 => \N__25434\,
            in1 => \N__27557\,
            in2 => \N__23619\,
            in3 => \N__25413\,
            lcout => \M_this_sprites_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32593\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_22_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23616\,
            in1 => \N__23598\,
            in2 => \_gnd_net_\,
            in3 => \N__30056\,
            lcout => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIL33L3_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__30480\,
            in1 => \N__28127\,
            in2 => \N__27659\,
            in3 => \N__27601\,
            lcout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIOCPV6_LC_22_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__23796\,
            in1 => \N__24608\,
            in2 => \N__23572\,
            in3 => \N__23531\,
            lcout => un30_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI0V2C3_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__25033\,
            in1 => \N__25300\,
            in2 => \N__32903\,
            in3 => \N__25352\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_2_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111110001111"
        )
    port map (
            in0 => \N__25032\,
            in1 => \N__27558\,
            in2 => \N__23514\,
            in3 => \N__25008\,
            lcout => \M_this_sprites_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI0T8G3_0_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23889\,
            in2 => \_gnd_net_\,
            in3 => \N__23652\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_913_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_7_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__26222\,
            in1 => \N__24622\,
            in2 => \N__23511\,
            in3 => \N__23957\,
            lcout => \M_this_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI213C3_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__24889\,
            in1 => \N__25301\,
            in2 => \N__31355\,
            in3 => \N__25353\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_3_LC_22_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111110001111"
        )
    port map (
            in0 => \N__24888\,
            in1 => \N__27559\,
            in2 => \N__23868\,
            in3 => \N__24864\,
            lcout => \M_this_sprites_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_13_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31919\,
            in1 => \N__32141\,
            in2 => \N__23865\,
            in3 => \N__23841\,
            lcout => \this_sprites_ram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI12SC4_LC_22_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000000000000"
        )
    port map (
            in0 => \N__32858\,
            in1 => \N__24445\,
            in2 => \N__28040\,
            in3 => \N__23828\,
            lcout => \this_start_data_delay.N_149\,
            ltout => \this_start_data_delay.N_149_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIF2NL5_LC_22_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__24281\,
            in1 => \N__24178\,
            in2 => \N__23802\,
            in3 => \N__23797\,
            lcout => \this_start_data_delay.M_this_data_count_qlde_i_2_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNITK893_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23732\,
            in2 => \_gnd_net_\,
            in3 => \N__26851\,
            lcout => \this_start_data_delay.N_820_0\,
            ltout => \this_start_data_delay.N_820_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI281SC_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110101"
        )
    port map (
            in0 => \N__23694\,
            in1 => \N__23685\,
            in2 => \N__23679\,
            in3 => \N__23676\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_data_count_qlde_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIC4IPK_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100101111"
        )
    port map (
            in0 => \N__24647\,
            in1 => \N__23656\,
            in2 => \N__23628\,
            in3 => \N__26201\,
            lcout => \N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_5_LC_22_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__24327\,
            in1 => \N__24179\,
            in2 => \N__24301\,
            in3 => \N__26202\,
            lcout => \M_this_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_d62_11_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28910\,
            in1 => \N__28939\,
            in2 => \N__28886\,
            in3 => \N__29136\,
            lcout => \this_start_data_delay.M_this_state_d62Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_5_LC_22_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__29195\,
            in1 => \N__28926\,
            in2 => \_gnd_net_\,
            in3 => \N__28940\,
            lcout => \M_this_data_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32618\,
            ce => \N__29104\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_7_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__28866\,
            in1 => \N__29196\,
            in2 => \_gnd_net_\,
            in3 => \N__28882\,
            lcout => \M_this_data_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32618\,
            ce => \N__29104\,
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIOU691_0_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__24285\,
            in1 => \N__26198\,
            in2 => \_gnd_net_\,
            in3 => \N__24226\,
            lcout => OPEN,
            ltout => \this_start_data_delay_M_this_data_count_q_3_0_a3_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_6_LC_22_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__28899\,
            in1 => \N__26765\,
            in2 => \N__24051\,
            in3 => \N__29194\,
            lcout => \M_this_data_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32618\,
            ce => \N__29104\,
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNII9RA6_LC_22_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__24019\,
            in1 => \N__26971\,
            in2 => \N__32884\,
            in3 => \N__26197\,
            lcout => \M_this_data_count_q_3_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_13_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001000100111"
        )
    port map (
            in0 => \N__29235\,
            in1 => \N__23970\,
            in2 => \N__29859\,
            in3 => \N__29879\,
            lcout => \M_this_data_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32626\,
            ce => \N__29081\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_9_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__29979\,
            in1 => \N__26974\,
            in2 => \N__30914\,
            in3 => \N__29234\,
            lcout => \M_this_data_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32626\,
            ce => \N__29081\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_8_LC_22_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__28833\,
            in1 => \N__26973\,
            in2 => \N__28470\,
            in3 => \N__29233\,
            lcout => \M_this_data_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32626\,
            ce => \N__29081\,
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un1_M_this_substate_q4_1_i_0_286_i_i_LC_22_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26192\,
            in2 => \_gnd_net_\,
            in3 => \N__24690\,
            lcout => \N_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIEGBV8_LC_22_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24669\,
            in1 => \N__26193\,
            in2 => \N__24654\,
            in3 => \N__24636\,
            lcout => \N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNINT691_LC_22_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26270\,
            in2 => \_gnd_net_\,
            in3 => \N__26190\,
            lcout => \M_this_external_address_d_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI86F36_LC_22_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010111111"
        )
    port map (
            in0 => \N__26191\,
            in1 => \N__26273\,
            in2 => \N__24498\,
            in3 => \N__24623\,
            lcout => \M_this_external_address_q_3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNISDEC3_LC_23_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__28419\,
            in1 => \N__27980\,
            in2 => \N__28320\,
            in3 => \N__27823\,
            lcout => \N_813_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI653C3_LC_23_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__27069\,
            in1 => \N__25302\,
            in2 => \N__24497\,
            in3 => \N__25343\,
            lcout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI873C3_LC_23_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__25345\,
            in1 => \N__28109\,
            in2 => \N__25313\,
            in3 => \N__25720\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_6_LC_23_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111110001111"
        )
    port map (
            in0 => \N__25719\,
            in1 => \N__27543\,
            in2 => \N__24330\,
            in3 => \N__25698\,
            lcout => \M_this_sprites_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIUS2C3_LC_23_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__25346\,
            in1 => \N__30930\,
            in2 => \N__25314\,
            in3 => \N__25168\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_1_LC_23_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111100001111"
        )
    port map (
            in0 => \N__25167\,
            in1 => \N__25146\,
            in2 => \N__25356\,
            in3 => \N__27542\,
            lcout => \M_this_sprites_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNISQ2C3_LC_23_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__25344\,
            in1 => \N__28472\,
            in2 => \N__25312\,
            in3 => \N__26457\,
            lcout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_0_c_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25367\,
            in2 => \N__26459\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_23_17_0_\,
            carryout => \un1_M_this_sprites_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_0_THRU_LUT4_0_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25175\,
            in3 => \N__25140\,
            lcout => \un1_M_this_sprites_address_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_0\,
            carryout => \un1_M_this_sprites_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_1_THRU_LUT4_0_LC_23_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25040\,
            in2 => \_gnd_net_\,
            in3 => \N__24999\,
            lcout => \un1_M_this_sprites_address_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_1\,
            carryout => \un1_M_this_sprites_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_2_THRU_LUT4_0_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24902\,
            in2 => \_gnd_net_\,
            in3 => \N__24855\,
            lcout => \un1_M_this_sprites_address_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_2\,
            carryout => \un1_M_this_sprites_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_3_THRU_LUT4_0_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24752\,
            in2 => \_gnd_net_\,
            in3 => \N__24696\,
            lcout => \un1_M_this_sprites_address_q_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_3\,
            carryout => \un1_M_this_sprites_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_4_THRU_LUT4_0_LC_23_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27070\,
            in2 => \_gnd_net_\,
            in3 => \N__24693\,
            lcout => \un1_M_this_sprites_address_q_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_4\,
            carryout => \un1_M_this_sprites_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_5_THRU_LUT4_0_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25721\,
            in2 => \_gnd_net_\,
            in3 => \N__25692\,
            lcout => \un1_M_this_sprites_address_q_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_5\,
            carryout => \un1_M_this_sprites_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_6_THRU_LUT4_0_LC_23_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25578\,
            in2 => \_gnd_net_\,
            in3 => \N__25548\,
            lcout => \un1_M_this_sprites_address_q_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_6\,
            carryout => \un1_M_this_sprites_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_7_THRU_LUT4_0_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27380\,
            in2 => \_gnd_net_\,
            in3 => \N__25545\,
            lcout => \un1_M_this_sprites_address_q_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_23_18_0_\,
            carryout => \un1_M_this_sprites_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_8_THRU_LUT4_0_LC_23_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26301\,
            in2 => \_gnd_net_\,
            in3 => \N__25542\,
            lcout => \un1_M_this_sprites_address_q_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_8\,
            carryout => \un1_M_this_sprites_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_9_THRU_LUT4_0_LC_23_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25436\,
            in2 => \_gnd_net_\,
            in3 => \N__25407\,
            lcout => \un1_M_this_sprites_address_q_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_9\,
            carryout => \un1_M_this_sprites_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_10_THRU_LUT4_0_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30572\,
            in2 => \_gnd_net_\,
            in3 => \N__25398\,
            lcout => \un1_M_this_sprites_address_q_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_10\,
            carryout => \un1_M_this_sprites_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_11_THRU_LUT4_0_LC_23_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30653\,
            in2 => \_gnd_net_\,
            in3 => \N__25389\,
            lcout => \un1_M_this_sprites_address_q_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_11\,
            carryout => \un1_M_this_sprites_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_13_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101110110011"
        )
    port map (
            in0 => \N__27562\,
            in1 => \N__25386\,
            in2 => \N__30513\,
            in3 => \N__25380\,
            lcout => \M_this_sprites_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_0_LC_23_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110111010101"
        )
    port map (
            in0 => \N__25377\,
            in1 => \N__27561\,
            in2 => \N__26458\,
            in3 => \N__25368\,
            lcout => \M_this_sprites_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_9_LC_23_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101110110011"
        )
    port map (
            in0 => \N__27563\,
            in1 => \N__26424\,
            in2 => \N__26309\,
            in3 => \N__26415\,
            lcout => \M_this_sprites_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI96JM1_LC_23_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__27933\,
            in1 => \N__26274\,
            in2 => \_gnd_net_\,
            in3 => \N__26200\,
            lcout => \this_start_data_delay_M_this_external_address_q_3_i_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25851\,
            in1 => \N__25839\,
            in2 => \_gnd_net_\,
            in3 => \N__30088\,
            lcout => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_12_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__29226\,
            in1 => \N__29892\,
            in2 => \N__28294\,
            in3 => \N__26975\,
            lcout => \M_this_data_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32619\,
            ce => \N__29109\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_0_LC_23_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29225\,
            in2 => \_gnd_net_\,
            in3 => \N__28512\,
            lcout => \M_this_data_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32619\,
            ce => \N__29109\,
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_d62_10_LC_23_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29020\,
            in1 => \N__28492\,
            in2 => \N__28995\,
            in3 => \N__28510\,
            lcout => \this_start_data_delay.M_this_state_d62Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_15_LC_23_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__29256\,
            in1 => \N__26972\,
            in2 => \N__27941\,
            in3 => \N__29227\,
            lcout => \M_this_data_count_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32627\,
            ce => \N__29101\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_1_LC_23_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__28493\,
            in1 => \_gnd_net_\,
            in2 => \N__29238\,
            in3 => \N__28479\,
            lcout => \M_this_data_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32627\,
            ce => \N__29101\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_2_LC_23_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__29021\,
            in1 => \N__29007\,
            in2 => \_gnd_net_\,
            in3 => \N__29231\,
            lcout => \M_this_data_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32627\,
            ce => \N__29101\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_11_LC_23_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__29236\,
            in1 => \N__29922\,
            in2 => \N__26979\,
            in3 => \N__31296\,
            lcout => \M_this_data_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32632\,
            ce => \N__29085\,
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_d62_8_LC_23_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29959\,
            in1 => \N__28817\,
            in2 => \N__29937\,
            in3 => \N__28844\,
            lcout => \this_start_data_delay.M_this_state_d62Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_d62_9_LC_23_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29315\,
            in1 => \N__29875\,
            in2 => \N__29274\,
            in3 => \N__29909\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_state_d62Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_d62_LC_23_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26898\,
            in1 => \N__26892\,
            in2 => \N__26886\,
            in3 => \N__26883\,
            lcout => \this_start_data_delay.M_this_state_dZ0Z62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_10_LC_23_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010011001"
        )
    port map (
            in0 => \N__29960\,
            in1 => \N__29946\,
            in2 => \N__26811\,
            in3 => \N__29237\,
            lcout => \M_this_data_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32632\,
            ce => \N__29085\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_8_LC_23_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__30969\,
            in1 => \N__32932\,
            in2 => \N__28455\,
            in3 => \N__32735\,
            lcout => \M_this_external_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32641\,
            ce => \N__32220\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_15_LC_23_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__26802\,
            in1 => \N__26787\,
            in2 => \N__31377\,
            in3 => \N__32734\,
            lcout => \M_this_external_address_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32641\,
            ce => \N__32220\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_13_LC_23_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010010111110"
        )
    port map (
            in0 => \N__32733\,
            in1 => \N__31486\,
            in2 => \N__31467\,
            in3 => \N__26703\,
            lcout => \M_this_external_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32641\,
            ce => \N__32220\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI5F621_2_LC_23_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__26697\,
            in1 => \N__26676\,
            in2 => \N__31964\,
            in3 => \N__32131\,
            lcout => \M_this_ppu_sprites_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__30519\,
            in1 => \N__30606\,
            in2 => \N__30697\,
            in3 => \N__30751\,
            lcout => \this_sprites_ram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__30752\,
            in1 => \N__30520\,
            in2 => \N__30614\,
            in3 => \N__30681\,
            lcout => \this_sprites_ram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__30754\,
            in1 => \N__30685\,
            in2 => \N__30526\,
            in3 => \N__30594\,
            lcout => \this_sprites_ram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__30593\,
            in1 => \N__30515\,
            in2 => \N__30698\,
            in3 => \N__30753\,
            lcout => \this_sprites_ram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI0IEC3_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__32904\,
            in1 => \N__27984\,
            in2 => \N__28108\,
            in3 => \N__27830\,
            lcout => \N_811_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_5_LC_24_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110111010101"
        )
    port map (
            in0 => \N__27186\,
            in1 => \N__27560\,
            in2 => \N__27074\,
            in3 => \N__27180\,
            lcout => \M_this_sprites_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__30481\,
            in1 => \N__30591\,
            in2 => \N__30699\,
            in3 => \N__30739\,
            lcout => \this_sprites_ram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_24_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27018\,
            in1 => \N__27006\,
            in2 => \_gnd_net_\,
            in3 => \N__30105\,
            lcout => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_3_0_LC_24_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28473\,
            in1 => \N__28285\,
            in2 => \N__30936\,
            in3 => \N__28096\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_ns_0_o4_0_a2_4_a2_4_o2_0_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27916\,
            in2 => \N__28047\,
            in3 => \N__31323\,
            lcout => \this_start_data_delay.N_902_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI2KEC3_LC_24_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__31322\,
            in1 => \N__27978\,
            in2 => \N__27929\,
            in3 => \N__27834\,
            lcout => \N_41_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_24_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30089\,
            in1 => \N__27732\,
            in2 => \_gnd_net_\,
            in3 => \N__27726\,
            lcout => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_24_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30090\,
            in1 => \N__27711\,
            in2 => \_gnd_net_\,
            in3 => \N__27705\,
            lcout => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_24_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30091\,
            in1 => \N__27687\,
            in2 => \_gnd_net_\,
            in3 => \N__27675\,
            lcout => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI433C3_0_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__27379\,
            in1 => \N__27663\,
            in2 => \N__30934\,
            in3 => \N__27612\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_sprites_address_q_0_0_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_8_LC_24_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111100001111"
        )
    port map (
            in0 => \N__27378\,
            in1 => \N__27573\,
            in2 => \N__27567\,
            in3 => \N__27564\,
            lcout => \M_this_sprites_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__28667\,
            in1 => \N__27354\,
            in2 => \N__28728\,
            in3 => \N__28806\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__28676\,
            in1 => \N__29991\,
            in2 => \N__28800\,
            in3 => \N__28797\,
            lcout => \M_this_ppu_vram_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30076\,
            in1 => \N__28755\,
            in2 => \_gnd_net_\,
            in3 => \N__28743\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__28720\,
            in1 => \N__28686\,
            in2 => \N__28680\,
            in3 => \N__28666\,
            lcout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_24_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30095\,
            in1 => \N__28614\,
            in2 => \_gnd_net_\,
            in3 => \N__28602\,
            lcout => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__30755\,
            in1 => \N__30514\,
            in2 => \N__30704\,
            in3 => \N__30605\,
            lcout => \this_sprites_ram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28554\,
            in1 => \N__28539\,
            in2 => \_gnd_net_\,
            in3 => \N__30096\,
            lcout => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_c_0_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28511\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_24_21_0_\,
            carryout => \M_this_data_count_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_0_THRU_LUT4_0_LC_24_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28494\,
            in2 => \N__29682\,
            in3 => \N__29025\,
            lcout => \M_this_data_count_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_0\,
            carryout => \M_this_data_count_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_1_THRU_LUT4_0_LC_24_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29022\,
            in2 => \N__29680\,
            in3 => \N__28998\,
            lcout => \M_this_data_count_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_1\,
            carryout => \M_this_data_count_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_2_THRU_LUT4_0_LC_24_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28994\,
            in2 => \N__29683\,
            in3 => \N__28950\,
            lcout => \M_this_data_count_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_2\,
            carryout => \M_this_data_count_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_3_THRU_LUT4_0_LC_24_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29135\,
            in2 => \N__29681\,
            in3 => \N__28947\,
            lcout => \M_this_data_count_q_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_3\,
            carryout => \M_this_data_count_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_4_THRU_LUT4_0_LC_24_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28944\,
            in2 => \N__29684\,
            in3 => \N__28917\,
            lcout => \M_this_data_count_q_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_4\,
            carryout => \M_this_data_count_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_6_LC_24_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28914\,
            in2 => \N__29679\,
            in3 => \N__28890\,
            lcout => \M_this_data_count_q_s_6\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_5\,
            carryout => \M_this_data_count_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_6_THRU_LUT4_0_LC_24_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28887\,
            in2 => \N__29685\,
            in3 => \N__28857\,
            lcout => \M_this_data_count_q_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_6\,
            carryout => \M_this_data_count_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_8_LC_24_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29691\,
            in2 => \N__28854\,
            in3 => \N__28824\,
            lcout => \M_this_data_count_q_s_8\,
            ltout => OPEN,
            carryin => \bfn_24_22_0_\,
            carryout => \M_this_data_count_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_9_LC_24_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28821\,
            in2 => \N__29752\,
            in3 => \N__29970\,
            lcout => \M_this_data_count_q_s_9\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_8\,
            carryout => \M_this_data_count_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_9_THRU_LUT4_0_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29698\,
            in2 => \N__29967\,
            in3 => \N__29940\,
            lcout => \M_this_data_count_q_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_9\,
            carryout => \M_this_data_count_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_11_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29936\,
            in2 => \N__29751\,
            in3 => \N__29916\,
            lcout => \M_this_data_count_q_s_11\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_10\,
            carryout => \M_this_data_count_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_12_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29689\,
            in2 => \N__29913\,
            in3 => \N__29883\,
            lcout => \M_this_data_count_q_s_12\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_11\,
            carryout => \M_this_data_count_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_12_THRU_LUT4_0_LC_24_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29880\,
            in2 => \N__29753\,
            in3 => \N__29847\,
            lcout => \M_this_data_count_q_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_12\,
            carryout => \M_this_data_count_q_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_14_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29690\,
            in2 => \N__29319\,
            in3 => \N__29277\,
            lcout => \M_this_data_count_q_s_14\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_13\,
            carryout => \M_this_data_count_q_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_15_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29273\,
            in2 => \_gnd_net_\,
            in3 => \N__29259\,
            lcout => \M_this_data_count_q_s_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_4_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__29247\,
            in1 => \N__29232\,
            in2 => \_gnd_net_\,
            in3 => \N__29131\,
            lcout => \M_this_data_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32642\,
            ce => \N__29102\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_12_LC_24_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101011010"
        )
    port map (
            in0 => \N__31512\,
            in1 => \N__30954\,
            in2 => \N__31538\,
            in3 => \N__32760\,
            lcout => \M_this_external_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32644\,
            ce => \N__32235\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_14_LC_24_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111000010100"
        )
    port map (
            in0 => \N__32758\,
            in1 => \N__31416\,
            in2 => \N__31442\,
            in3 => \N__30945\,
            lcout => \M_this_external_address_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32644\,
            ce => \N__32235\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_9_LC_24_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__31560\,
            in1 => \N__32941\,
            in2 => \N__30915\,
            in3 => \N__32759\,
            lcout => \M_this_external_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32644\,
            ce => \N__32235\,
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__30527\,
            in1 => \N__30610\,
            in2 => \N__30705\,
            in3 => \N__30761\,
            lcout => \this_sprites_ram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30762\,
            in1 => \N__30700\,
            in2 => \N__30615\,
            in3 => \N__30528\,
            lcout => \this_sprites_ram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIP0T41_2_LC_24_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__32129\,
            in1 => \N__31960\,
            in2 => \N__30429\,
            in3 => \N__30405\,
            lcout => \M_this_ppu_sprites_addr_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNI2HC01_2_LC_24_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__30291\,
            in1 => \N__32128\,
            in2 => \N__31969\,
            in3 => \N__30249\,
            lcout => \M_this_ppu_sprites_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_26_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30135\,
            in1 => \N__30117\,
            in2 => \_gnd_net_\,
            in3 => \N__30107\,
            lcout => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_0_LC_26_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32752\,
            in1 => \N__31178\,
            in2 => \_gnd_net_\,
            in3 => \N__31167\,
            lcout => \M_this_external_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_26_23_0_\,
            carryout => \M_this_external_address_q_cry_0\,
            clk => \N__32648\,
            ce => \N__32233\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_1_LC_26_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32748\,
            in1 => \N__31157\,
            in2 => \_gnd_net_\,
            in3 => \N__31146\,
            lcout => \M_this_external_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_0\,
            carryout => \M_this_external_address_q_cry_1\,
            clk => \N__32648\,
            ce => \N__32233\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_2_LC_26_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32753\,
            in1 => \N__31130\,
            in2 => \_gnd_net_\,
            in3 => \N__31119\,
            lcout => \M_this_external_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_1\,
            carryout => \M_this_external_address_q_cry_2\,
            clk => \N__32648\,
            ce => \N__32233\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_3_LC_26_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32749\,
            in1 => \N__31103\,
            in2 => \_gnd_net_\,
            in3 => \N__31092\,
            lcout => \M_this_external_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_2\,
            carryout => \M_this_external_address_q_cry_3\,
            clk => \N__32648\,
            ce => \N__32233\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_4_LC_26_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32754\,
            in1 => \N__31085\,
            in2 => \_gnd_net_\,
            in3 => \N__31074\,
            lcout => \M_this_external_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_3\,
            carryout => \M_this_external_address_q_cry_4\,
            clk => \N__32648\,
            ce => \N__32233\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_5_LC_26_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32750\,
            in1 => \N__31061\,
            in2 => \_gnd_net_\,
            in3 => \N__31050\,
            lcout => \M_this_external_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_4\,
            carryout => \M_this_external_address_q_cry_5\,
            clk => \N__32648\,
            ce => \N__32233\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_6_LC_26_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32755\,
            in1 => \N__31040\,
            in2 => \_gnd_net_\,
            in3 => \N__31029\,
            lcout => \M_this_external_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_5\,
            carryout => \M_this_external_address_q_cry_6\,
            clk => \N__32648\,
            ce => \N__32233\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_7_LC_26_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32751\,
            in1 => \N__31010\,
            in2 => \_gnd_net_\,
            in3 => \N__30999\,
            lcout => \M_this_external_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_6\,
            carryout => \M_this_external_address_q_cry_7\,
            clk => \N__32648\,
            ce => \N__32233\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_RNO_0_8_LC_26_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30986\,
            in2 => \_gnd_net_\,
            in3 => \N__30957\,
            lcout => \M_this_external_address_q_s_8\,
            ltout => OPEN,
            carryin => \bfn_26_24_0_\,
            carryout => \M_this_external_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_RNO_0_9_LC_26_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31577\,
            in2 => \_gnd_net_\,
            in3 => \N__31551\,
            lcout => \M_this_external_address_q_s_9\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_8\,
            carryout => \M_this_external_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_RNO_0_10_LC_26_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32675\,
            in2 => \_gnd_net_\,
            in3 => \N__31548\,
            lcout => \M_this_external_address_q_s_10\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_9\,
            carryout => \M_this_external_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_RNO_0_11_LC_26_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31202\,
            in2 => \_gnd_net_\,
            in3 => \N__31545\,
            lcout => \M_this_external_address_q_s_11\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_10\,
            carryout => \M_this_external_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_cry_11_THRU_LUT4_0_LC_26_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31537\,
            in2 => \_gnd_net_\,
            in3 => \N__31503\,
            lcout => \M_this_external_address_q_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_11\,
            carryout => \M_this_external_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_cry_12_THRU_LUT4_0_LC_26_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31490\,
            in2 => \_gnd_net_\,
            in3 => \N__31455\,
            lcout => \M_this_external_address_q_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_12\,
            carryout => \M_this_external_address_q_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_cry_13_THRU_LUT4_0_LC_26_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31441\,
            in2 => \_gnd_net_\,
            in3 => \N__31407\,
            lcout => \M_this_external_address_q_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_13\,
            carryout => \M_this_external_address_q_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_RNO_0_15_LC_26_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31397\,
            in2 => \_gnd_net_\,
            in3 => \N__31380\,
            lcout => \M_this_external_address_q_s_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_11_LC_26_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__32756\,
            in1 => \N__31365\,
            in2 => \N__31295\,
            in3 => \N__32949\,
            lcout => \M_this_external_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32654\,
            ce => \N__32234\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_10_LC_26_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__32955\,
            in1 => \N__32948\,
            in2 => \N__32819\,
            in3 => \N__32757\,
            lcout => \M_this_external_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32654\,
            ce => \N__32234\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIVCB01_1_LC_26_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__32187\,
            in1 => \N__32130\,
            in2 => \N__31970\,
            in3 => \N__31806\,
            lcout => \M_this_ppu_sprites_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un1_M_this_state_q_17_i_o2_1_4_LC_32_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31689\,
            in1 => \N__31668\,
            in2 => \N__31656\,
            in3 => \N__31608\,
            lcout => \this_start_data_delay.un1_M_this_state_q_17_i_o2_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
