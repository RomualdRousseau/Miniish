-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     May 21 2022 22:52:11

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : inout std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    debug : out std_logic_vector(1 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : inout std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__25733\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \VCCG0\ : std_logic;
signal \this_vga_signals.N_517_1\ : std_logic;
signal \N_205_i\ : std_logic;
signal \this_vga_ramdac.M_this_rgb_d_3_0_dreg\ : std_logic;
signal \this_vga_ramdac.m5_cascade_\ : std_logic;
signal \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_0\ : std_logic;
signal \this_vga_ramdac.m16\ : std_logic;
signal \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_2\ : std_logic;
signal \this_vga_ramdac.m19\ : std_logic;
signal \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_3\ : std_logic;
signal \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_1\ : std_logic;
signal \this_vga_ramdac.i2_mux\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \this_vga_ramdac.N_706_0\ : std_logic;
signal \this_vga_ramdac.i2_mux_0\ : std_logic;
signal \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_4\ : std_logic;
signal \N_94\ : std_logic;
signal \N_274_i\ : std_logic;
signal \this_vga_signals.if_N_6_mux_0_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_8\ : std_logic;
signal \M_this_vga_signals_address_11\ : std_logic;
signal \this_vga_signals.g0_0_a2_1\ : std_logic;
signal \M_this_vga_signals_address_9\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.g2_0_x1\ : std_logic;
signal \this_vga_signals.g2_0_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0_0\ : std_logic;
signal \this_vga_signals.g2_0\ : std_logic;
signal \M_this_vga_signals_address_12\ : std_logic;
signal \this_vga_signals.g0_2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_1\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_cry_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_cry_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_cry_2\ : std_logic;
signal \N_70_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_cry_1_THRU_CO\ : std_logic;
signal \G_501\ : std_logic;
signal \N_70\ : std_logic;
signal \N_26\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_cry_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_cry_1_s\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_cry_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axb_3\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_cry_2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb_2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb_1_l_fx\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_cry_2_THRU_CO\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_s_3\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_cry_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_cry_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_cry_2\ : std_logic;
signal \this_vga_signals.N_70_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_i_3\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_cry_1_s\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_cry_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_cry_1_s\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb_3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_cry_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb_3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_cry_2\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_s_3\ : std_logic;
signal \this_vga_signals.M_hcounter_q_i_0_5\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_s_3\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_i_3\ : std_logic;
signal \this_ppu.M_N_6_0_cascade_\ : std_logic;
signal \this_ppu.M_N_13_mux\ : std_logic;
signal \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_c_0\ : std_logic;
signal \this_ppu.M_N_15_mux_cascade_\ : std_logic;
signal \this_ppu.M_m12_0_x3_s_0_1Z0Z_0_cascade_\ : std_logic;
signal \this_ppu.M_m12_0_x3_out_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m12_cascade_\ : std_logic;
signal \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_c3_0_cascade_\ : std_logic;
signal \this_ppu.N_277\ : std_logic;
signal \this_ppu.M_mZ0Z1_cascade_\ : std_logic;
signal \N_92\ : std_logic;
signal \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axb1_cascade_\ : std_logic;
signal this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_c3_0 : std_logic;
signal this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axb1 : std_logic;
signal \this_ppu.M_N_16_1_cascade_\ : std_logic;
signal \this_ppu.M_m9_i_x3Z0Z_0\ : std_logic;
signal \this_ppu.M_mZ0Z1\ : std_logic;
signal \this_ppu.M_m1_e_0_1_0_cascade_\ : std_logic;
signal \this_ppu.M_m1_e_0_1_1\ : std_logic;
signal \this_ppu.M_m12_0_x3_out_0\ : std_logic;
signal \this_ppu.M_N_16_1\ : std_logic;
signal \this_ppu.M_m1_e_0_0\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \this_ppu.un1_M_current_q_cry_0\ : std_logic;
signal \this_ppu.un1_M_current_q_cry_1\ : std_logic;
signal \this_ppu.un1_M_current_q_cry_2\ : std_logic;
signal \this_ppu.un1_M_current_q_cry_3\ : std_logic;
signal \this_ppu.un1_M_current_q_cry_4\ : std_logic;
signal \this_ppu.un1_M_current_q_cry_5\ : std_logic;
signal \this_ppu.N_256_1_i\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_0\ : std_logic;
signal \M_this_vga_signals_address_10\ : std_logic;
signal \this_vga_signals.N_9_0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3Z0Z_5_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_0Z0Z_5\ : std_logic;
signal \this_vga_signals.N_5\ : std_logic;
signal \this_vga_signals.g0_0_x2_0_0_a3_3_cascade_\ : std_logic;
signal \this_vga_signals.N_9_i_0_0_cascade_\ : std_logic;
signal \this_vga_signals.N_9_i_0_0\ : std_logic;
signal \this_vga_signals.g0_2_x0_cascade_\ : std_logic;
signal \this_vga_signals.g0_2_x1\ : std_logic;
signal \this_vga_signals.N_3_1\ : std_logic;
signal \this_vga_signals.m6_2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_0_0\ : std_logic;
signal \this_vga_signals.if_i3_mux_0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNI820378Z0Z_2\ : std_logic;
signal \this_vga_signals.N_3_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNI820378_0Z0Z_2\ : std_logic;
signal \this_vga_signals.g0_3_0_a3_2_cascade_\ : std_logic;
signal \this_vga_signals.g2_1\ : std_logic;
signal \this_vga_signals.g1_0_0_0\ : std_logic;
signal \this_vga_signals.N_188_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m10_0_a4_0_0\ : std_logic;
signal \this_vga_signals.g1_3_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m10_0_a4_1_1\ : std_logic;
signal \this_vga_signals.if_N_18_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_1_0_0\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_9\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_x1_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_x0_3\ : std_logic;
signal \this_vga_signals.CO1_5_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum0_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_ns_2_cascade_\ : std_logic;
signal \this_vga_signals.N_196_0\ : std_logic;
signal \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0_cascade_\ : std_logic;
signal this_vga_signals_un4_lcounter_if_generate_plus_mult1_un54_sum_axb1 : std_logic;
signal \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un54_sum_axb1_cascade_\ : std_logic;
signal this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_c3_0 : std_logic;
signal \this_vga_signals_un4_lcounter_if_i1_mux_cascade_\ : std_logic;
signal this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0 : std_logic;
signal \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_cascade_\ : std_logic;
signal this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_1 : std_logic;
signal \this_ppu.M_m7Z0Z_1\ : std_logic;
signal \this_ppu.M_m12_0_o2_381_10Z0Z_1\ : std_logic;
signal \this_ppu.M_N_11_mux_cascade_\ : std_logic;
signal \this_ppu.M_m12_0_o2_381_10\ : std_logic;
signal this_vga_signals_un4_lcounter_if_i1_mux : std_logic;
signal this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1 : std_logic;
signal this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_1 : std_logic;
signal \this_vga_signals_un4_lcounter_if_N_7_i_i\ : std_logic;
signal \M_this_ppu_vram_addr_5\ : std_logic;
signal \M_this_ppu_vram_addr_4\ : std_logic;
signal \M_this_ppu_vram_addr_6\ : std_logic;
signal \M_this_ppu_vram_addr_2\ : std_logic;
signal \this_ppu.un1_M_state_d8_4_0_cascade_\ : std_logic;
signal \this_ppu.M_N_3_mux_0_0\ : std_logic;
signal \M_this_ppu_vram_addr_0\ : std_logic;
signal \M_this_ppu_vram_addr_3\ : std_logic;
signal \M_this_ppu_vram_addr_1\ : std_logic;
signal \this_ppu.un1_M_state_d8_5_0\ : std_logic;
signal \M_this_sprites_ram_read_data_0_cascade_\ : std_logic;
signal \M_this_vram_write_data_0\ : std_logic;
signal port_clk_c : std_logic;
signal \this_vga_signals.vsync_1_0_a2_6_a2_1_0\ : std_logic;
signal this_vga_signals_vsync_1_i : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_0\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_1\ : std_logic;
signal \this_vga_signals.g0_16_x0_cascade_\ : std_logic;
signal \this_vga_signals.g3_0\ : std_logic;
signal \this_vga_signals.N_57_i_i_0_0\ : std_logic;
signal \this_vga_signals.g0_1_0_cascade_\ : std_logic;
signal \this_vga_signals.N_5_0_0_1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_3_0_0_0_cascade_\ : std_logic;
signal this_vga_signals_address_0_i_7 : std_logic;
signal \this_vga_signals.N_6_0_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c2_0_0_0_1\ : std_logic;
signal \this_vga_signals.g3_3_0\ : std_logic;
signal \this_vga_signals.g3_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_i_cascade_\ : std_logic;
signal \this_vga_signals.g1_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_1\ : std_logic;
signal \this_vga_signals.N_4_i_0_x\ : std_logic;
signal \this_vga_signals.N_4_i_0_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m10_0_x2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m2_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc1\ : std_logic;
signal \this_vga_signals.if_m10_0_a4_1_0_x1\ : std_logic;
signal \this_vga_signals.if_m10_0_a4_1_0_x0_cascade_\ : std_logic;
signal \this_vga_signals.if_m10_0_a4_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c2_0\ : std_logic;
signal \this_vga_signals.g0_0_a3_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNISGOSZ0Z_4_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_1_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_1_x1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_c\ : std_logic;
signal \N_475_cascade_\ : std_logic;
signal \this_vga_signals.if_N_3_mux_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axb2_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_x1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axb2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_x0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_ns\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_1_0_x1\ : std_logic;
signal \this_vga_signals_M_vcounter_q_fast_6\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_1_0_x0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb2_i\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \this_vga_signals.if_m5_0_1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41Z0Z_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_axb1_i_cascade_\ : std_logic;
signal \this_vga_signals.N_81_0\ : std_logic;
signal \this_vga_signals.N_370_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum1_2\ : std_logic;
signal \this_vga_signals_M_vcounter_q_7_rep1\ : std_logic;
signal \this_vga_signals_M_vcounter_q_8_rep1\ : std_logic;
signal \this_vga_signals.N_330_0\ : std_logic;
signal \this_vga_signals.vsync_1_0_a2_6_a2_0\ : std_logic;
signal \this_vga_signals.if_m11_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_i_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_2_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_1_0_x1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_2_2_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_2_2_1_cascade_\ : std_logic;
signal this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0 : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_ns_2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_sx\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_2_4_tz\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_ns_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_2_cascade_\ : std_logic;
signal this_vga_signals_un4_lcounter_if_i3_mux : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_2\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_i\ : std_logic;
signal \this_vga_signals.g0_16_x1\ : std_logic;
signal \this_vga_signals.N_81_1\ : std_logic;
signal \this_vga_signals.g1_2\ : std_logic;
signal \this_vga_signals.if_N_7_i\ : std_logic;
signal \this_vga_signals.if_N_11\ : std_logic;
signal \this_vga_signals.if_i3_mux_0_1_cascade_\ : std_logic;
signal \this_vga_signals.m48_i_x4_3\ : std_logic;
signal \this_vga_signals.if_i3_mux_0_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_0_0\ : std_logic;
signal \this_vga_signals.N_57_0\ : std_logic;
signal \this_vga_signals.N_57_i_i_0\ : std_logic;
signal \this_vga_signals.g1_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_6_mux_0_0_0\ : std_logic;
signal \this_vga_signals.g2_1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0\ : std_logic;
signal \this_vga_signals.N_5_i_1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i\ : std_logic;
signal \this_vga_signals.g0_10_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.if_N_18_1\ : std_logic;
signal \this_vga_signals.m48_i_x4_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_0\ : std_logic;
signal \this_vga_signals.g4_1_0\ : std_logic;
signal \this_vga_signals.g0_1\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_cry_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_cry_1_s\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_cry_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb_3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_cry_2\ : std_logic;
signal \this_vga_signals.vaddress_8\ : std_logic;
signal \this_vga_signals.N_3_2\ : std_logic;
signal \this_vga_signals.g1_4\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_s_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_i_3\ : std_logic;
signal \this_vga_signals.if_N_3_mux\ : std_logic;
signal \this_vga_signals.g6_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0\ : std_logic;
signal \M_this_vga_signals_address_13\ : std_logic;
signal \this_vga_signals.g0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0ASZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_9_repZ0Z1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\ : std_logic;
signal \this_vga_signals.vaddress_7\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.vaddress_6\ : std_logic;
signal \this_vga_signals.N_188_0\ : std_logic;
signal \this_vga_signals.M_this_vga_ramdac_en_i_o2_0_0\ : std_logic;
signal \this_vga_signals.M_this_vga_ramdac_en_i_o2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.N_188_0_0_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_1_0_3\ : std_logic;
signal \this_vga_signals.N_188_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_1_0_2_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_1\ : std_logic;
signal \N_183_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_5_repZ0Z1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_axb1_i\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axb1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_x0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_x1_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_ns_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_ns_1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_repZ0Z1\ : std_logic;
signal \this_vga_signals.if_N_8_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_i_0\ : std_logic;
signal \N_31\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals_M_vcounter_q_6\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.N_177_0_cascade_\ : std_logic;
signal \this_vga_signals.CO0_i_0\ : std_logic;
signal \this_vga_signals.N_269_0\ : std_logic;
signal \this_vga_signals.N_286\ : std_logic;
signal \this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1_cascade_\ : std_logic;
signal \M_this_delay_clk_out_0\ : std_logic;
signal port_enb_c : std_logic;
signal \this_start_data_delay_M_last_q\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_i_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1_0\ : std_logic;
signal \N_90_0\ : std_logic;
signal \this_vga_signals_M_vcounter_q_2\ : std_logic;
signal \this_vga_signals_M_vcounter_q_3\ : std_logic;
signal \N_184_0\ : std_logic;
signal \this_vga_signals_M_vcounter_q_1\ : std_logic;
signal \N_184_0_cascade_\ : std_logic;
signal \this_vga_signals_M_vcounter_q_0\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \G_504\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_cry_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_cry_1_s\ : std_logic;
signal \G_503\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_cry_1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb_3\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_cry_2\ : std_logic;
signal \this_ppu.M_m12_0_o2_381Z0Z_4_cascade_\ : std_logic;
signal \N_275\ : std_logic;
signal \this_ppu.M_m12_0_o2_381_5_cascade_\ : std_logic;
signal \N_190_0\ : std_logic;
signal \this_ppu.M_m12_0_o2_381_8\ : std_logic;
signal \this_vga_signals.N_336_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.N_287\ : std_logic;
signal \this_vga_signals.N_287_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_2_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_\ : std_logic;
signal \this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_1_cascade_\ : std_logic;
signal \this_vga_signals.SUM_7_i_1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_x1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_2\ : std_logic;
signal \this_vga_signals.N_336_0\ : std_logic;
signal \this_vga_signals.N_3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_s_3\ : std_logic;
signal \M_this_vga_signals_pixel_clk_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\ : std_logic;
signal \this_vga_signals.N_517_1_g\ : std_logic;
signal \this_vga_signals.N_684_g\ : std_logic;
signal \this_vga_signals.N_272_0\ : std_logic;
signal \this_vga_signals_M_vcounter_q_4\ : std_logic;
signal \N_475\ : std_logic;
signal \this_vga_signals_M_vcounter_q_5\ : std_logic;
signal \this_vga_signals.N_404_0\ : std_logic;
signal \N_204_0\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_1_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_1_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_1_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_1_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_1_cry_5\ : std_logic;
signal \this_vga_signals_M_hcounter_q_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_1_cry_6\ : std_logic;
signal \this_vga_signals_M_hcounter_q_8\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_1_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_1_cry_8\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \this_vga_signals_M_hcounter_q_9\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUFZ0\ : std_logic;
signal \this_vga_signals_M_hcounter_q_6\ : std_logic;
signal \this_vga_signals.N_517_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc1\ : std_logic;
signal \this_ppu.sprites_addr_1_i_2_1Z0Z_9\ : std_logic;
signal \this_ppu.sprites_addr_1_i_0_0Z0Z_9_cascade_\ : std_logic;
signal \this_ppu.sprites_addr_1_i_a0_2Z0Z_9\ : std_logic;
signal \this_ppu.sprites_addr_1_i_0_2Z0Z_9_cascade_\ : std_logic;
signal \N_138_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_0_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_x0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_x1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_1\ : std_logic;
signal \if_generate_plus_mult1_un68_sum_axbxc3_ns_cascade_\ : std_logic;
signal \this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_cascade_\ : std_logic;
signal \this_vga_signals_M_hcounter_q_5\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_0\ : std_logic;
signal \this_vga_signals_M_hcounter_q_4\ : std_logic;
signal \this_vga_signals.if_N_8_i_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_1\ : std_logic;
signal \M_counter_q_RNIFKS8_0\ : std_logic;
signal \M_counter_q_RNIFKS8_0_cascade_\ : std_logic;
signal \this_pixel_clk_M_counter_q_i_1\ : std_logic;
signal \this_vga_signals.N_455\ : std_logic;
signal \this_vga_signals.N_459\ : std_logic;
signal \this_vga_signals.GZ0Z_210_cascade_\ : std_logic;
signal \this_vga_signals_M_vcounter_q_9\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNIIRV75Z0Z_9\ : std_logic;
signal \this_pixel_clk.M_counter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0\ : std_logic;
signal \if_generate_plus_mult1_un75_sum_axbxc3_cascade_\ : std_logic;
signal \this_ppu.un5_sprites_addr_1_c2_cascade_\ : std_logic;
signal \this_ppu.N_4_0_1\ : std_logic;
signal \this_ppu.sprites_addr_1_i_7_tz_0_9\ : std_logic;
signal \this_ppu.sprites_addr_1_i_a7Z0Z_9\ : std_logic;
signal this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3 : std_logic;
signal \this_ppu.un5_sprites_addr1_4\ : std_logic;
signal this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_c3 : std_logic;
signal this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0 : std_logic;
signal \this_vga_signals.GZ0Z_210\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI4UBI1Z0Z_9\ : std_logic;
signal \this_vga_signals_M_hcounter_q_3\ : std_logic;
signal \this_vga_signals.if_N_9_1\ : std_logic;
signal \this_ppu.sprites_m1_0_xZ0Z1\ : std_logic;
signal \this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3_cascade_\ : std_logic;
signal \this_ppu.sprites_m1_0_xZ0Z0\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_2\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_9\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_3_cascade_\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_8\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \un1_M_this_data_count_q_cry_0\ : std_logic;
signal \un1_M_this_data_count_q_cry_1\ : std_logic;
signal \un1_M_this_data_count_q_cry_2\ : std_logic;
signal \un1_M_this_data_count_q_cry_3\ : std_logic;
signal \un1_M_this_data_count_q_cry_4\ : std_logic;
signal \un1_M_this_data_count_q_cry_5\ : std_logic;
signal \un1_M_this_data_count_q_cry_6\ : std_logic;
signal \un1_M_this_data_count_q_cry_7\ : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal \un1_M_this_data_count_q_cry_8\ : std_logic;
signal \un1_M_this_data_count_q_cry_9\ : std_logic;
signal \un1_M_this_data_count_q_cry_10\ : std_logic;
signal \un1_M_this_data_count_q_cry_11\ : std_logic;
signal \M_this_state_q_RNI20CEZ0Z_0\ : std_logic;
signal \un1_M_this_data_count_q_cry_12\ : std_logic;
signal \un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO\ : std_logic;
signal \un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO\ : std_logic;
signal \bfn_15_25_0_\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \N_13_0\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \this_ppu.un5_sprites_addr_1_c4\ : std_logic;
signal \this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_c3_0_cascade_\ : std_logic;
signal if_generate_plus_mult1_un89_sum_axbxc3 : std_logic;
signal \this_ppu.sprites_N_7_0_cascade_\ : std_logic;
signal \this_ppu.un5_sprites_addr_1_c2\ : std_logic;
signal \this_ppu.sprites_m7Z0Z_0_cascade_\ : std_logic;
signal if_generate_plus_mult1_un68_sum_axbxc3_ns : std_logic;
signal \N_140_i\ : std_logic;
signal \this_vga_signals_M_hcounter_q_2\ : std_logic;
signal this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1 : std_logic;
signal this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3 : std_logic;
signal if_generate_plus_mult1_un75_sum_axbxc3 : std_logic;
signal this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0 : std_logic;
signal \this_vga_signals_M_hcounter_q_1\ : std_logic;
signal \this_vga_signals_M_hcounter_q_0\ : std_logic;
signal \this_ppu.sprites_mZ0Z1_cascade_\ : std_logic;
signal this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axb1 : std_logic;
signal \M_this_internal_address_q_3_ns_1_10_cascade_\ : std_logic;
signal \bfn_16_21_0_\ : std_logic;
signal \un1_M_this_internal_address_q_cry_0\ : std_logic;
signal \M_this_internal_address_qZ0Z_2\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_2\ : std_logic;
signal \un1_M_this_internal_address_q_cry_1\ : std_logic;
signal \M_this_internal_address_qZ0Z_3\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_3\ : std_logic;
signal \un1_M_this_internal_address_q_cry_2\ : std_logic;
signal \un1_M_this_internal_address_q_cry_3\ : std_logic;
signal \un1_M_this_internal_address_q_cry_4\ : std_logic;
signal \un1_M_this_internal_address_q_cry_5\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_7\ : std_logic;
signal \un1_M_this_internal_address_q_cry_6\ : std_logic;
signal \un1_M_this_internal_address_q_cry_7\ : std_logic;
signal \M_this_internal_address_qZ0Z_8\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_8\ : std_logic;
signal \bfn_16_22_0_\ : std_logic;
signal \M_this_internal_address_qZ0Z_9\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_9\ : std_logic;
signal \un1_M_this_internal_address_q_cry_8\ : std_logic;
signal \M_this_internal_address_qZ0Z_10\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_10\ : std_logic;
signal \un1_M_this_internal_address_q_cry_9\ : std_logic;
signal \un1_M_this_internal_address_q_cry_10\ : std_logic;
signal \un1_M_this_internal_address_q_cry_11\ : std_logic;
signal \un1_M_this_internal_address_q_cry_12\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_13\ : std_logic;
signal \M_this_internal_address_qZ0Z_7\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_7\ : std_logic;
signal \N_235_0_i\ : std_logic;
signal \M_this_data_count_qZ0Z_13\ : std_logic;
signal \M_this_data_count_qZ0Z_0\ : std_logic;
signal \M_this_data_count_qZ0Z_11\ : std_logic;
signal \M_this_data_count_qZ0Z_9\ : std_logic;
signal \M_this_data_count_qZ0Z_8\ : std_logic;
signal \M_this_data_count_qZ0Z_12\ : std_logic;
signal \M_this_data_count_qZ0Z_6\ : std_logic;
signal \M_this_data_count_qZ0Z_5\ : std_logic;
signal \M_this_data_count_qZ0Z_7\ : std_logic;
signal \M_this_data_count_qZ0Z_4\ : std_logic;
signal \M_this_data_count_qZ0Z_3\ : std_logic;
signal \M_this_data_count_qZ0Z_2\ : std_logic;
signal \M_this_data_count_qZ0Z_10\ : std_logic;
signal \M_this_data_count_qZ0Z_1\ : std_logic;
signal \M_this_state_q_srsts_0_a2_1_9_4\ : std_logic;
signal \M_this_state_q_srsts_0_a2_1_7_4\ : std_logic;
signal \M_this_state_q_srsts_0_a2_1_8_4_cascade_\ : std_logic;
signal \M_this_state_q_srsts_0_a2_1_6_4\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_c3_0 : std_logic;
signal \this_ppu_sprites_N_2_1\ : std_logic;
signal \N_134_0\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_4\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_4_cascade_\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_i_1Z0Z_4\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_i_0Z0Z_4\ : std_logic;
signal \this_vga_signals.N_224_0\ : std_logic;
signal \M_this_state_q_nss_0\ : std_logic;
signal \N_235_0\ : std_logic;
signal \this_vga_signals.N_319\ : std_logic;
signal un19_i_i_i_a2 : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_11\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_0\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_0\ : std_logic;
signal \M_this_internal_address_qZ0Z_0\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_1\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_1\ : std_logic;
signal \M_this_internal_address_qZ0Z_1\ : std_logic;
signal \N_476\ : std_logic;
signal \N_240\ : std_logic;
signal \M_this_state_qZ0Z_1\ : std_logic;
signal \this_vga_signals.N_343_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_2\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_5\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_6\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_12\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_11\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_4\ : std_logic;
signal \M_this_internal_address_q_RNO_1Z0Z_4\ : std_logic;
signal \M_this_internal_address_qZ0Z_4\ : std_logic;
signal \M_this_vram_write_data_1\ : std_logic;
signal port_address_in_7 : std_logic;
signal port_address_in_6 : std_logic;
signal port_rw_in : std_logic;
signal \this_vga_signals.N_185_0\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_i_o4_4Z0Z_4\ : std_logic;
signal \M_this_state_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_i_o4_4Z0Z_4_cascade_\ : std_logic;
signal \this_vga_signals.N_490_cascade_\ : std_logic;
signal \this_vga_signals.N_386_cascade_\ : std_logic;
signal \this_vga_signals.N_387_cascade_\ : std_logic;
signal port_address_in_1 : std_logic;
signal port_address_in_0 : std_logic;
signal \this_vga_signals.N_391_cascade_\ : std_logic;
signal \this_vga_signals.N_490\ : std_logic;
signal \M_this_state_qZ0Z_5\ : std_logic;
signal \M_this_state_qZ0Z_6\ : std_logic;
signal \N_14_0\ : std_logic;
signal \M_this_internal_address_qZ0Z_5\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_5\ : std_logic;
signal \M_this_internal_address_qZ0Z_6\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_6\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_13\ : std_logic;
signal \N_355\ : std_logic;
signal \M_this_internal_address_q_3_ns_1_12\ : std_logic;
signal \M_this_state_qZ0Z_7\ : std_logic;
signal port_data_c_5 : std_logic;
signal port_data_c_1 : std_logic;
signal \M_this_sprites_ram_write_data_1\ : std_logic;
signal port_data_c_0 : std_logic;
signal port_data_c_4 : std_logic;
signal \M_this_sprites_ram_write_data_0\ : std_logic;
signal \M_this_vram_write_data_2\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_2\ : std_logic;
signal \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\ : std_logic;
signal \M_this_sprites_ram_read_data_2\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\ : std_logic;
signal \M_this_sprites_ram_read_data_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_1\ : std_logic;
signal \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_0\ : std_logic;
signal \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0\ : std_logic;
signal \M_this_sprites_ram_read_data_3_cascade_\ : std_logic;
signal \M_this_ppu_vram_en_0\ : std_logic;
signal \M_this_vram_write_data_3\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_11\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_12\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_0\ : std_logic;
signal \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_0\ : std_logic;
signal \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\ : std_logic;
signal \this_vga_signals.N_483\ : std_logic;
signal \N_175_0\ : std_logic;
signal \this_sprites_ram.mem_WE_0\ : std_logic;
signal \this_sprites_ram.mem_WE_14\ : std_logic;
signal \this_sprites_ram.mem_WE_10\ : std_logic;
signal \this_sprites_ram.mem_WE_12\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_2\ : std_logic;
signal \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_1\ : std_logic;
signal \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_2\ : std_logic;
signal \this_sprites_ram.mem_mem_0_1_RNIL62PZ0\ : std_logic;
signal \this_sprites_ram.mem_WE_8\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_2\ : std_logic;
signal \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_1\ : std_logic;
signal \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_1\ : std_logic;
signal \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_3\ : std_logic;
signal \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_WE_6\ : std_logic;
signal port_data_c_3 : std_logic;
signal port_data_c_7 : std_logic;
signal \M_this_sprites_ram_write_data_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_3\ : std_logic;
signal \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_3\ : std_logic;
signal \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_3\ : std_logic;
signal \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_0\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_13\ : std_logic;
signal \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\ : std_logic;
signal \this_vga_signals.N_481\ : std_logic;
signal port_data_c_2 : std_logic;
signal port_data_c_6 : std_logic;
signal \this_vga_signals.N_479\ : std_logic;
signal \M_this_sprites_ram_write_data_2\ : std_logic;
signal \this_sprites_ram.mem_WE_4\ : std_logic;
signal \M_this_internal_address_qZ0Z_12\ : std_logic;
signal \M_this_internal_address_qZ0Z_11\ : std_logic;
signal \M_this_internal_address_qZ0Z_13\ : std_logic;
signal \N_24_0\ : std_logic;
signal \this_sprites_ram.mem_WE_2\ : std_logic;
signal \N_192_0\ : std_logic;
signal this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2 : std_logic;
signal \this_ppu.sprites_N_6\ : std_logic;
signal sprites_m7 : std_logic;
signal \M_this_state_qZ0Z_3\ : std_logic;
signal \M_this_external_address_qZ0Z_0\ : std_logic;
signal \bfn_31_23_0_\ : std_logic;
signal \M_this_external_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_external_address_q_cry_0\ : std_logic;
signal \M_this_external_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_external_address_q_cry_1\ : std_logic;
signal \M_this_external_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_external_address_q_cry_2\ : std_logic;
signal \M_this_external_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_external_address_q_cry_3\ : std_logic;
signal \M_this_external_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_external_address_q_cry_4\ : std_logic;
signal \M_this_external_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_external_address_q_cry_5\ : std_logic;
signal \M_this_external_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_external_address_q_cry_6\ : std_logic;
signal \un1_M_this_external_address_q_cry_7\ : std_logic;
signal \M_this_external_address_qZ0Z_8\ : std_logic;
signal \bfn_31_24_0_\ : std_logic;
signal \M_this_external_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_external_address_q_cry_8\ : std_logic;
signal \M_this_external_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_external_address_q_cry_9\ : std_logic;
signal \M_this_external_address_qZ0Z_11\ : std_logic;
signal \un1_M_this_external_address_q_cry_10\ : std_logic;
signal \M_this_external_address_qZ0Z_12\ : std_logic;
signal \un1_M_this_external_address_q_cry_11\ : std_logic;
signal \M_this_external_address_qZ0Z_13\ : std_logic;
signal \un1_M_this_external_address_q_cry_12\ : std_logic;
signal \M_this_external_address_qZ0Z_14\ : std_logic;
signal \un1_M_this_external_address_q_cry_13\ : std_logic;
signal \M_this_state_qZ0Z_0\ : std_logic;
signal \un1_M_this_external_address_q_cry_14\ : std_logic;
signal \M_this_external_address_qZ0Z_15\ : std_logic;
signal clk_0_c_g : std_logic;
signal \M_this_state_q_nss_g_0\ : std_logic;
signal port_address_in_2 : std_logic;
signal port_address_in_3 : std_logic;
signal port_address_in_4 : std_logic;
signal port_address_in_5 : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_i_o4_5Z0Z_4\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic_vector(1 downto 0);
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \this_sprites_ram.mem_out_bus0_1\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_0\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ <= \N__18215\&\N__16481\&\N__23654\&\N__19736\&\N__10196\&\N__10478\&\N__10340\&\N__10970\&\N__10049\&\N__10835\&\N__11111\;
    \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ <= \N__19058\&\N__19187\&\N__19313\&\N__18899\&\N__21374\&\N__21506\&\N__20366\&\N__18443\&\N__18575\&\N__19964\&\N__20105\;
    \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20966\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20789\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus0_3\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_2\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ <= \N__18209\&\N__16475\&\N__23648\&\N__19730\&\N__10190\&\N__10472\&\N__10334\&\N__10964\&\N__10043\&\N__10829\&\N__11105\;
    \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ <= \N__19052\&\N__19181\&\N__19307\&\N__18893\&\N__21368\&\N__21500\&\N__20360\&\N__18437\&\N__18569\&\N__19958\&\N__20099\;
    \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__23107\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24314\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_1\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_0\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ <= \N__18203\&\N__16469\&\N__23642\&\N__19724\&\N__10184\&\N__10466\&\N__10328\&\N__10958\&\N__10037\&\N__10823\&\N__11099\;
    \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ <= \N__19046\&\N__19175\&\N__19301\&\N__18887\&\N__21362\&\N__21494\&\N__20354\&\N__18431\&\N__18563\&\N__19952\&\N__20093\;
    \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20972\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20785\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_3\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_2\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ <= \N__18197\&\N__16463\&\N__23636\&\N__19718\&\N__10178\&\N__10460\&\N__10322\&\N__10952\&\N__10031\&\N__10817\&\N__11093\;
    \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ <= \N__19040\&\N__19169\&\N__19295\&\N__18881\&\N__21356\&\N__21488\&\N__20348\&\N__18425\&\N__18557\&\N__19946\&\N__20087\;
    \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__23099\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24310\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_1\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_0\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ <= \N__18191\&\N__16457\&\N__23630\&\N__19712\&\N__10172\&\N__10454\&\N__10316\&\N__10946\&\N__10025\&\N__10811\&\N__11087\;
    \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ <= \N__19034\&\N__19163\&\N__19289\&\N__18875\&\N__21350\&\N__21482\&\N__20342\&\N__18419\&\N__18551\&\N__19940\&\N__20081\;
    \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20968\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20778\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_3\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_2\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ <= \N__18185\&\N__16451\&\N__23624\&\N__19706\&\N__10166\&\N__10448\&\N__10310\&\N__10940\&\N__10019\&\N__10805\&\N__11081\;
    \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ <= \N__19028\&\N__19157\&\N__19283\&\N__18869\&\N__21344\&\N__21476\&\N__20336\&\N__18413\&\N__18545\&\N__19934\&\N__20075\;
    \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__23085\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24302\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_1\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_0\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ <= \N__18179\&\N__16445\&\N__23618\&\N__19700\&\N__10160\&\N__10442\&\N__10304\&\N__10934\&\N__10013\&\N__10799\&\N__11075\;
    \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ <= \N__19022\&\N__19151\&\N__19277\&\N__18863\&\N__21338\&\N__21470\&\N__20330\&\N__18407\&\N__18539\&\N__19928\&\N__20069\;
    \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20952\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20767\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_3\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_2\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ <= \N__18173\&\N__16439\&\N__23612\&\N__19694\&\N__10154\&\N__10436\&\N__10298\&\N__10928\&\N__10007\&\N__10793\&\N__11069\;
    \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ <= \N__19016\&\N__19145\&\N__19271\&\N__18857\&\N__21332\&\N__21464\&\N__20324\&\N__18401\&\N__18533\&\N__19922\&\N__20063\;
    \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__23067\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24288\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_1\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_0\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ <= \N__18167\&\N__16433\&\N__23606\&\N__19688\&\N__10148\&\N__10430\&\N__10292\&\N__10922\&\N__10001\&\N__10787\&\N__11063\;
    \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ <= \N__19010\&\N__19139\&\N__19265\&\N__18851\&\N__21326\&\N__21458\&\N__20318\&\N__18395\&\N__18527\&\N__19916\&\N__20057\;
    \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20938\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20745\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_3\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_2\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ <= \N__18161\&\N__16427\&\N__23600\&\N__19682\&\N__10142\&\N__10424\&\N__10286\&\N__10916\&\N__9995\&\N__10781\&\N__11057\;
    \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ <= \N__19004\&\N__19133\&\N__19259\&\N__18845\&\N__21320\&\N__21452\&\N__20312\&\N__18389\&\N__18521\&\N__19910\&\N__20051\;
    \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__23076\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24248\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_1\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_0\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ <= \N__18155\&\N__16421\&\N__23594\&\N__19676\&\N__10136\&\N__10418\&\N__10280\&\N__10910\&\N__9989\&\N__10775\&\N__11051\;
    \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ <= \N__18998\&\N__19127\&\N__19253\&\N__18839\&\N__21314\&\N__21446\&\N__20306\&\N__18383\&\N__18515\&\N__19904\&\N__20045\;
    \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20939\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20744\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_3\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_2\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ <= \N__18149\&\N__16415\&\N__23588\&\N__19670\&\N__10130\&\N__10412\&\N__10274\&\N__10904\&\N__9983\&\N__10769\&\N__11045\;
    \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ <= \N__18992\&\N__19121\&\N__19247\&\N__18833\&\N__21308\&\N__21440\&\N__20300\&\N__18377\&\N__18509\&\N__19898\&\N__20039\;
    \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__23092\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24281\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_1\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_0\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ <= \N__18143\&\N__16409\&\N__23582\&\N__19664\&\N__10124\&\N__10406\&\N__10268\&\N__10898\&\N__9977\&\N__10763\&\N__11039\;
    \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ <= \N__18986\&\N__19115\&\N__19241\&\N__18827\&\N__21302\&\N__21434\&\N__20294\&\N__18371\&\N__18503\&\N__19892\&\N__20033\;
    \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20956\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20763\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_3\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_2\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ <= \N__18137\&\N__16403\&\N__23576\&\N__19658\&\N__10118\&\N__10400\&\N__10262\&\N__10892\&\N__9971\&\N__10757\&\N__11033\;
    \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ <= \N__18980\&\N__19109\&\N__19235\&\N__18821\&\N__21296\&\N__21428\&\N__20288\&\N__18365\&\N__18497\&\N__19886\&\N__20027\;
    \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__23103\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24298\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_1\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_0\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ <= \N__18131\&\N__16397\&\N__23570\&\N__19652\&\N__10112\&\N__10394\&\N__10256\&\N__10886\&\N__9965\&\N__10751\&\N__11027\;
    \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ <= \N__18974\&\N__19103\&\N__19229\&\N__18815\&\N__21290\&\N__21422\&\N__20282\&\N__18359\&\N__18491\&\N__19880\&\N__20021\;
    \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20967\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20777\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_3\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_2\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ <= \N__18125\&\N__16391\&\N__23564\&\N__19646\&\N__10106\&\N__10388\&\N__10250\&\N__10879\&\N__9959\&\N__10745\&\N__11021\;
    \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ <= \N__18968\&\N__19097\&\N__19223\&\N__18809\&\N__21284\&\N__21416\&\N__20276\&\N__18353\&\N__18485\&\N__19874\&\N__20015\;
    \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__23108\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24309\&'0'&'0'&'0';
    \M_this_vram_read_data_3\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_vram_read_data_2\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_vram_read_data_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_vram_read_data_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__12761\&\N__9050\&\N__9002\&\N__9491\&\N__8987\&\N__9011\&\N__11156\&\N__17309\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__14597\&\N__10099\&\N__10381\&\N__10246\&\N__10882\&\N__9952\&\N__10738\&\N__11017\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22322\&\N__21836\&\N__20240\&\N__10682\;

    \this_sprites_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24961\,
            RE => \N__17674\,
            WCLKE => \N__21866\,
            WCLK => \N__24962\,
            WE => \N__17492\
        );

    \this_sprites_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24963\,
            RE => \N__17673\,
            WCLKE => \N__21865\,
            WCLK => \N__24964\,
            WE => \N__17675\
        );

    \this_sprites_ram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24967\,
            RE => \N__17661\,
            WCLKE => \N__22661\,
            WCLK => \N__24968\,
            WE => \N__17672\
        );

    \this_sprites_ram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24971\,
            RE => \N__17660\,
            WCLKE => \N__22660\,
            WCLK => \N__24972\,
            WE => \N__17671\
        );

    \this_sprites_ram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24980\,
            RE => \N__17637\,
            WCLKE => \N__22676\,
            WCLK => \N__24979\,
            WE => \N__17659\
        );

    \this_sprites_ram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24992\,
            RE => \N__17636\,
            WCLKE => \N__22675\,
            WCLK => \N__24993\,
            WE => \N__17658\
        );

    \this_sprites_ram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__25000\,
            RE => \N__17604\,
            WCLKE => \N__22537\,
            WCLK => \N__25001\,
            WE => \N__17631\
        );

    \this_sprites_ram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__25010\,
            RE => \N__17603\,
            WCLKE => \N__22538\,
            WCLK => \N__25011\,
            WE => \N__17629\
        );

    \this_sprites_ram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__25019\,
            RE => \N__17560\,
            WCLKE => \N__23209\,
            WCLK => \N__25020\,
            WE => \N__17591\
        );

    \this_sprites_ram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__25022\,
            RE => \N__17559\,
            WCLKE => \N__23213\,
            WCLK => \N__25023\,
            WE => \N__17549\
        );

    \this_sprites_ram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__25024\,
            RE => \N__17503\,
            WCLKE => \N__24226\,
            WCLK => \N__25025\,
            WE => \N__17540\
        );

    \this_sprites_ram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__25026\,
            RE => \N__17502\,
            WCLKE => \N__24230\,
            WCLK => \N__25027\,
            WE => \N__17458\
        );

    \this_sprites_ram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__25028\,
            RE => \N__17522\,
            WCLKE => \N__23878\,
            WCLK => \N__25029\,
            WE => \N__17533\
        );

    \this_sprites_ram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__25030\,
            RE => \N__17523\,
            WCLKE => \N__23882\,
            WCLK => \N__25031\,
            WE => \N__17589\
        );

    \this_sprites_ram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__25032\,
            RE => \N__17584\,
            WCLKE => \N__21886\,
            WCLK => \N__25033\,
            WE => \N__17590\
        );

    \this_sprites_ram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__25036\,
            RE => \N__17585\,
            WCLKE => \N__21890\,
            WCLK => \N__25037\,
            WE => \N__17630\
        );

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__24976\,
            RE => \N__17635\,
            WCLKE => \N__9116\,
            WCLK => \N__24975\,
            WE => \N__17598\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__25731\,
            GLOBALBUFFEROUTPUT => clk_0_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25733\,
            DIN => \N__25732\,
            DOUT => \N__25731\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__25733\,
            PADOUT => \N__25732\,
            PADIN => \N__25731\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25722\,
            DIN => \N__25721\,
            DOUT => \N__25720\,
            PACKAGEPIN => debug_wire(0)
        );

    \debug_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__25722\,
            PADOUT => \N__25721\,
            PADIN => \N__25720\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25713\,
            DIN => \N__25712\,
            DOUT => \N__25711\,
            PACKAGEPIN => debug_wire(1)
        );

    \debug_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__25713\,
            PADOUT => \N__25712\,
            PADIN => \N__25711\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25704\,
            DIN => \N__25703\,
            DOUT => \N__25702\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__25704\,
            PADOUT => \N__25703\,
            PADIN => \N__25702\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__9464\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25695\,
            DIN => \N__25694\,
            DOUT => \N__25693\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__25695\,
            PADOUT => \N__25694\,
            PADIN => \N__25693\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13829\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25686\,
            DIN => \N__25685\,
            DOUT => \N__25684\,
            PACKAGEPIN => port_address(0)
        );

    \port_address_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25686\,
            PADOUT => \N__25685\,
            PADIN => \N__25684\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__23363\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18673\
        );

    \port_address_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25677\,
            DIN => \N__25676\,
            DOUT => \N__25675\,
            PACKAGEPIN => port_address(1)
        );

    \port_address_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25677\,
            PADOUT => \N__25676\,
            PADIN => \N__25675\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__23336\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18749\
        );

    \port_address_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25668\,
            DIN => \N__25667\,
            DOUT => \N__25666\,
            PACKAGEPIN => port_address(2)
        );

    \port_address_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25668\,
            PADOUT => \N__25667\,
            PADIN => \N__25666\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__23315\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18729\
        );

    \port_address_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25659\,
            DIN => \N__25658\,
            DOUT => \N__25657\,
            PACKAGEPIN => port_address(3)
        );

    \port_address_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25659\,
            PADOUT => \N__25658\,
            PADIN => \N__25657\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__23285\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18758\
        );

    \port_address_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25650\,
            DIN => \N__25649\,
            DOUT => \N__25648\,
            PACKAGEPIN => port_address(4)
        );

    \port_address_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25650\,
            PADOUT => \N__25649\,
            PADIN => \N__25648\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__23261\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18642\
        );

    \port_address_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25641\,
            DIN => \N__25640\,
            DOUT => \N__25639\,
            PACKAGEPIN => port_address(5)
        );

    \port_address_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25641\,
            PADOUT => \N__25640\,
            PADIN => \N__25639\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__24563\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18715\
        );

    \port_address_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25632\,
            DIN => \N__25631\,
            DOUT => \N__25630\,
            PACKAGEPIN => port_address(6)
        );

    \port_address_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25632\,
            PADOUT => \N__25631\,
            PADIN => \N__25630\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__24542\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18740\
        );

    \port_address_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25623\,
            DIN => \N__25622\,
            DOUT => \N__25621\,
            PACKAGEPIN => port_address(7)
        );

    \port_address_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25623\,
            PADOUT => \N__25622\,
            PADIN => \N__25621\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__24521\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18767\
        );

    \port_address_obuft_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25614\,
            DIN => \N__25613\,
            DOUT => \N__25612\,
            PACKAGEPIN => port_address(10)
        );

    \port_address_obuft_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25614\,
            PADOUT => \N__25613\,
            PADIN => \N__25612\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__24434\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18653\
        );

    \port_address_obuft_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25605\,
            DIN => \N__25604\,
            DOUT => \N__25603\,
            PACKAGEPIN => port_address(11)
        );

    \port_address_obuft_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25605\,
            PADOUT => \N__25604\,
            PADIN => \N__25603\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__24404\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18759\
        );

    \port_address_obuft_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25596\,
            DIN => \N__25595\,
            DOUT => \N__25594\,
            PACKAGEPIN => port_address(12)
        );

    \port_address_obuft_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25596\,
            PADOUT => \N__25595\,
            PADIN => \N__25594\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__24377\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18714\
        );

    \port_address_obuft_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25587\,
            DIN => \N__25586\,
            DOUT => \N__25585\,
            PACKAGEPIN => port_address(13)
        );

    \port_address_obuft_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25587\,
            PADOUT => \N__25586\,
            PADIN => \N__25585\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__25325\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18716\
        );

    \port_address_obuft_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25578\,
            DIN => \N__25577\,
            DOUT => \N__25576\,
            PACKAGEPIN => port_address(14)
        );

    \port_address_obuft_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25578\,
            PADOUT => \N__25577\,
            PADIN => \N__25576\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__25301\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18741\
        );

    \port_address_obuft_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25569\,
            DIN => \N__25568\,
            DOUT => \N__25567\,
            PACKAGEPIN => port_address(15)
        );

    \port_address_obuft_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25569\,
            PADOUT => \N__25568\,
            PADIN => \N__25567\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__25061\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18766\
        );

    \port_address_obuft_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25560\,
            DIN => \N__25559\,
            DOUT => \N__25558\,
            PACKAGEPIN => port_address(8)
        );

    \port_address_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25560\,
            PADOUT => \N__25559\,
            PADIN => \N__25558\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__24494\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18638\
        );

    \port_address_obuft_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25551\,
            DIN => \N__25550\,
            DOUT => \N__25549\,
            PACKAGEPIN => port_address(9)
        );

    \port_address_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25551\,
            PADOUT => \N__25550\,
            PADIN => \N__25549\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__24464\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18748\
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25542\,
            DIN => \N__25541\,
            DOUT => \N__25540\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__25542\,
            PADOUT => \N__25541\,
            PADIN => \N__25540\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25533\,
            DIN => \N__25532\,
            DOUT => \N__25531\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__25533\,
            PADOUT => \N__25532\,
            PADIN => \N__25531\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25524\,
            DIN => \N__25523\,
            DOUT => \N__25522\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__25524\,
            PADOUT => \N__25523\,
            PADIN => \N__25522\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25515\,
            DIN => \N__25514\,
            DOUT => \N__25513\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__25515\,
            PADOUT => \N__25514\,
            PADIN => \N__25513\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25506\,
            DIN => \N__25505\,
            DOUT => \N__25504\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__25506\,
            PADOUT => \N__25505\,
            PADIN => \N__25504\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25497\,
            DIN => \N__25496\,
            DOUT => \N__25495\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__25497\,
            PADOUT => \N__25496\,
            PADIN => \N__25495\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25488\,
            DIN => \N__25487\,
            DOUT => \N__25486\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__25488\,
            PADOUT => \N__25487\,
            PADIN => \N__25486\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25479\,
            DIN => \N__25478\,
            DOUT => \N__25477\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__25479\,
            PADOUT => \N__25478\,
            PADIN => \N__25477\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25470\,
            DIN => \N__25469\,
            DOUT => \N__25468\,
            PACKAGEPIN => port_data_wire(7)
        );

    \port_data_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__25470\,
            PADOUT => \N__25469\,
            PADIN => \N__25468\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25461\,
            DIN => \N__25460\,
            DOUT => \N__25459\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__25461\,
            PADOUT => \N__25460\,
            PADIN => \N__25459\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8609\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25452\,
            DIN => \N__25451\,
            DOUT => \N__25450\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__25452\,
            PADOUT => \N__25451\,
            PADIN => \N__25450\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__20222\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25443\,
            DIN => \N__25442\,
            DOUT => \N__25441\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__25443\,
            PADOUT => \N__25442\,
            PADIN => \N__25441\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25434\,
            DIN => \N__25433\,
            DOUT => \N__25432\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__25434\,
            PADOUT => \N__25433\,
            PADIN => \N__25432\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8651\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25425\,
            DIN => \N__25424\,
            DOUT => \N__25423\,
            PACKAGEPIN => port_rw
        );

    \port_rw_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__25425\,
            PADOUT => \N__25424\,
            PADIN => \N__25423\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_in,
            DIN1 => OPEN,
            DOUT0 => \N__17602\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18739\
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25416\,
            DIN => \N__25415\,
            DOUT => \N__25414\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__25416\,
            PADOUT => \N__25415\,
            PADIN => \N__25414\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8603\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__15620\,
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25407\,
            DIN => \N__25406\,
            DOUT => \N__25405\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__25407\,
            PADOUT => \N__25406\,
            PADIN => \N__25405\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8585\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__15609\,
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25398\,
            DIN => \N__25397\,
            DOUT => \N__25396\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__25398\,
            PADOUT => \N__25397\,
            PADIN => \N__25396\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8927\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__15613\,
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25389\,
            DIN => \N__25388\,
            DOUT => \N__25387\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__25389\,
            PADOUT => \N__25388\,
            PADIN => \N__25387\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8969\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__15622\,
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25380\,
            DIN => \N__25379\,
            DOUT => \N__25378\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__25380\,
            PADOUT => \N__25379\,
            PADIN => \N__25378\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8945\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__15621\,
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25371\,
            DIN => \N__25370\,
            DOUT => \N__25369\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "010101"
        )
    port map (
            PADOEN => \N__25371\,
            PADOUT => \N__25370\,
            PADIN => \N__25369\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8672\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => \N__15623\,
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25362\,
            DIN => \N__25361\,
            DOUT => \N__25360\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__25362\,
            PADOUT => \N__25361\,
            PADIN => \N__25360\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25353\,
            DIN => \N__25352\,
            DOUT => \N__25351\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__25353\,
            PADOUT => \N__25352\,
            PADIN => \N__25351\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8636\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25344\,
            DIN => \N__25343\,
            DOUT => \N__25342\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__25344\,
            PADOUT => \N__25343\,
            PADIN => \N__25342\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__10646\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__6214\ : IoInMux
    port map (
            O => \N__25325\,
            I => \N__25322\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__25322\,
            I => \N__25319\
        );

    \I__6212\ : IoSpan4Mux
    port map (
            O => \N__25319\,
            I => \N__25316\
        );

    \I__6211\ : Span4Mux_s1_h
    port map (
            O => \N__25316\,
            I => \N__25312\
        );

    \I__6210\ : InMux
    port map (
            O => \N__25315\,
            I => \N__25309\
        );

    \I__6209\ : Odrv4
    port map (
            O => \N__25312\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__25309\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__6207\ : InMux
    port map (
            O => \N__25304\,
            I => \un1_M_this_external_address_q_cry_12\
        );

    \I__6206\ : IoInMux
    port map (
            O => \N__25301\,
            I => \N__25298\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__25298\,
            I => \N__25295\
        );

    \I__6204\ : Span4Mux_s1_h
    port map (
            O => \N__25295\,
            I => \N__25292\
        );

    \I__6203\ : Sp12to4
    port map (
            O => \N__25292\,
            I => \N__25288\
        );

    \I__6202\ : InMux
    port map (
            O => \N__25291\,
            I => \N__25285\
        );

    \I__6201\ : Odrv12
    port map (
            O => \N__25288\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__25285\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__6199\ : InMux
    port map (
            O => \N__25280\,
            I => \un1_M_this_external_address_q_cry_13\
        );

    \I__6198\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25265\
        );

    \I__6197\ : InMux
    port map (
            O => \N__25276\,
            I => \N__25265\
        );

    \I__6196\ : InMux
    port map (
            O => \N__25275\,
            I => \N__25265\
        );

    \I__6195\ : InMux
    port map (
            O => \N__25274\,
            I => \N__25265\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__25265\,
            I => \N__25248\
        );

    \I__6193\ : InMux
    port map (
            O => \N__25264\,
            I => \N__25239\
        );

    \I__6192\ : InMux
    port map (
            O => \N__25263\,
            I => \N__25239\
        );

    \I__6191\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25239\
        );

    \I__6190\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25239\
        );

    \I__6189\ : InMux
    port map (
            O => \N__25260\,
            I => \N__25230\
        );

    \I__6188\ : InMux
    port map (
            O => \N__25259\,
            I => \N__25230\
        );

    \I__6187\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25230\
        );

    \I__6186\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25230\
        );

    \I__6185\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25221\
        );

    \I__6184\ : InMux
    port map (
            O => \N__25255\,
            I => \N__25221\
        );

    \I__6183\ : InMux
    port map (
            O => \N__25254\,
            I => \N__25221\
        );

    \I__6182\ : InMux
    port map (
            O => \N__25253\,
            I => \N__25221\
        );

    \I__6181\ : CascadeMux
    port map (
            O => \N__25252\,
            I => \N__25216\
        );

    \I__6180\ : InMux
    port map (
            O => \N__25251\,
            I => \N__25209\
        );

    \I__6179\ : Span4Mux_h
    port map (
            O => \N__25248\,
            I => \N__25204\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__25239\,
            I => \N__25204\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__25230\,
            I => \N__25201\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__25221\,
            I => \N__25198\
        );

    \I__6175\ : InMux
    port map (
            O => \N__25220\,
            I => \N__25193\
        );

    \I__6174\ : InMux
    port map (
            O => \N__25219\,
            I => \N__25190\
        );

    \I__6173\ : InMux
    port map (
            O => \N__25216\,
            I => \N__25187\
        );

    \I__6172\ : InMux
    port map (
            O => \N__25215\,
            I => \N__25182\
        );

    \I__6171\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25182\
        );

    \I__6170\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25179\
        );

    \I__6169\ : InMux
    port map (
            O => \N__25212\,
            I => \N__25176\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__25209\,
            I => \N__25173\
        );

    \I__6167\ : Span4Mux_v
    port map (
            O => \N__25204\,
            I => \N__25170\
        );

    \I__6166\ : Span4Mux_v
    port map (
            O => \N__25201\,
            I => \N__25165\
        );

    \I__6165\ : Span4Mux_v
    port map (
            O => \N__25198\,
            I => \N__25165\
        );

    \I__6164\ : InMux
    port map (
            O => \N__25197\,
            I => \N__25162\
        );

    \I__6163\ : CascadeMux
    port map (
            O => \N__25196\,
            I => \N__25156\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__25193\,
            I => \N__25147\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__25190\,
            I => \N__25147\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__25187\,
            I => \N__25144\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__25182\,
            I => \N__25135\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__25179\,
            I => \N__25135\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__25176\,
            I => \N__25135\
        );

    \I__6156\ : Span4Mux_v
    port map (
            O => \N__25173\,
            I => \N__25135\
        );

    \I__6155\ : Span4Mux_h
    port map (
            O => \N__25170\,
            I => \N__25132\
        );

    \I__6154\ : Sp12to4
    port map (
            O => \N__25165\,
            I => \N__25129\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__25162\,
            I => \N__25126\
        );

    \I__6152\ : InMux
    port map (
            O => \N__25161\,
            I => \N__25121\
        );

    \I__6151\ : InMux
    port map (
            O => \N__25160\,
            I => \N__25121\
        );

    \I__6150\ : InMux
    port map (
            O => \N__25159\,
            I => \N__25118\
        );

    \I__6149\ : InMux
    port map (
            O => \N__25156\,
            I => \N__25115\
        );

    \I__6148\ : InMux
    port map (
            O => \N__25155\,
            I => \N__25110\
        );

    \I__6147\ : InMux
    port map (
            O => \N__25154\,
            I => \N__25110\
        );

    \I__6146\ : InMux
    port map (
            O => \N__25153\,
            I => \N__25107\
        );

    \I__6145\ : InMux
    port map (
            O => \N__25152\,
            I => \N__25104\
        );

    \I__6144\ : Span4Mux_v
    port map (
            O => \N__25147\,
            I => \N__25097\
        );

    \I__6143\ : Span4Mux_v
    port map (
            O => \N__25144\,
            I => \N__25097\
        );

    \I__6142\ : Span4Mux_v
    port map (
            O => \N__25135\,
            I => \N__25097\
        );

    \I__6141\ : Sp12to4
    port map (
            O => \N__25132\,
            I => \N__25092\
        );

    \I__6140\ : Span12Mux_s3_h
    port map (
            O => \N__25129\,
            I => \N__25092\
        );

    \I__6139\ : Span4Mux_h
    port map (
            O => \N__25126\,
            I => \N__25089\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__25121\,
            I => \N__25082\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__25118\,
            I => \N__25082\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__25115\,
            I => \N__25082\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__25110\,
            I => \N__25079\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__25107\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__25104\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__6132\ : Odrv4
    port map (
            O => \N__25097\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__6131\ : Odrv12
    port map (
            O => \N__25092\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__6130\ : Odrv4
    port map (
            O => \N__25089\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__6129\ : Odrv4
    port map (
            O => \N__25082\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__6128\ : Odrv4
    port map (
            O => \N__25079\,
            I => \M_this_state_qZ0Z_0\
        );

    \I__6127\ : InMux
    port map (
            O => \N__25064\,
            I => \un1_M_this_external_address_q_cry_14\
        );

    \I__6126\ : IoInMux
    port map (
            O => \N__25061\,
            I => \N__25058\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__25058\,
            I => \N__25055\
        );

    \I__6124\ : Span4Mux_s1_h
    port map (
            O => \N__25055\,
            I => \N__25052\
        );

    \I__6123\ : Sp12to4
    port map (
            O => \N__25052\,
            I => \N__25049\
        );

    \I__6122\ : Span12Mux_v
    port map (
            O => \N__25049\,
            I => \N__25045\
        );

    \I__6121\ : InMux
    port map (
            O => \N__25048\,
            I => \N__25042\
        );

    \I__6120\ : Odrv12
    port map (
            O => \N__25045\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__25042\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__6118\ : ClkMux
    port map (
            O => \N__25037\,
            I => \N__24806\
        );

    \I__6117\ : ClkMux
    port map (
            O => \N__25036\,
            I => \N__24806\
        );

    \I__6116\ : ClkMux
    port map (
            O => \N__25035\,
            I => \N__24806\
        );

    \I__6115\ : ClkMux
    port map (
            O => \N__25034\,
            I => \N__24806\
        );

    \I__6114\ : ClkMux
    port map (
            O => \N__25033\,
            I => \N__24806\
        );

    \I__6113\ : ClkMux
    port map (
            O => \N__25032\,
            I => \N__24806\
        );

    \I__6112\ : ClkMux
    port map (
            O => \N__25031\,
            I => \N__24806\
        );

    \I__6111\ : ClkMux
    port map (
            O => \N__25030\,
            I => \N__24806\
        );

    \I__6110\ : ClkMux
    port map (
            O => \N__25029\,
            I => \N__24806\
        );

    \I__6109\ : ClkMux
    port map (
            O => \N__25028\,
            I => \N__24806\
        );

    \I__6108\ : ClkMux
    port map (
            O => \N__25027\,
            I => \N__24806\
        );

    \I__6107\ : ClkMux
    port map (
            O => \N__25026\,
            I => \N__24806\
        );

    \I__6106\ : ClkMux
    port map (
            O => \N__25025\,
            I => \N__24806\
        );

    \I__6105\ : ClkMux
    port map (
            O => \N__25024\,
            I => \N__24806\
        );

    \I__6104\ : ClkMux
    port map (
            O => \N__25023\,
            I => \N__24806\
        );

    \I__6103\ : ClkMux
    port map (
            O => \N__25022\,
            I => \N__24806\
        );

    \I__6102\ : ClkMux
    port map (
            O => \N__25021\,
            I => \N__24806\
        );

    \I__6101\ : ClkMux
    port map (
            O => \N__25020\,
            I => \N__24806\
        );

    \I__6100\ : ClkMux
    port map (
            O => \N__25019\,
            I => \N__24806\
        );

    \I__6099\ : ClkMux
    port map (
            O => \N__25018\,
            I => \N__24806\
        );

    \I__6098\ : ClkMux
    port map (
            O => \N__25017\,
            I => \N__24806\
        );

    \I__6097\ : ClkMux
    port map (
            O => \N__25016\,
            I => \N__24806\
        );

    \I__6096\ : ClkMux
    port map (
            O => \N__25015\,
            I => \N__24806\
        );

    \I__6095\ : ClkMux
    port map (
            O => \N__25014\,
            I => \N__24806\
        );

    \I__6094\ : ClkMux
    port map (
            O => \N__25013\,
            I => \N__24806\
        );

    \I__6093\ : ClkMux
    port map (
            O => \N__25012\,
            I => \N__24806\
        );

    \I__6092\ : ClkMux
    port map (
            O => \N__25011\,
            I => \N__24806\
        );

    \I__6091\ : ClkMux
    port map (
            O => \N__25010\,
            I => \N__24806\
        );

    \I__6090\ : ClkMux
    port map (
            O => \N__25009\,
            I => \N__24806\
        );

    \I__6089\ : ClkMux
    port map (
            O => \N__25008\,
            I => \N__24806\
        );

    \I__6088\ : ClkMux
    port map (
            O => \N__25007\,
            I => \N__24806\
        );

    \I__6087\ : ClkMux
    port map (
            O => \N__25006\,
            I => \N__24806\
        );

    \I__6086\ : ClkMux
    port map (
            O => \N__25005\,
            I => \N__24806\
        );

    \I__6085\ : ClkMux
    port map (
            O => \N__25004\,
            I => \N__24806\
        );

    \I__6084\ : ClkMux
    port map (
            O => \N__25003\,
            I => \N__24806\
        );

    \I__6083\ : ClkMux
    port map (
            O => \N__25002\,
            I => \N__24806\
        );

    \I__6082\ : ClkMux
    port map (
            O => \N__25001\,
            I => \N__24806\
        );

    \I__6081\ : ClkMux
    port map (
            O => \N__25000\,
            I => \N__24806\
        );

    \I__6080\ : ClkMux
    port map (
            O => \N__24999\,
            I => \N__24806\
        );

    \I__6079\ : ClkMux
    port map (
            O => \N__24998\,
            I => \N__24806\
        );

    \I__6078\ : ClkMux
    port map (
            O => \N__24997\,
            I => \N__24806\
        );

    \I__6077\ : ClkMux
    port map (
            O => \N__24996\,
            I => \N__24806\
        );

    \I__6076\ : ClkMux
    port map (
            O => \N__24995\,
            I => \N__24806\
        );

    \I__6075\ : ClkMux
    port map (
            O => \N__24994\,
            I => \N__24806\
        );

    \I__6074\ : ClkMux
    port map (
            O => \N__24993\,
            I => \N__24806\
        );

    \I__6073\ : ClkMux
    port map (
            O => \N__24992\,
            I => \N__24806\
        );

    \I__6072\ : ClkMux
    port map (
            O => \N__24991\,
            I => \N__24806\
        );

    \I__6071\ : ClkMux
    port map (
            O => \N__24990\,
            I => \N__24806\
        );

    \I__6070\ : ClkMux
    port map (
            O => \N__24989\,
            I => \N__24806\
        );

    \I__6069\ : ClkMux
    port map (
            O => \N__24988\,
            I => \N__24806\
        );

    \I__6068\ : ClkMux
    port map (
            O => \N__24987\,
            I => \N__24806\
        );

    \I__6067\ : ClkMux
    port map (
            O => \N__24986\,
            I => \N__24806\
        );

    \I__6066\ : ClkMux
    port map (
            O => \N__24985\,
            I => \N__24806\
        );

    \I__6065\ : ClkMux
    port map (
            O => \N__24984\,
            I => \N__24806\
        );

    \I__6064\ : ClkMux
    port map (
            O => \N__24983\,
            I => \N__24806\
        );

    \I__6063\ : ClkMux
    port map (
            O => \N__24982\,
            I => \N__24806\
        );

    \I__6062\ : ClkMux
    port map (
            O => \N__24981\,
            I => \N__24806\
        );

    \I__6061\ : ClkMux
    port map (
            O => \N__24980\,
            I => \N__24806\
        );

    \I__6060\ : ClkMux
    port map (
            O => \N__24979\,
            I => \N__24806\
        );

    \I__6059\ : ClkMux
    port map (
            O => \N__24978\,
            I => \N__24806\
        );

    \I__6058\ : ClkMux
    port map (
            O => \N__24977\,
            I => \N__24806\
        );

    \I__6057\ : ClkMux
    port map (
            O => \N__24976\,
            I => \N__24806\
        );

    \I__6056\ : ClkMux
    port map (
            O => \N__24975\,
            I => \N__24806\
        );

    \I__6055\ : ClkMux
    port map (
            O => \N__24974\,
            I => \N__24806\
        );

    \I__6054\ : ClkMux
    port map (
            O => \N__24973\,
            I => \N__24806\
        );

    \I__6053\ : ClkMux
    port map (
            O => \N__24972\,
            I => \N__24806\
        );

    \I__6052\ : ClkMux
    port map (
            O => \N__24971\,
            I => \N__24806\
        );

    \I__6051\ : ClkMux
    port map (
            O => \N__24970\,
            I => \N__24806\
        );

    \I__6050\ : ClkMux
    port map (
            O => \N__24969\,
            I => \N__24806\
        );

    \I__6049\ : ClkMux
    port map (
            O => \N__24968\,
            I => \N__24806\
        );

    \I__6048\ : ClkMux
    port map (
            O => \N__24967\,
            I => \N__24806\
        );

    \I__6047\ : ClkMux
    port map (
            O => \N__24966\,
            I => \N__24806\
        );

    \I__6046\ : ClkMux
    port map (
            O => \N__24965\,
            I => \N__24806\
        );

    \I__6045\ : ClkMux
    port map (
            O => \N__24964\,
            I => \N__24806\
        );

    \I__6044\ : ClkMux
    port map (
            O => \N__24963\,
            I => \N__24806\
        );

    \I__6043\ : ClkMux
    port map (
            O => \N__24962\,
            I => \N__24806\
        );

    \I__6042\ : ClkMux
    port map (
            O => \N__24961\,
            I => \N__24806\
        );

    \I__6041\ : GlobalMux
    port map (
            O => \N__24806\,
            I => \N__24803\
        );

    \I__6040\ : gio2CtrlBuf
    port map (
            O => \N__24803\,
            I => clk_0_c_g
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__24800\,
            I => \N__24795\
        );

    \I__6038\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24781\
        );

    \I__6037\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24778\
        );

    \I__6036\ : InMux
    port map (
            O => \N__24795\,
            I => \N__24775\
        );

    \I__6035\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24770\
        );

    \I__6034\ : InMux
    port map (
            O => \N__24793\,
            I => \N__24770\
        );

    \I__6033\ : InMux
    port map (
            O => \N__24792\,
            I => \N__24765\
        );

    \I__6032\ : InMux
    port map (
            O => \N__24791\,
            I => \N__24765\
        );

    \I__6031\ : InMux
    port map (
            O => \N__24790\,
            I => \N__24762\
        );

    \I__6030\ : InMux
    port map (
            O => \N__24789\,
            I => \N__24757\
        );

    \I__6029\ : InMux
    port map (
            O => \N__24788\,
            I => \N__24757\
        );

    \I__6028\ : InMux
    port map (
            O => \N__24787\,
            I => \N__24754\
        );

    \I__6027\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24751\
        );

    \I__6026\ : InMux
    port map (
            O => \N__24785\,
            I => \N__24746\
        );

    \I__6025\ : InMux
    port map (
            O => \N__24784\,
            I => \N__24746\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__24781\,
            I => \N__24728\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__24778\,
            I => \N__24725\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__24775\,
            I => \N__24722\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__24770\,
            I => \N__24719\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__24765\,
            I => \N__24716\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__24762\,
            I => \N__24713\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__24757\,
            I => \N__24710\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__24754\,
            I => \N__24707\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__24751\,
            I => \N__24704\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__24746\,
            I => \N__24701\
        );

    \I__6014\ : SRMux
    port map (
            O => \N__24745\,
            I => \N__24650\
        );

    \I__6013\ : SRMux
    port map (
            O => \N__24744\,
            I => \N__24650\
        );

    \I__6012\ : SRMux
    port map (
            O => \N__24743\,
            I => \N__24650\
        );

    \I__6011\ : SRMux
    port map (
            O => \N__24742\,
            I => \N__24650\
        );

    \I__6010\ : SRMux
    port map (
            O => \N__24741\,
            I => \N__24650\
        );

    \I__6009\ : SRMux
    port map (
            O => \N__24740\,
            I => \N__24650\
        );

    \I__6008\ : SRMux
    port map (
            O => \N__24739\,
            I => \N__24650\
        );

    \I__6007\ : SRMux
    port map (
            O => \N__24738\,
            I => \N__24650\
        );

    \I__6006\ : SRMux
    port map (
            O => \N__24737\,
            I => \N__24650\
        );

    \I__6005\ : SRMux
    port map (
            O => \N__24736\,
            I => \N__24650\
        );

    \I__6004\ : SRMux
    port map (
            O => \N__24735\,
            I => \N__24650\
        );

    \I__6003\ : SRMux
    port map (
            O => \N__24734\,
            I => \N__24650\
        );

    \I__6002\ : SRMux
    port map (
            O => \N__24733\,
            I => \N__24650\
        );

    \I__6001\ : SRMux
    port map (
            O => \N__24732\,
            I => \N__24650\
        );

    \I__6000\ : SRMux
    port map (
            O => \N__24731\,
            I => \N__24650\
        );

    \I__5999\ : Glb2LocalMux
    port map (
            O => \N__24728\,
            I => \N__24650\
        );

    \I__5998\ : Glb2LocalMux
    port map (
            O => \N__24725\,
            I => \N__24650\
        );

    \I__5997\ : Glb2LocalMux
    port map (
            O => \N__24722\,
            I => \N__24650\
        );

    \I__5996\ : Glb2LocalMux
    port map (
            O => \N__24719\,
            I => \N__24650\
        );

    \I__5995\ : Glb2LocalMux
    port map (
            O => \N__24716\,
            I => \N__24650\
        );

    \I__5994\ : Glb2LocalMux
    port map (
            O => \N__24713\,
            I => \N__24650\
        );

    \I__5993\ : Glb2LocalMux
    port map (
            O => \N__24710\,
            I => \N__24650\
        );

    \I__5992\ : Glb2LocalMux
    port map (
            O => \N__24707\,
            I => \N__24650\
        );

    \I__5991\ : Glb2LocalMux
    port map (
            O => \N__24704\,
            I => \N__24650\
        );

    \I__5990\ : Glb2LocalMux
    port map (
            O => \N__24701\,
            I => \N__24650\
        );

    \I__5989\ : GlobalMux
    port map (
            O => \N__24650\,
            I => \N__24647\
        );

    \I__5988\ : gio2CtrlBuf
    port map (
            O => \N__24647\,
            I => \M_this_state_q_nss_g_0\
        );

    \I__5987\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24641\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__24641\,
            I => \N__24638\
        );

    \I__5985\ : Span12Mux_s10_h
    port map (
            O => \N__24638\,
            I => \N__24635\
        );

    \I__5984\ : Odrv12
    port map (
            O => \N__24635\,
            I => port_address_in_2
        );

    \I__5983\ : InMux
    port map (
            O => \N__24632\,
            I => \N__24629\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__24629\,
            I => \N__24626\
        );

    \I__5981\ : Span12Mux_v
    port map (
            O => \N__24626\,
            I => \N__24623\
        );

    \I__5980\ : Odrv12
    port map (
            O => \N__24623\,
            I => port_address_in_3
        );

    \I__5979\ : CascadeMux
    port map (
            O => \N__24620\,
            I => \N__24617\
        );

    \I__5978\ : InMux
    port map (
            O => \N__24617\,
            I => \N__24614\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__24614\,
            I => port_address_in_4
        );

    \I__5976\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__24608\,
            I => \N__24605\
        );

    \I__5974\ : Span4Mux_v
    port map (
            O => \N__24605\,
            I => \N__24602\
        );

    \I__5973\ : Odrv4
    port map (
            O => \N__24602\,
            I => port_address_in_5
        );

    \I__5972\ : InMux
    port map (
            O => \N__24599\,
            I => \N__24596\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__24596\,
            I => \N__24592\
        );

    \I__5970\ : InMux
    port map (
            O => \N__24595\,
            I => \N__24589\
        );

    \I__5969\ : Span4Mux_h
    port map (
            O => \N__24592\,
            I => \N__24586\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__24589\,
            I => \N__24583\
        );

    \I__5967\ : Sp12to4
    port map (
            O => \N__24586\,
            I => \N__24580\
        );

    \I__5966\ : Span4Mux_v
    port map (
            O => \N__24583\,
            I => \N__24577\
        );

    \I__5965\ : Span12Mux_v
    port map (
            O => \N__24580\,
            I => \N__24572\
        );

    \I__5964\ : Sp12to4
    port map (
            O => \N__24577\,
            I => \N__24572\
        );

    \I__5963\ : Span12Mux_h
    port map (
            O => \N__24572\,
            I => \N__24569\
        );

    \I__5962\ : Odrv12
    port map (
            O => \N__24569\,
            I => \this_vga_signals.M_this_state_q_srsts_0_i_o4_5Z0Z_4\
        );

    \I__5961\ : InMux
    port map (
            O => \N__24566\,
            I => \un1_M_this_external_address_q_cry_3\
        );

    \I__5960\ : IoInMux
    port map (
            O => \N__24563\,
            I => \N__24560\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__24560\,
            I => \N__24557\
        );

    \I__5958\ : Span4Mux_s1_h
    port map (
            O => \N__24557\,
            I => \N__24553\
        );

    \I__5957\ : InMux
    port map (
            O => \N__24556\,
            I => \N__24550\
        );

    \I__5956\ : Odrv4
    port map (
            O => \N__24553\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__24550\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__5954\ : InMux
    port map (
            O => \N__24545\,
            I => \un1_M_this_external_address_q_cry_4\
        );

    \I__5953\ : IoInMux
    port map (
            O => \N__24542\,
            I => \N__24539\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__5951\ : Span12Mux_s1_h
    port map (
            O => \N__24536\,
            I => \N__24532\
        );

    \I__5950\ : InMux
    port map (
            O => \N__24535\,
            I => \N__24529\
        );

    \I__5949\ : Odrv12
    port map (
            O => \N__24532\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__24529\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__5947\ : InMux
    port map (
            O => \N__24524\,
            I => \un1_M_this_external_address_q_cry_5\
        );

    \I__5946\ : IoInMux
    port map (
            O => \N__24521\,
            I => \N__24518\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__24518\,
            I => \N__24515\
        );

    \I__5944\ : Span4Mux_s1_h
    port map (
            O => \N__24515\,
            I => \N__24512\
        );

    \I__5943\ : Sp12to4
    port map (
            O => \N__24512\,
            I => \N__24509\
        );

    \I__5942\ : Span12Mux_v
    port map (
            O => \N__24509\,
            I => \N__24505\
        );

    \I__5941\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24502\
        );

    \I__5940\ : Odrv12
    port map (
            O => \N__24505\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__24502\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__5938\ : InMux
    port map (
            O => \N__24497\,
            I => \un1_M_this_external_address_q_cry_6\
        );

    \I__5937\ : IoInMux
    port map (
            O => \N__24494\,
            I => \N__24491\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__24491\,
            I => \N__24488\
        );

    \I__5935\ : Span4Mux_s0_v
    port map (
            O => \N__24488\,
            I => \N__24485\
        );

    \I__5934\ : Span4Mux_h
    port map (
            O => \N__24485\,
            I => \N__24482\
        );

    \I__5933\ : Sp12to4
    port map (
            O => \N__24482\,
            I => \N__24479\
        );

    \I__5932\ : Span12Mux_h
    port map (
            O => \N__24479\,
            I => \N__24475\
        );

    \I__5931\ : InMux
    port map (
            O => \N__24478\,
            I => \N__24472\
        );

    \I__5930\ : Odrv12
    port map (
            O => \N__24475\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__24472\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__5928\ : InMux
    port map (
            O => \N__24467\,
            I => \bfn_31_24_0_\
        );

    \I__5927\ : IoInMux
    port map (
            O => \N__24464\,
            I => \N__24461\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__24461\,
            I => \N__24458\
        );

    \I__5925\ : IoSpan4Mux
    port map (
            O => \N__24458\,
            I => \N__24455\
        );

    \I__5924\ : IoSpan4Mux
    port map (
            O => \N__24455\,
            I => \N__24452\
        );

    \I__5923\ : IoSpan4Mux
    port map (
            O => \N__24452\,
            I => \N__24449\
        );

    \I__5922\ : IoSpan4Mux
    port map (
            O => \N__24449\,
            I => \N__24445\
        );

    \I__5921\ : InMux
    port map (
            O => \N__24448\,
            I => \N__24442\
        );

    \I__5920\ : Odrv4
    port map (
            O => \N__24445\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__24442\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__5918\ : InMux
    port map (
            O => \N__24437\,
            I => \un1_M_this_external_address_q_cry_8\
        );

    \I__5917\ : IoInMux
    port map (
            O => \N__24434\,
            I => \N__24431\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__24431\,
            I => \N__24428\
        );

    \I__5915\ : Span4Mux_s2_v
    port map (
            O => \N__24428\,
            I => \N__24425\
        );

    \I__5914\ : Span4Mux_v
    port map (
            O => \N__24425\,
            I => \N__24422\
        );

    \I__5913\ : Sp12to4
    port map (
            O => \N__24422\,
            I => \N__24419\
        );

    \I__5912\ : Span12Mux_h
    port map (
            O => \N__24419\,
            I => \N__24415\
        );

    \I__5911\ : InMux
    port map (
            O => \N__24418\,
            I => \N__24412\
        );

    \I__5910\ : Odrv12
    port map (
            O => \N__24415\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__24412\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__5908\ : InMux
    port map (
            O => \N__24407\,
            I => \un1_M_this_external_address_q_cry_9\
        );

    \I__5907\ : IoInMux
    port map (
            O => \N__24404\,
            I => \N__24401\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__24401\,
            I => \N__24398\
        );

    \I__5905\ : Span4Mux_s0_v
    port map (
            O => \N__24398\,
            I => \N__24395\
        );

    \I__5904\ : Span4Mux_v
    port map (
            O => \N__24395\,
            I => \N__24392\
        );

    \I__5903\ : Span4Mux_v
    port map (
            O => \N__24392\,
            I => \N__24388\
        );

    \I__5902\ : InMux
    port map (
            O => \N__24391\,
            I => \N__24385\
        );

    \I__5901\ : Odrv4
    port map (
            O => \N__24388\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__24385\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__5899\ : InMux
    port map (
            O => \N__24380\,
            I => \un1_M_this_external_address_q_cry_10\
        );

    \I__5898\ : IoInMux
    port map (
            O => \N__24377\,
            I => \N__24374\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__24374\,
            I => \N__24370\
        );

    \I__5896\ : InMux
    port map (
            O => \N__24373\,
            I => \N__24367\
        );

    \I__5895\ : Odrv12
    port map (
            O => \N__24370\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__24367\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__5893\ : InMux
    port map (
            O => \N__24362\,
            I => \un1_M_this_external_address_q_cry_11\
        );

    \I__5892\ : InMux
    port map (
            O => \N__24359\,
            I => \N__24355\
        );

    \I__5891\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24351\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__24355\,
            I => \N__24348\
        );

    \I__5889\ : InMux
    port map (
            O => \N__24354\,
            I => \N__24345\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__24351\,
            I => \N__24341\
        );

    \I__5887\ : Span4Mux_h
    port map (
            O => \N__24348\,
            I => \N__24338\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__24345\,
            I => \N__24335\
        );

    \I__5885\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24332\
        );

    \I__5884\ : Span12Mux_h
    port map (
            O => \N__24341\,
            I => \N__24329\
        );

    \I__5883\ : Span4Mux_h
    port map (
            O => \N__24338\,
            I => \N__24326\
        );

    \I__5882\ : Span4Mux_v
    port map (
            O => \N__24335\,
            I => \N__24321\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__24332\,
            I => \N__24321\
        );

    \I__5880\ : Odrv12
    port map (
            O => \N__24329\,
            I => \this_vga_signals.N_479\
        );

    \I__5879\ : Odrv4
    port map (
            O => \N__24326\,
            I => \this_vga_signals.N_479\
        );

    \I__5878\ : Odrv4
    port map (
            O => \N__24321\,
            I => \this_vga_signals.N_479\
        );

    \I__5877\ : InMux
    port map (
            O => \N__24314\,
            I => \N__24311\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__24311\,
            I => \N__24306\
        );

    \I__5875\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24303\
        );

    \I__5874\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24299\
        );

    \I__5873\ : Span4Mux_h
    port map (
            O => \N__24306\,
            I => \N__24295\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__24303\,
            I => \N__24292\
        );

    \I__5871\ : InMux
    port map (
            O => \N__24302\,
            I => \N__24289\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__24299\,
            I => \N__24285\
        );

    \I__5869\ : InMux
    port map (
            O => \N__24298\,
            I => \N__24282\
        );

    \I__5868\ : Span4Mux_v
    port map (
            O => \N__24295\,
            I => \N__24276\
        );

    \I__5867\ : Span4Mux_h
    port map (
            O => \N__24292\,
            I => \N__24276\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__24289\,
            I => \N__24273\
        );

    \I__5865\ : InMux
    port map (
            O => \N__24288\,
            I => \N__24270\
        );

    \I__5864\ : Span4Mux_v
    port map (
            O => \N__24285\,
            I => \N__24265\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__24282\,
            I => \N__24265\
        );

    \I__5862\ : InMux
    port map (
            O => \N__24281\,
            I => \N__24262\
        );

    \I__5861\ : Span4Mux_v
    port map (
            O => \N__24276\,
            I => \N__24257\
        );

    \I__5860\ : Span4Mux_h
    port map (
            O => \N__24273\,
            I => \N__24257\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__24270\,
            I => \N__24254\
        );

    \I__5858\ : Span4Mux_v
    port map (
            O => \N__24265\,
            I => \N__24249\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__24262\,
            I => \N__24249\
        );

    \I__5856\ : Span4Mux_v
    port map (
            O => \N__24257\,
            I => \N__24243\
        );

    \I__5855\ : Span4Mux_h
    port map (
            O => \N__24254\,
            I => \N__24243\
        );

    \I__5854\ : Span4Mux_v
    port map (
            O => \N__24249\,
            I => \N__24240\
        );

    \I__5853\ : InMux
    port map (
            O => \N__24248\,
            I => \N__24237\
        );

    \I__5852\ : Odrv4
    port map (
            O => \N__24243\,
            I => \M_this_sprites_ram_write_data_2\
        );

    \I__5851\ : Odrv4
    port map (
            O => \N__24240\,
            I => \M_this_sprites_ram_write_data_2\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__24237\,
            I => \M_this_sprites_ram_write_data_2\
        );

    \I__5849\ : CEMux
    port map (
            O => \N__24230\,
            I => \N__24227\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__24227\,
            I => \N__24223\
        );

    \I__5847\ : CEMux
    port map (
            O => \N__24226\,
            I => \N__24220\
        );

    \I__5846\ : Span4Mux_h
    port map (
            O => \N__24223\,
            I => \N__24217\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__24220\,
            I => \N__24214\
        );

    \I__5844\ : Odrv4
    port map (
            O => \N__24217\,
            I => \this_sprites_ram.mem_WE_4\
        );

    \I__5843\ : Odrv12
    port map (
            O => \N__24214\,
            I => \this_sprites_ram.mem_WE_4\
        );

    \I__5842\ : InMux
    port map (
            O => \N__24209\,
            I => \N__24203\
        );

    \I__5841\ : InMux
    port map (
            O => \N__24208\,
            I => \N__24198\
        );

    \I__5840\ : InMux
    port map (
            O => \N__24207\,
            I => \N__24198\
        );

    \I__5839\ : InMux
    port map (
            O => \N__24206\,
            I => \N__24195\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__24203\,
            I => \N__24191\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__24198\,
            I => \N__24186\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__24195\,
            I => \N__24186\
        );

    \I__5835\ : InMux
    port map (
            O => \N__24194\,
            I => \N__24183\
        );

    \I__5834\ : Span4Mux_v
    port map (
            O => \N__24191\,
            I => \N__24176\
        );

    \I__5833\ : Span4Mux_v
    port map (
            O => \N__24186\,
            I => \N__24176\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__24183\,
            I => \N__24176\
        );

    \I__5831\ : Span4Mux_v
    port map (
            O => \N__24176\,
            I => \N__24170\
        );

    \I__5830\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24164\
        );

    \I__5829\ : InMux
    port map (
            O => \N__24174\,
            I => \N__24164\
        );

    \I__5828\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24161\
        );

    \I__5827\ : Span4Mux_v
    port map (
            O => \N__24170\,
            I => \N__24157\
        );

    \I__5826\ : InMux
    port map (
            O => \N__24169\,
            I => \N__24154\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__24164\,
            I => \N__24149\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__24161\,
            I => \N__24149\
        );

    \I__5823\ : InMux
    port map (
            O => \N__24160\,
            I => \N__24146\
        );

    \I__5822\ : Span4Mux_h
    port map (
            O => \N__24157\,
            I => \N__24141\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__24154\,
            I => \N__24141\
        );

    \I__5820\ : Odrv12
    port map (
            O => \N__24149\,
            I => \M_this_internal_address_qZ0Z_12\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__24146\,
            I => \M_this_internal_address_qZ0Z_12\
        );

    \I__5818\ : Odrv4
    port map (
            O => \N__24141\,
            I => \M_this_internal_address_qZ0Z_12\
        );

    \I__5817\ : CascadeMux
    port map (
            O => \N__24134\,
            I => \N__24131\
        );

    \I__5816\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24124\
        );

    \I__5815\ : InMux
    port map (
            O => \N__24130\,
            I => \N__24124\
        );

    \I__5814\ : InMux
    port map (
            O => \N__24129\,
            I => \N__24121\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__24124\,
            I => \N__24115\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__24121\,
            I => \N__24115\
        );

    \I__5811\ : InMux
    port map (
            O => \N__24120\,
            I => \N__24112\
        );

    \I__5810\ : Span4Mux_v
    port map (
            O => \N__24115\,
            I => \N__24107\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__24112\,
            I => \N__24107\
        );

    \I__5808\ : Span4Mux_h
    port map (
            O => \N__24107\,
            I => \N__24104\
        );

    \I__5807\ : Span4Mux_v
    port map (
            O => \N__24104\,
            I => \N__24100\
        );

    \I__5806\ : InMux
    port map (
            O => \N__24103\,
            I => \N__24097\
        );

    \I__5805\ : Sp12to4
    port map (
            O => \N__24100\,
            I => \N__24089\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__24097\,
            I => \N__24089\
        );

    \I__5803\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24084\
        );

    \I__5802\ : InMux
    port map (
            O => \N__24095\,
            I => \N__24084\
        );

    \I__5801\ : InMux
    port map (
            O => \N__24094\,
            I => \N__24081\
        );

    \I__5800\ : Span12Mux_h
    port map (
            O => \N__24089\,
            I => \N__24076\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__24084\,
            I => \N__24071\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__24081\,
            I => \N__24071\
        );

    \I__5797\ : InMux
    port map (
            O => \N__24080\,
            I => \N__24068\
        );

    \I__5796\ : InMux
    port map (
            O => \N__24079\,
            I => \N__24065\
        );

    \I__5795\ : Odrv12
    port map (
            O => \N__24076\,
            I => \M_this_internal_address_qZ0Z_11\
        );

    \I__5794\ : Odrv12
    port map (
            O => \N__24071\,
            I => \M_this_internal_address_qZ0Z_11\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__24068\,
            I => \M_this_internal_address_qZ0Z_11\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__24065\,
            I => \M_this_internal_address_qZ0Z_11\
        );

    \I__5791\ : CascadeMux
    port map (
            O => \N__24056\,
            I => \N__24048\
        );

    \I__5790\ : CascadeMux
    port map (
            O => \N__24055\,
            I => \N__24045\
        );

    \I__5789\ : CascadeMux
    port map (
            O => \N__24054\,
            I => \N__24042\
        );

    \I__5788\ : CascadeMux
    port map (
            O => \N__24053\,
            I => \N__24038\
        );

    \I__5787\ : CascadeMux
    port map (
            O => \N__24052\,
            I => \N__24035\
        );

    \I__5786\ : CascadeMux
    port map (
            O => \N__24051\,
            I => \N__24031\
        );

    \I__5785\ : InMux
    port map (
            O => \N__24048\,
            I => \N__24027\
        );

    \I__5784\ : InMux
    port map (
            O => \N__24045\,
            I => \N__24022\
        );

    \I__5783\ : InMux
    port map (
            O => \N__24042\,
            I => \N__24022\
        );

    \I__5782\ : CascadeMux
    port map (
            O => \N__24041\,
            I => \N__24019\
        );

    \I__5781\ : InMux
    port map (
            O => \N__24038\,
            I => \N__24016\
        );

    \I__5780\ : InMux
    port map (
            O => \N__24035\,
            I => \N__24013\
        );

    \I__5779\ : InMux
    port map (
            O => \N__24034\,
            I => \N__24008\
        );

    \I__5778\ : InMux
    port map (
            O => \N__24031\,
            I => \N__24008\
        );

    \I__5777\ : InMux
    port map (
            O => \N__24030\,
            I => \N__24005\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__24027\,
            I => \N__24002\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__24022\,
            I => \N__23999\
        );

    \I__5774\ : InMux
    port map (
            O => \N__24019\,
            I => \N__23996\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__24016\,
            I => \N__23989\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__24013\,
            I => \N__23989\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__24008\,
            I => \N__23989\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__24005\,
            I => \N__23985\
        );

    \I__5769\ : Span4Mux_h
    port map (
            O => \N__24002\,
            I => \N__23982\
        );

    \I__5768\ : Span4Mux_v
    port map (
            O => \N__23999\,
            I => \N__23979\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__23996\,
            I => \N__23976\
        );

    \I__5766\ : Span4Mux_v
    port map (
            O => \N__23989\,
            I => \N__23973\
        );

    \I__5765\ : InMux
    port map (
            O => \N__23988\,
            I => \N__23970\
        );

    \I__5764\ : Span4Mux_v
    port map (
            O => \N__23985\,
            I => \N__23963\
        );

    \I__5763\ : Span4Mux_v
    port map (
            O => \N__23982\,
            I => \N__23963\
        );

    \I__5762\ : Span4Mux_h
    port map (
            O => \N__23979\,
            I => \N__23963\
        );

    \I__5761\ : Span4Mux_v
    port map (
            O => \N__23976\,
            I => \N__23960\
        );

    \I__5760\ : Sp12to4
    port map (
            O => \N__23973\,
            I => \N__23957\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__23970\,
            I => \N__23950\
        );

    \I__5758\ : Sp12to4
    port map (
            O => \N__23963\,
            I => \N__23950\
        );

    \I__5757\ : Sp12to4
    port map (
            O => \N__23960\,
            I => \N__23950\
        );

    \I__5756\ : Span12Mux_h
    port map (
            O => \N__23957\,
            I => \N__23947\
        );

    \I__5755\ : Odrv12
    port map (
            O => \N__23950\,
            I => \M_this_internal_address_qZ0Z_13\
        );

    \I__5754\ : Odrv12
    port map (
            O => \N__23947\,
            I => \M_this_internal_address_qZ0Z_13\
        );

    \I__5753\ : InMux
    port map (
            O => \N__23942\,
            I => \N__23935\
        );

    \I__5752\ : InMux
    port map (
            O => \N__23941\,
            I => \N__23935\
        );

    \I__5751\ : InMux
    port map (
            O => \N__23940\,
            I => \N__23932\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__23935\,
            I => \N__23926\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__23932\,
            I => \N__23923\
        );

    \I__5748\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23920\
        );

    \I__5747\ : InMux
    port map (
            O => \N__23930\,
            I => \N__23913\
        );

    \I__5746\ : InMux
    port map (
            O => \N__23929\,
            I => \N__23913\
        );

    \I__5745\ : Span4Mux_v
    port map (
            O => \N__23926\,
            I => \N__23906\
        );

    \I__5744\ : Span4Mux_h
    port map (
            O => \N__23923\,
            I => \N__23906\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__23920\,
            I => \N__23906\
        );

    \I__5742\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23903\
        );

    \I__5741\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23900\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__23913\,
            I => \N__23897\
        );

    \I__5739\ : Span4Mux_v
    port map (
            O => \N__23906\,
            I => \N__23892\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__23903\,
            I => \N__23892\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__23900\,
            I => \N__23889\
        );

    \I__5736\ : Odrv4
    port map (
            O => \N__23897\,
            I => \N_24_0\
        );

    \I__5735\ : Odrv4
    port map (
            O => \N__23892\,
            I => \N_24_0\
        );

    \I__5734\ : Odrv4
    port map (
            O => \N__23889\,
            I => \N_24_0\
        );

    \I__5733\ : CEMux
    port map (
            O => \N__23882\,
            I => \N__23879\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__23879\,
            I => \N__23875\
        );

    \I__5731\ : CEMux
    port map (
            O => \N__23878\,
            I => \N__23872\
        );

    \I__5730\ : Span4Mux_v
    port map (
            O => \N__23875\,
            I => \N__23867\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__23872\,
            I => \N__23867\
        );

    \I__5728\ : Span4Mux_v
    port map (
            O => \N__23867\,
            I => \N__23864\
        );

    \I__5727\ : Odrv4
    port map (
            O => \N__23864\,
            I => \this_sprites_ram.mem_WE_2\
        );

    \I__5726\ : CascadeMux
    port map (
            O => \N__23861\,
            I => \N__23847\
        );

    \I__5725\ : InMux
    port map (
            O => \N__23860\,
            I => \N__23844\
        );

    \I__5724\ : InMux
    port map (
            O => \N__23859\,
            I => \N__23839\
        );

    \I__5723\ : InMux
    port map (
            O => \N__23858\,
            I => \N__23834\
        );

    \I__5722\ : InMux
    port map (
            O => \N__23857\,
            I => \N__23834\
        );

    \I__5721\ : CascadeMux
    port map (
            O => \N__23856\,
            I => \N__23831\
        );

    \I__5720\ : InMux
    port map (
            O => \N__23855\,
            I => \N__23827\
        );

    \I__5719\ : InMux
    port map (
            O => \N__23854\,
            I => \N__23824\
        );

    \I__5718\ : InMux
    port map (
            O => \N__23853\,
            I => \N__23818\
        );

    \I__5717\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23818\
        );

    \I__5716\ : InMux
    port map (
            O => \N__23851\,
            I => \N__23815\
        );

    \I__5715\ : InMux
    port map (
            O => \N__23850\,
            I => \N__23812\
        );

    \I__5714\ : InMux
    port map (
            O => \N__23847\,
            I => \N__23809\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__23844\,
            I => \N__23806\
        );

    \I__5712\ : CascadeMux
    port map (
            O => \N__23843\,
            I => \N__23803\
        );

    \I__5711\ : InMux
    port map (
            O => \N__23842\,
            I => \N__23800\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__23839\,
            I => \N__23797\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__23834\,
            I => \N__23794\
        );

    \I__5708\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23789\
        );

    \I__5707\ : InMux
    port map (
            O => \N__23830\,
            I => \N__23789\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__23827\,
            I => \N__23786\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__23824\,
            I => \N__23783\
        );

    \I__5704\ : InMux
    port map (
            O => \N__23823\,
            I => \N__23780\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__23818\,
            I => \N__23777\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__23815\,
            I => \N__23772\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__23812\,
            I => \N__23772\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__23809\,
            I => \N__23769\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__23806\,
            I => \N__23766\
        );

    \I__5698\ : InMux
    port map (
            O => \N__23803\,
            I => \N__23763\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__23800\,
            I => \N__23760\
        );

    \I__5696\ : Span4Mux_v
    port map (
            O => \N__23797\,
            I => \N__23753\
        );

    \I__5695\ : Span4Mux_v
    port map (
            O => \N__23794\,
            I => \N__23753\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__23789\,
            I => \N__23753\
        );

    \I__5693\ : Span12Mux_s7_v
    port map (
            O => \N__23786\,
            I => \N__23750\
        );

    \I__5692\ : Sp12to4
    port map (
            O => \N__23783\,
            I => \N__23747\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__23780\,
            I => \N__23744\
        );

    \I__5690\ : Span4Mux_v
    port map (
            O => \N__23777\,
            I => \N__23739\
        );

    \I__5689\ : Span4Mux_v
    port map (
            O => \N__23772\,
            I => \N__23739\
        );

    \I__5688\ : Span4Mux_v
    port map (
            O => \N__23769\,
            I => \N__23736\
        );

    \I__5687\ : Span4Mux_h
    port map (
            O => \N__23766\,
            I => \N__23731\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__23763\,
            I => \N__23731\
        );

    \I__5685\ : Span4Mux_v
    port map (
            O => \N__23760\,
            I => \N__23728\
        );

    \I__5684\ : Span4Mux_h
    port map (
            O => \N__23753\,
            I => \N__23725\
        );

    \I__5683\ : Span12Mux_h
    port map (
            O => \N__23750\,
            I => \N__23718\
        );

    \I__5682\ : Span12Mux_v
    port map (
            O => \N__23747\,
            I => \N__23718\
        );

    \I__5681\ : Span12Mux_s11_h
    port map (
            O => \N__23744\,
            I => \N__23718\
        );

    \I__5680\ : Span4Mux_v
    port map (
            O => \N__23739\,
            I => \N__23709\
        );

    \I__5679\ : Span4Mux_h
    port map (
            O => \N__23736\,
            I => \N__23709\
        );

    \I__5678\ : Span4Mux_v
    port map (
            O => \N__23731\,
            I => \N__23709\
        );

    \I__5677\ : Span4Mux_h
    port map (
            O => \N__23728\,
            I => \N__23709\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__23725\,
            I => \N_192_0\
        );

    \I__5675\ : Odrv12
    port map (
            O => \N__23718\,
            I => \N_192_0\
        );

    \I__5674\ : Odrv4
    port map (
            O => \N__23709\,
            I => \N_192_0\
        );

    \I__5673\ : InMux
    port map (
            O => \N__23702\,
            I => \N__23699\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__23699\,
            I => \N__23696\
        );

    \I__5671\ : Span12Mux_h
    port map (
            O => \N__23696\,
            I => \N__23693\
        );

    \I__5670\ : Span12Mux_v
    port map (
            O => \N__23693\,
            I => \N__23687\
        );

    \I__5669\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23684\
        );

    \I__5668\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23681\
        );

    \I__5667\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23678\
        );

    \I__5666\ : Odrv12
    port map (
            O => \N__23687\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__23684\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__23681\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__23678\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2
        );

    \I__5662\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23666\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__23666\,
            I => \N__23663\
        );

    \I__5660\ : Span12Mux_h
    port map (
            O => \N__23663\,
            I => \N__23660\
        );

    \I__5659\ : Span12Mux_v
    port map (
            O => \N__23660\,
            I => \N__23657\
        );

    \I__5658\ : Odrv12
    port map (
            O => \N__23657\,
            I => \this_ppu.sprites_N_6\
        );

    \I__5657\ : CascadeMux
    port map (
            O => \N__23654\,
            I => \N__23651\
        );

    \I__5656\ : CascadeBuf
    port map (
            O => \N__23651\,
            I => \N__23648\
        );

    \I__5655\ : CascadeMux
    port map (
            O => \N__23648\,
            I => \N__23645\
        );

    \I__5654\ : CascadeBuf
    port map (
            O => \N__23645\,
            I => \N__23642\
        );

    \I__5653\ : CascadeMux
    port map (
            O => \N__23642\,
            I => \N__23639\
        );

    \I__5652\ : CascadeBuf
    port map (
            O => \N__23639\,
            I => \N__23636\
        );

    \I__5651\ : CascadeMux
    port map (
            O => \N__23636\,
            I => \N__23633\
        );

    \I__5650\ : CascadeBuf
    port map (
            O => \N__23633\,
            I => \N__23630\
        );

    \I__5649\ : CascadeMux
    port map (
            O => \N__23630\,
            I => \N__23627\
        );

    \I__5648\ : CascadeBuf
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__23624\,
            I => \N__23621\
        );

    \I__5646\ : CascadeBuf
    port map (
            O => \N__23621\,
            I => \N__23618\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__5644\ : CascadeBuf
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__5643\ : CascadeMux
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__5642\ : CascadeBuf
    port map (
            O => \N__23609\,
            I => \N__23606\
        );

    \I__5641\ : CascadeMux
    port map (
            O => \N__23606\,
            I => \N__23603\
        );

    \I__5640\ : CascadeBuf
    port map (
            O => \N__23603\,
            I => \N__23600\
        );

    \I__5639\ : CascadeMux
    port map (
            O => \N__23600\,
            I => \N__23597\
        );

    \I__5638\ : CascadeBuf
    port map (
            O => \N__23597\,
            I => \N__23594\
        );

    \I__5637\ : CascadeMux
    port map (
            O => \N__23594\,
            I => \N__23591\
        );

    \I__5636\ : CascadeBuf
    port map (
            O => \N__23591\,
            I => \N__23588\
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__23588\,
            I => \N__23585\
        );

    \I__5634\ : CascadeBuf
    port map (
            O => \N__23585\,
            I => \N__23582\
        );

    \I__5633\ : CascadeMux
    port map (
            O => \N__23582\,
            I => \N__23579\
        );

    \I__5632\ : CascadeBuf
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__5631\ : CascadeMux
    port map (
            O => \N__23576\,
            I => \N__23573\
        );

    \I__5630\ : CascadeBuf
    port map (
            O => \N__23573\,
            I => \N__23570\
        );

    \I__5629\ : CascadeMux
    port map (
            O => \N__23570\,
            I => \N__23567\
        );

    \I__5628\ : CascadeBuf
    port map (
            O => \N__23567\,
            I => \N__23564\
        );

    \I__5627\ : CascadeMux
    port map (
            O => \N__23564\,
            I => \N__23561\
        );

    \I__5626\ : InMux
    port map (
            O => \N__23561\,
            I => \N__23558\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__23558\,
            I => \N__23555\
        );

    \I__5624\ : Odrv4
    port map (
            O => \N__23555\,
            I => sprites_m7
        );

    \I__5623\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23549\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__23549\,
            I => \N__23537\
        );

    \I__5621\ : CascadeMux
    port map (
            O => \N__23548\,
            I => \N__23531\
        );

    \I__5620\ : CascadeMux
    port map (
            O => \N__23547\,
            I => \N__23527\
        );

    \I__5619\ : CascadeMux
    port map (
            O => \N__23546\,
            I => \N__23523\
        );

    \I__5618\ : CascadeMux
    port map (
            O => \N__23545\,
            I => \N__23519\
        );

    \I__5617\ : CascadeMux
    port map (
            O => \N__23544\,
            I => \N__23516\
        );

    \I__5616\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23513\
        );

    \I__5615\ : CascadeMux
    port map (
            O => \N__23542\,
            I => \N__23510\
        );

    \I__5614\ : CascadeMux
    port map (
            O => \N__23541\,
            I => \N__23506\
        );

    \I__5613\ : CascadeMux
    port map (
            O => \N__23540\,
            I => \N__23502\
        );

    \I__5612\ : Span4Mux_h
    port map (
            O => \N__23537\,
            I => \N__23497\
        );

    \I__5611\ : InMux
    port map (
            O => \N__23536\,
            I => \N__23494\
        );

    \I__5610\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23491\
        );

    \I__5609\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23474\
        );

    \I__5608\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23474\
        );

    \I__5607\ : InMux
    port map (
            O => \N__23530\,
            I => \N__23474\
        );

    \I__5606\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23474\
        );

    \I__5605\ : InMux
    port map (
            O => \N__23526\,
            I => \N__23474\
        );

    \I__5604\ : InMux
    port map (
            O => \N__23523\,
            I => \N__23474\
        );

    \I__5603\ : InMux
    port map (
            O => \N__23522\,
            I => \N__23474\
        );

    \I__5602\ : InMux
    port map (
            O => \N__23519\,
            I => \N__23474\
        );

    \I__5601\ : InMux
    port map (
            O => \N__23516\,
            I => \N__23471\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__23513\,
            I => \N__23467\
        );

    \I__5599\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23456\
        );

    \I__5598\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23456\
        );

    \I__5597\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23456\
        );

    \I__5596\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23456\
        );

    \I__5595\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23456\
        );

    \I__5594\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23453\
        );

    \I__5593\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23450\
        );

    \I__5592\ : Span4Mux_h
    port map (
            O => \N__23497\,
            I => \N__23447\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__23494\,
            I => \N__23444\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__23491\,
            I => \N__23441\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__23474\,
            I => \N__23438\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__23471\,
            I => \N__23435\
        );

    \I__5587\ : InMux
    port map (
            O => \N__23470\,
            I => \N__23432\
        );

    \I__5586\ : Span4Mux_v
    port map (
            O => \N__23467\,
            I => \N__23425\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__23456\,
            I => \N__23425\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__23453\,
            I => \N__23422\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23415\
        );

    \I__5582\ : Span4Mux_h
    port map (
            O => \N__23447\,
            I => \N__23415\
        );

    \I__5581\ : Span4Mux_h
    port map (
            O => \N__23444\,
            I => \N__23415\
        );

    \I__5580\ : Sp12to4
    port map (
            O => \N__23441\,
            I => \N__23408\
        );

    \I__5579\ : Span12Mux_h
    port map (
            O => \N__23438\,
            I => \N__23408\
        );

    \I__5578\ : Span12Mux_s2_h
    port map (
            O => \N__23435\,
            I => \N__23408\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__23432\,
            I => \N__23404\
        );

    \I__5576\ : InMux
    port map (
            O => \N__23431\,
            I => \N__23401\
        );

    \I__5575\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23398\
        );

    \I__5574\ : Span4Mux_v
    port map (
            O => \N__23425\,
            I => \N__23395\
        );

    \I__5573\ : Span12Mux_h
    port map (
            O => \N__23422\,
            I => \N__23392\
        );

    \I__5572\ : Span4Mux_v
    port map (
            O => \N__23415\,
            I => \N__23389\
        );

    \I__5571\ : Span12Mux_h
    port map (
            O => \N__23408\,
            I => \N__23386\
        );

    \I__5570\ : InMux
    port map (
            O => \N__23407\,
            I => \N__23383\
        );

    \I__5569\ : Span12Mux_v
    port map (
            O => \N__23404\,
            I => \N__23380\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__23401\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__23398\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5566\ : Odrv4
    port map (
            O => \N__23395\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5565\ : Odrv12
    port map (
            O => \N__23392\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5564\ : Odrv4
    port map (
            O => \N__23389\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5563\ : Odrv12
    port map (
            O => \N__23386\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__23383\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5561\ : Odrv12
    port map (
            O => \N__23380\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5560\ : IoInMux
    port map (
            O => \N__23363\,
            I => \N__23360\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__23360\,
            I => \N__23357\
        );

    \I__5558\ : IoSpan4Mux
    port map (
            O => \N__23357\,
            I => \N__23354\
        );

    \I__5557\ : Span4Mux_s1_v
    port map (
            O => \N__23354\,
            I => \N__23351\
        );

    \I__5556\ : Sp12to4
    port map (
            O => \N__23351\,
            I => \N__23348\
        );

    \I__5555\ : Span12Mux_h
    port map (
            O => \N__23348\,
            I => \N__23344\
        );

    \I__5554\ : InMux
    port map (
            O => \N__23347\,
            I => \N__23341\
        );

    \I__5553\ : Odrv12
    port map (
            O => \N__23344\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__23341\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__5551\ : IoInMux
    port map (
            O => \N__23336\,
            I => \N__23333\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__23333\,
            I => \N__23330\
        );

    \I__5549\ : Span12Mux_s9_v
    port map (
            O => \N__23330\,
            I => \N__23326\
        );

    \I__5548\ : InMux
    port map (
            O => \N__23329\,
            I => \N__23323\
        );

    \I__5547\ : Odrv12
    port map (
            O => \N__23326\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__23323\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__5545\ : InMux
    port map (
            O => \N__23318\,
            I => \un1_M_this_external_address_q_cry_0\
        );

    \I__5544\ : IoInMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__23312\,
            I => \N__23309\
        );

    \I__5542\ : Span4Mux_s3_v
    port map (
            O => \N__23309\,
            I => \N__23306\
        );

    \I__5541\ : Span4Mux_v
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__5540\ : Sp12to4
    port map (
            O => \N__23303\,
            I => \N__23300\
        );

    \I__5539\ : Span12Mux_h
    port map (
            O => \N__23300\,
            I => \N__23296\
        );

    \I__5538\ : InMux
    port map (
            O => \N__23299\,
            I => \N__23293\
        );

    \I__5537\ : Odrv12
    port map (
            O => \N__23296\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__23293\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__5535\ : InMux
    port map (
            O => \N__23288\,
            I => \un1_M_this_external_address_q_cry_1\
        );

    \I__5534\ : IoInMux
    port map (
            O => \N__23285\,
            I => \N__23282\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__23282\,
            I => \N__23279\
        );

    \I__5532\ : Span4Mux_s1_h
    port map (
            O => \N__23279\,
            I => \N__23276\
        );

    \I__5531\ : Span4Mux_v
    port map (
            O => \N__23276\,
            I => \N__23272\
        );

    \I__5530\ : InMux
    port map (
            O => \N__23275\,
            I => \N__23269\
        );

    \I__5529\ : Odrv4
    port map (
            O => \N__23272\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__23269\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__5527\ : InMux
    port map (
            O => \N__23264\,
            I => \un1_M_this_external_address_q_cry_2\
        );

    \I__5526\ : IoInMux
    port map (
            O => \N__23261\,
            I => \N__23258\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__23258\,
            I => \N__23254\
        );

    \I__5524\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23251\
        );

    \I__5523\ : Odrv4
    port map (
            O => \N__23254\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__23251\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__5521\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23243\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__23243\,
            I => \N__23240\
        );

    \I__5519\ : Span4Mux_v
    port map (
            O => \N__23240\,
            I => \N__23237\
        );

    \I__5518\ : Span4Mux_v
    port map (
            O => \N__23237\,
            I => \N__23234\
        );

    \I__5517\ : Span4Mux_v
    port map (
            O => \N__23234\,
            I => \N__23231\
        );

    \I__5516\ : Odrv4
    port map (
            O => \N__23231\,
            I => \this_sprites_ram.mem_out_bus7_3\
        );

    \I__5515\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23225\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__23225\,
            I => \N__23222\
        );

    \I__5513\ : Odrv4
    port map (
            O => \N__23222\,
            I => \this_sprites_ram.mem_out_bus3_3\
        );

    \I__5512\ : InMux
    port map (
            O => \N__23219\,
            I => \N__23216\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__23216\,
            I => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\
        );

    \I__5510\ : CEMux
    port map (
            O => \N__23213\,
            I => \N__23210\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__23210\,
            I => \N__23206\
        );

    \I__5508\ : CEMux
    port map (
            O => \N__23209\,
            I => \N__23203\
        );

    \I__5507\ : Odrv4
    port map (
            O => \N__23206\,
            I => \this_sprites_ram.mem_WE_6\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__23203\,
            I => \this_sprites_ram.mem_WE_6\
        );

    \I__5505\ : CascadeMux
    port map (
            O => \N__23198\,
            I => \N__23195\
        );

    \I__5504\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23189\
        );

    \I__5503\ : CascadeMux
    port map (
            O => \N__23194\,
            I => \N__23186\
        );

    \I__5502\ : InMux
    port map (
            O => \N__23193\,
            I => \N__23183\
        );

    \I__5501\ : InMux
    port map (
            O => \N__23192\,
            I => \N__23180\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__23189\,
            I => \N__23177\
        );

    \I__5499\ : InMux
    port map (
            O => \N__23186\,
            I => \N__23174\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__23183\,
            I => \N__23171\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__23180\,
            I => \N__23168\
        );

    \I__5496\ : Span4Mux_h
    port map (
            O => \N__23177\,
            I => \N__23163\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__23174\,
            I => \N__23163\
        );

    \I__5494\ : Span4Mux_h
    port map (
            O => \N__23171\,
            I => \N__23160\
        );

    \I__5493\ : Span4Mux_v
    port map (
            O => \N__23168\,
            I => \N__23157\
        );

    \I__5492\ : Sp12to4
    port map (
            O => \N__23163\,
            I => \N__23154\
        );

    \I__5491\ : Span4Mux_h
    port map (
            O => \N__23160\,
            I => \N__23151\
        );

    \I__5490\ : Span4Mux_h
    port map (
            O => \N__23157\,
            I => \N__23148\
        );

    \I__5489\ : Span12Mux_v
    port map (
            O => \N__23154\,
            I => \N__23145\
        );

    \I__5488\ : Sp12to4
    port map (
            O => \N__23151\,
            I => \N__23140\
        );

    \I__5487\ : Sp12to4
    port map (
            O => \N__23148\,
            I => \N__23140\
        );

    \I__5486\ : Span12Mux_h
    port map (
            O => \N__23145\,
            I => \N__23137\
        );

    \I__5485\ : Span12Mux_v
    port map (
            O => \N__23140\,
            I => \N__23134\
        );

    \I__5484\ : Odrv12
    port map (
            O => \N__23137\,
            I => port_data_c_3
        );

    \I__5483\ : Odrv12
    port map (
            O => \N__23134\,
            I => port_data_c_3
        );

    \I__5482\ : CascadeMux
    port map (
            O => \N__23129\,
            I => \N__23126\
        );

    \I__5481\ : InMux
    port map (
            O => \N__23126\,
            I => \N__23123\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__23123\,
            I => \N__23120\
        );

    \I__5479\ : Span4Mux_v
    port map (
            O => \N__23120\,
            I => \N__23117\
        );

    \I__5478\ : Span4Mux_h
    port map (
            O => \N__23117\,
            I => \N__23114\
        );

    \I__5477\ : IoSpan4Mux
    port map (
            O => \N__23114\,
            I => \N__23111\
        );

    \I__5476\ : Odrv4
    port map (
            O => \N__23111\,
            I => port_data_c_7
        );

    \I__5475\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23104\
        );

    \I__5474\ : InMux
    port map (
            O => \N__23107\,
            I => \N__23100\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__23104\,
            I => \N__23096\
        );

    \I__5472\ : InMux
    port map (
            O => \N__23103\,
            I => \N__23093\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__23100\,
            I => \N__23089\
        );

    \I__5470\ : InMux
    port map (
            O => \N__23099\,
            I => \N__23086\
        );

    \I__5469\ : Span4Mux_v
    port map (
            O => \N__23096\,
            I => \N__23080\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__23093\,
            I => \N__23080\
        );

    \I__5467\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23077\
        );

    \I__5466\ : Span4Mux_v
    port map (
            O => \N__23089\,
            I => \N__23071\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__23086\,
            I => \N__23071\
        );

    \I__5464\ : InMux
    port map (
            O => \N__23085\,
            I => \N__23068\
        );

    \I__5463\ : Span4Mux_v
    port map (
            O => \N__23080\,
            I => \N__23062\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__23077\,
            I => \N__23062\
        );

    \I__5461\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23059\
        );

    \I__5460\ : Span4Mux_v
    port map (
            O => \N__23071\,
            I => \N__23054\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__23068\,
            I => \N__23054\
        );

    \I__5458\ : InMux
    port map (
            O => \N__23067\,
            I => \N__23051\
        );

    \I__5457\ : Span4Mux_v
    port map (
            O => \N__23062\,
            I => \N__23046\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__23059\,
            I => \N__23046\
        );

    \I__5455\ : Span4Mux_v
    port map (
            O => \N__23054\,
            I => \N__23041\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__23051\,
            I => \N__23041\
        );

    \I__5453\ : Odrv4
    port map (
            O => \N__23046\,
            I => \M_this_sprites_ram_write_data_3\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__23041\,
            I => \M_this_sprites_ram_write_data_3\
        );

    \I__5451\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23033\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__23033\,
            I => \N__23030\
        );

    \I__5449\ : Span4Mux_v
    port map (
            O => \N__23030\,
            I => \N__23027\
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__23027\,
            I => \this_sprites_ram.mem_out_bus5_3\
        );

    \I__5447\ : InMux
    port map (
            O => \N__23024\,
            I => \N__23021\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__23021\,
            I => \N__23018\
        );

    \I__5445\ : Span4Mux_v
    port map (
            O => \N__23018\,
            I => \N__23015\
        );

    \I__5444\ : Span4Mux_v
    port map (
            O => \N__23015\,
            I => \N__23012\
        );

    \I__5443\ : Odrv4
    port map (
            O => \N__23012\,
            I => \this_sprites_ram.mem_out_bus1_3\
        );

    \I__5442\ : InMux
    port map (
            O => \N__23009\,
            I => \N__23006\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__23006\,
            I => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\
        );

    \I__5440\ : InMux
    port map (
            O => \N__23003\,
            I => \N__23000\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__23000\,
            I => \N__22997\
        );

    \I__5438\ : Sp12to4
    port map (
            O => \N__22997\,
            I => \N__22994\
        );

    \I__5437\ : Span12Mux_v
    port map (
            O => \N__22994\,
            I => \N__22991\
        );

    \I__5436\ : Odrv12
    port map (
            O => \N__22991\,
            I => \this_sprites_ram.mem_out_bus0_3\
        );

    \I__5435\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22985\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__22985\,
            I => \this_sprites_ram.mem_out_bus4_3\
        );

    \I__5433\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22979\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__22979\,
            I => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\
        );

    \I__5431\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22973\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__22973\,
            I => \N__22970\
        );

    \I__5429\ : Sp12to4
    port map (
            O => \N__22970\,
            I => \N__22967\
        );

    \I__5428\ : Odrv12
    port map (
            O => \N__22967\,
            I => \this_sprites_ram.mem_out_bus6_3\
        );

    \I__5427\ : InMux
    port map (
            O => \N__22964\,
            I => \N__22961\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__22961\,
            I => \N__22958\
        );

    \I__5425\ : Span4Mux_v
    port map (
            O => \N__22958\,
            I => \N__22955\
        );

    \I__5424\ : Span4Mux_v
    port map (
            O => \N__22955\,
            I => \N__22952\
        );

    \I__5423\ : Odrv4
    port map (
            O => \N__22952\,
            I => \this_sprites_ram.mem_out_bus2_3\
        );

    \I__5422\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22946\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__22946\,
            I => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\
        );

    \I__5420\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22940\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__22940\,
            I => \N__22937\
        );

    \I__5418\ : Span4Mux_v
    port map (
            O => \N__22937\,
            I => \N__22934\
        );

    \I__5417\ : Span4Mux_v
    port map (
            O => \N__22934\,
            I => \N__22931\
        );

    \I__5416\ : Odrv4
    port map (
            O => \N__22931\,
            I => \this_sprites_ram.mem_out_bus7_0\
        );

    \I__5415\ : InMux
    port map (
            O => \N__22928\,
            I => \N__22925\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__22925\,
            I => \N__22922\
        );

    \I__5413\ : Span4Mux_v
    port map (
            O => \N__22922\,
            I => \N__22919\
        );

    \I__5412\ : Odrv4
    port map (
            O => \N__22919\,
            I => \this_sprites_ram.mem_out_bus3_0\
        );

    \I__5411\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22911\
        );

    \I__5410\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22899\
        );

    \I__5409\ : InMux
    port map (
            O => \N__22914\,
            I => \N__22899\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__22911\,
            I => \N__22891\
        );

    \I__5407\ : InMux
    port map (
            O => \N__22910\,
            I => \N__22888\
        );

    \I__5406\ : InMux
    port map (
            O => \N__22909\,
            I => \N__22883\
        );

    \I__5405\ : InMux
    port map (
            O => \N__22908\,
            I => \N__22883\
        );

    \I__5404\ : InMux
    port map (
            O => \N__22907\,
            I => \N__22880\
        );

    \I__5403\ : InMux
    port map (
            O => \N__22906\,
            I => \N__22873\
        );

    \I__5402\ : InMux
    port map (
            O => \N__22905\,
            I => \N__22873\
        );

    \I__5401\ : InMux
    port map (
            O => \N__22904\,
            I => \N__22873\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__22899\,
            I => \N__22870\
        );

    \I__5399\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22867\
        );

    \I__5398\ : InMux
    port map (
            O => \N__22897\,
            I => \N__22862\
        );

    \I__5397\ : InMux
    port map (
            O => \N__22896\,
            I => \N__22862\
        );

    \I__5396\ : InMux
    port map (
            O => \N__22895\,
            I => \N__22859\
        );

    \I__5395\ : InMux
    port map (
            O => \N__22894\,
            I => \N__22856\
        );

    \I__5394\ : Span4Mux_v
    port map (
            O => \N__22891\,
            I => \N__22850\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__22888\,
            I => \N__22850\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__22883\,
            I => \N__22841\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__22880\,
            I => \N__22841\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__22873\,
            I => \N__22841\
        );

    \I__5389\ : Span4Mux_h
    port map (
            O => \N__22870\,
            I => \N__22841\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__22867\,
            I => \N__22832\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__22862\,
            I => \N__22832\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__22859\,
            I => \N__22832\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__22856\,
            I => \N__22832\
        );

    \I__5384\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22829\
        );

    \I__5383\ : Span4Mux_h
    port map (
            O => \N__22850\,
            I => \N__22826\
        );

    \I__5382\ : Span4Mux_v
    port map (
            O => \N__22841\,
            I => \N__22819\
        );

    \I__5381\ : Span4Mux_v
    port map (
            O => \N__22832\,
            I => \N__22819\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__22829\,
            I => \N__22819\
        );

    \I__5379\ : Span4Mux_v
    port map (
            O => \N__22826\,
            I => \N__22814\
        );

    \I__5378\ : Span4Mux_h
    port map (
            O => \N__22819\,
            I => \N__22814\
        );

    \I__5377\ : Odrv4
    port map (
            O => \N__22814\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__5376\ : InMux
    port map (
            O => \N__22811\,
            I => \N__22808\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__22808\,
            I => \N__22805\
        );

    \I__5374\ : Span12Mux_h
    port map (
            O => \N__22805\,
            I => \N__22802\
        );

    \I__5373\ : Odrv12
    port map (
            O => \N__22802\,
            I => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\
        );

    \I__5372\ : InMux
    port map (
            O => \N__22799\,
            I => \N__22796\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__22796\,
            I => \N__22792\
        );

    \I__5370\ : InMux
    port map (
            O => \N__22795\,
            I => \N__22789\
        );

    \I__5369\ : Span4Mux_v
    port map (
            O => \N__22792\,
            I => \N__22783\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__22789\,
            I => \N__22783\
        );

    \I__5367\ : InMux
    port map (
            O => \N__22788\,
            I => \N__22780\
        );

    \I__5366\ : Span4Mux_h
    port map (
            O => \N__22783\,
            I => \N__22774\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__22780\,
            I => \N__22774\
        );

    \I__5364\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22771\
        );

    \I__5363\ : Odrv4
    port map (
            O => \N__22774\,
            I => \this_vga_signals.N_481\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__22771\,
            I => \this_vga_signals.N_481\
        );

    \I__5361\ : CascadeMux
    port map (
            O => \N__22766\,
            I => \N__22763\
        );

    \I__5360\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22760\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__22760\,
            I => \N__22756\
        );

    \I__5358\ : CascadeMux
    port map (
            O => \N__22759\,
            I => \N__22751\
        );

    \I__5357\ : Span4Mux_h
    port map (
            O => \N__22756\,
            I => \N__22748\
        );

    \I__5356\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22745\
        );

    \I__5355\ : InMux
    port map (
            O => \N__22754\,
            I => \N__22740\
        );

    \I__5354\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22740\
        );

    \I__5353\ : Span4Mux_v
    port map (
            O => \N__22748\,
            I => \N__22735\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__22745\,
            I => \N__22735\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__22740\,
            I => \N__22732\
        );

    \I__5350\ : Span4Mux_v
    port map (
            O => \N__22735\,
            I => \N__22729\
        );

    \I__5349\ : Span12Mux_v
    port map (
            O => \N__22732\,
            I => \N__22726\
        );

    \I__5348\ : Sp12to4
    port map (
            O => \N__22729\,
            I => \N__22723\
        );

    \I__5347\ : Span12Mux_h
    port map (
            O => \N__22726\,
            I => \N__22720\
        );

    \I__5346\ : Span12Mux_h
    port map (
            O => \N__22723\,
            I => \N__22717\
        );

    \I__5345\ : Odrv12
    port map (
            O => \N__22720\,
            I => port_data_c_2
        );

    \I__5344\ : Odrv12
    port map (
            O => \N__22717\,
            I => port_data_c_2
        );

    \I__5343\ : CascadeMux
    port map (
            O => \N__22712\,
            I => \N__22708\
        );

    \I__5342\ : InMux
    port map (
            O => \N__22711\,
            I => \N__22703\
        );

    \I__5341\ : InMux
    port map (
            O => \N__22708\,
            I => \N__22703\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__22703\,
            I => \N__22700\
        );

    \I__5339\ : Span4Mux_v
    port map (
            O => \N__22700\,
            I => \N__22696\
        );

    \I__5338\ : CascadeMux
    port map (
            O => \N__22699\,
            I => \N__22693\
        );

    \I__5337\ : Span4Mux_h
    port map (
            O => \N__22696\,
            I => \N__22690\
        );

    \I__5336\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22687\
        );

    \I__5335\ : Sp12to4
    port map (
            O => \N__22690\,
            I => \N__22682\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__22687\,
            I => \N__22682\
        );

    \I__5333\ : Span12Mux_v
    port map (
            O => \N__22682\,
            I => \N__22679\
        );

    \I__5332\ : Odrv12
    port map (
            O => \N__22679\,
            I => port_data_c_6
        );

    \I__5331\ : CEMux
    port map (
            O => \N__22676\,
            I => \N__22672\
        );

    \I__5330\ : CEMux
    port map (
            O => \N__22675\,
            I => \N__22669\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__22672\,
            I => \N__22664\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__22669\,
            I => \N__22664\
        );

    \I__5327\ : Odrv4
    port map (
            O => \N__22664\,
            I => \this_sprites_ram.mem_WE_10\
        );

    \I__5326\ : CEMux
    port map (
            O => \N__22661\,
            I => \N__22657\
        );

    \I__5325\ : CEMux
    port map (
            O => \N__22660\,
            I => \N__22654\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__22657\,
            I => \N__22651\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__22654\,
            I => \N__22648\
        );

    \I__5322\ : Span4Mux_v
    port map (
            O => \N__22651\,
            I => \N__22645\
        );

    \I__5321\ : Span4Mux_h
    port map (
            O => \N__22648\,
            I => \N__22642\
        );

    \I__5320\ : Odrv4
    port map (
            O => \N__22645\,
            I => \this_sprites_ram.mem_WE_12\
        );

    \I__5319\ : Odrv4
    port map (
            O => \N__22642\,
            I => \this_sprites_ram.mem_WE_12\
        );

    \I__5318\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22634\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__22634\,
            I => \N__22631\
        );

    \I__5316\ : Span4Mux_v
    port map (
            O => \N__22631\,
            I => \N__22628\
        );

    \I__5315\ : Sp12to4
    port map (
            O => \N__22628\,
            I => \N__22625\
        );

    \I__5314\ : Odrv12
    port map (
            O => \N__22625\,
            I => \this_sprites_ram.mem_out_bus5_2\
        );

    \I__5313\ : InMux
    port map (
            O => \N__22622\,
            I => \N__22619\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__22619\,
            I => \N__22616\
        );

    \I__5311\ : Span4Mux_v
    port map (
            O => \N__22616\,
            I => \N__22613\
        );

    \I__5310\ : Odrv4
    port map (
            O => \N__22613\,
            I => \this_sprites_ram.mem_out_bus1_2\
        );

    \I__5309\ : InMux
    port map (
            O => \N__22610\,
            I => \N__22607\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__22607\,
            I => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\
        );

    \I__5307\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22601\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22598\
        );

    \I__5305\ : Span4Mux_h
    port map (
            O => \N__22598\,
            I => \N__22595\
        );

    \I__5304\ : Odrv4
    port map (
            O => \N__22595\,
            I => \this_sprites_ram.mem_out_bus4_1\
        );

    \I__5303\ : InMux
    port map (
            O => \N__22592\,
            I => \N__22589\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__22589\,
            I => \N__22586\
        );

    \I__5301\ : Sp12to4
    port map (
            O => \N__22586\,
            I => \N__22583\
        );

    \I__5300\ : Span12Mux_v
    port map (
            O => \N__22583\,
            I => \N__22580\
        );

    \I__5299\ : Odrv12
    port map (
            O => \N__22580\,
            I => \this_sprites_ram.mem_out_bus0_1\
        );

    \I__5298\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22574\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__22574\,
            I => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0\
        );

    \I__5296\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22568\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__5294\ : Span4Mux_v
    port map (
            O => \N__22565\,
            I => \N__22562\
        );

    \I__5293\ : Odrv4
    port map (
            O => \N__22562\,
            I => \this_sprites_ram.mem_out_bus4_2\
        );

    \I__5292\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22556\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__22556\,
            I => \N__22553\
        );

    \I__5290\ : Span4Mux_v
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__5289\ : Span4Mux_v
    port map (
            O => \N__22550\,
            I => \N__22547\
        );

    \I__5288\ : Odrv4
    port map (
            O => \N__22547\,
            I => \this_sprites_ram.mem_out_bus0_2\
        );

    \I__5287\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22541\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__22541\,
            I => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0\
        );

    \I__5285\ : CEMux
    port map (
            O => \N__22538\,
            I => \N__22534\
        );

    \I__5284\ : CEMux
    port map (
            O => \N__22537\,
            I => \N__22531\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__22534\,
            I => \N__22528\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__22531\,
            I => \N__22525\
        );

    \I__5281\ : Span4Mux_v
    port map (
            O => \N__22528\,
            I => \N__22522\
        );

    \I__5280\ : Span4Mux_h
    port map (
            O => \N__22525\,
            I => \N__22519\
        );

    \I__5279\ : Odrv4
    port map (
            O => \N__22522\,
            I => \this_sprites_ram.mem_WE_8\
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__22519\,
            I => \this_sprites_ram.mem_WE_8\
        );

    \I__5277\ : InMux
    port map (
            O => \N__22514\,
            I => \N__22511\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__22511\,
            I => \N__22508\
        );

    \I__5275\ : Sp12to4
    port map (
            O => \N__22508\,
            I => \N__22505\
        );

    \I__5274\ : Span12Mux_v
    port map (
            O => \N__22505\,
            I => \N__22502\
        );

    \I__5273\ : Span12Mux_v
    port map (
            O => \N__22502\,
            I => \N__22499\
        );

    \I__5272\ : Odrv12
    port map (
            O => \N__22499\,
            I => \this_sprites_ram.mem_out_bus7_2\
        );

    \I__5271\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22493\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__22493\,
            I => \N__22490\
        );

    \I__5269\ : Span4Mux_h
    port map (
            O => \N__22490\,
            I => \N__22487\
        );

    \I__5268\ : Odrv4
    port map (
            O => \N__22487\,
            I => \this_sprites_ram.mem_out_bus3_2\
        );

    \I__5267\ : InMux
    port map (
            O => \N__22484\,
            I => \N__22481\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__22481\,
            I => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\
        );

    \I__5265\ : InMux
    port map (
            O => \N__22478\,
            I => \N__22475\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__22475\,
            I => \N__22472\
        );

    \I__5263\ : Span4Mux_v
    port map (
            O => \N__22472\,
            I => \N__22469\
        );

    \I__5262\ : Span4Mux_v
    port map (
            O => \N__22469\,
            I => \N__22466\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__22466\,
            I => \N__22463\
        );

    \I__5260\ : Odrv4
    port map (
            O => \N__22463\,
            I => \this_sprites_ram.mem_out_bus7_1\
        );

    \I__5259\ : InMux
    port map (
            O => \N__22460\,
            I => \N__22457\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__22457\,
            I => \this_sprites_ram.mem_out_bus3_1\
        );

    \I__5257\ : InMux
    port map (
            O => \N__22454\,
            I => \N__22451\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__22451\,
            I => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\
        );

    \I__5255\ : InMux
    port map (
            O => \N__22448\,
            I => \N__22445\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__22445\,
            I => \N__22442\
        );

    \I__5253\ : Span4Mux_v
    port map (
            O => \N__22442\,
            I => \N__22439\
        );

    \I__5252\ : Span4Mux_v
    port map (
            O => \N__22439\,
            I => \N__22436\
        );

    \I__5251\ : Odrv4
    port map (
            O => \N__22436\,
            I => \this_sprites_ram.mem_out_bus6_1\
        );

    \I__5250\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22430\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__22430\,
            I => \N__22427\
        );

    \I__5248\ : Span4Mux_v
    port map (
            O => \N__22427\,
            I => \N__22424\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__22424\,
            I => \this_sprites_ram.mem_out_bus2_1\
        );

    \I__5246\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22418\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__22418\,
            I => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\
        );

    \I__5244\ : CascadeMux
    port map (
            O => \N__22415\,
            I => \M_this_sprites_ram_read_data_3_cascade_\
        );

    \I__5243\ : InMux
    port map (
            O => \N__22412\,
            I => \N__22408\
        );

    \I__5242\ : InMux
    port map (
            O => \N__22411\,
            I => \N__22405\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__22408\,
            I => \N__22401\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__22405\,
            I => \N__22398\
        );

    \I__5239\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22395\
        );

    \I__5238\ : Span4Mux_h
    port map (
            O => \N__22401\,
            I => \N__22392\
        );

    \I__5237\ : Span4Mux_h
    port map (
            O => \N__22398\,
            I => \N__22387\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__22395\,
            I => \N__22387\
        );

    \I__5235\ : Span4Mux_h
    port map (
            O => \N__22392\,
            I => \N__22379\
        );

    \I__5234\ : Span4Mux_v
    port map (
            O => \N__22387\,
            I => \N__22379\
        );

    \I__5233\ : InMux
    port map (
            O => \N__22386\,
            I => \N__22375\
        );

    \I__5232\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22372\
        );

    \I__5231\ : InMux
    port map (
            O => \N__22384\,
            I => \N__22369\
        );

    \I__5230\ : Span4Mux_h
    port map (
            O => \N__22379\,
            I => \N__22366\
        );

    \I__5229\ : CascadeMux
    port map (
            O => \N__22378\,
            I => \N__22360\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__22375\,
            I => \N__22357\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__22372\,
            I => \N__22354\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__22369\,
            I => \N__22351\
        );

    \I__5225\ : Span4Mux_h
    port map (
            O => \N__22366\,
            I => \N__22348\
        );

    \I__5224\ : InMux
    port map (
            O => \N__22365\,
            I => \N__22341\
        );

    \I__5223\ : InMux
    port map (
            O => \N__22364\,
            I => \N__22341\
        );

    \I__5222\ : InMux
    port map (
            O => \N__22363\,
            I => \N__22341\
        );

    \I__5221\ : InMux
    port map (
            O => \N__22360\,
            I => \N__22338\
        );

    \I__5220\ : Span4Mux_h
    port map (
            O => \N__22357\,
            I => \N__22331\
        );

    \I__5219\ : Span4Mux_v
    port map (
            O => \N__22354\,
            I => \N__22331\
        );

    \I__5218\ : Span4Mux_h
    port map (
            O => \N__22351\,
            I => \N__22331\
        );

    \I__5217\ : Odrv4
    port map (
            O => \N__22348\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__22341\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__22338\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__5214\ : Odrv4
    port map (
            O => \N__22331\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__5213\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__22319\,
            I => \N__22316\
        );

    \I__5211\ : Span4Mux_v
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__5210\ : Span4Mux_h
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__5209\ : Sp12to4
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__5208\ : Span12Mux_h
    port map (
            O => \N__22307\,
            I => \N__22304\
        );

    \I__5207\ : Odrv12
    port map (
            O => \N__22304\,
            I => \M_this_vram_write_data_3\
        );

    \I__5206\ : CascadeMux
    port map (
            O => \N__22301\,
            I => \N__22295\
        );

    \I__5205\ : CascadeMux
    port map (
            O => \N__22300\,
            I => \N__22292\
        );

    \I__5204\ : InMux
    port map (
            O => \N__22299\,
            I => \N__22289\
        );

    \I__5203\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22286\
        );

    \I__5202\ : InMux
    port map (
            O => \N__22295\,
            I => \N__22282\
        );

    \I__5201\ : InMux
    port map (
            O => \N__22292\,
            I => \N__22279\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__22289\,
            I => \N__22274\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__22286\,
            I => \N__22274\
        );

    \I__5198\ : InMux
    port map (
            O => \N__22285\,
            I => \N__22271\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__22282\,
            I => \N__22265\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__22279\,
            I => \N__22260\
        );

    \I__5195\ : Span4Mux_h
    port map (
            O => \N__22274\,
            I => \N__22260\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__22271\,
            I => \N__22257\
        );

    \I__5193\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22254\
        );

    \I__5192\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22251\
        );

    \I__5191\ : InMux
    port map (
            O => \N__22268\,
            I => \N__22248\
        );

    \I__5190\ : Span4Mux_v
    port map (
            O => \N__22265\,
            I => \N__22245\
        );

    \I__5189\ : Span4Mux_v
    port map (
            O => \N__22260\,
            I => \N__22238\
        );

    \I__5188\ : Span4Mux_h
    port map (
            O => \N__22257\,
            I => \N__22238\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__22254\,
            I => \N__22238\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__22251\,
            I => \N__22233\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__22248\,
            I => \N__22233\
        );

    \I__5184\ : Span4Mux_h
    port map (
            O => \N__22245\,
            I => \N__22228\
        );

    \I__5183\ : Span4Mux_h
    port map (
            O => \N__22238\,
            I => \N__22228\
        );

    \I__5182\ : Span12Mux_h
    port map (
            O => \N__22233\,
            I => \N__22225\
        );

    \I__5181\ : Span4Mux_h
    port map (
            O => \N__22228\,
            I => \N__22222\
        );

    \I__5180\ : Odrv12
    port map (
            O => \N__22225\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__22222\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__5178\ : CascadeMux
    port map (
            O => \N__22217\,
            I => \N__22214\
        );

    \I__5177\ : InMux
    port map (
            O => \N__22214\,
            I => \N__22208\
        );

    \I__5176\ : CascadeMux
    port map (
            O => \N__22213\,
            I => \N__22205\
        );

    \I__5175\ : CascadeMux
    port map (
            O => \N__22212\,
            I => \N__22202\
        );

    \I__5174\ : InMux
    port map (
            O => \N__22211\,
            I => \N__22199\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__22208\,
            I => \N__22196\
        );

    \I__5172\ : InMux
    port map (
            O => \N__22205\,
            I => \N__22193\
        );

    \I__5171\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22190\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__22199\,
            I => \N__22187\
        );

    \I__5169\ : Span4Mux_v
    port map (
            O => \N__22196\,
            I => \N__22182\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__22193\,
            I => \N__22182\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__22190\,
            I => \N__22179\
        );

    \I__5166\ : Span4Mux_h
    port map (
            O => \N__22187\,
            I => \N__22176\
        );

    \I__5165\ : Span4Mux_v
    port map (
            O => \N__22182\,
            I => \N__22173\
        );

    \I__5164\ : Span4Mux_v
    port map (
            O => \N__22179\,
            I => \N__22170\
        );

    \I__5163\ : Span4Mux_v
    port map (
            O => \N__22176\,
            I => \N__22165\
        );

    \I__5162\ : Span4Mux_h
    port map (
            O => \N__22173\,
            I => \N__22165\
        );

    \I__5161\ : Span4Mux_h
    port map (
            O => \N__22170\,
            I => \N__22162\
        );

    \I__5160\ : Odrv4
    port map (
            O => \N__22165\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__5159\ : Odrv4
    port map (
            O => \N__22162\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__5158\ : InMux
    port map (
            O => \N__22157\,
            I => \N__22154\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__22154\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3\
        );

    \I__5156\ : InMux
    port map (
            O => \N__22151\,
            I => \N__22148\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__22148\,
            I => \N__22145\
        );

    \I__5154\ : Span12Mux_h
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__5153\ : Odrv12
    port map (
            O => \N__22142\,
            I => \this_sprites_ram.mem_out_bus6_0\
        );

    \I__5152\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22136\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__22136\,
            I => \N__22133\
        );

    \I__5150\ : Span4Mux_v
    port map (
            O => \N__22133\,
            I => \N__22130\
        );

    \I__5149\ : Span4Mux_v
    port map (
            O => \N__22130\,
            I => \N__22127\
        );

    \I__5148\ : Odrv4
    port map (
            O => \N__22127\,
            I => \this_sprites_ram.mem_out_bus2_0\
        );

    \I__5147\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22121\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__22121\,
            I => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\
        );

    \I__5145\ : InMux
    port map (
            O => \N__22118\,
            I => \N__22115\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__22115\,
            I => \N__22112\
        );

    \I__5143\ : Span4Mux_v
    port map (
            O => \N__22112\,
            I => \N__22109\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__22109\,
            I => \this_sprites_ram.mem_out_bus5_0\
        );

    \I__5141\ : InMux
    port map (
            O => \N__22106\,
            I => \N__22103\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__22103\,
            I => \N__22100\
        );

    \I__5139\ : Span4Mux_v
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__5138\ : Span4Mux_v
    port map (
            O => \N__22097\,
            I => \N__22094\
        );

    \I__5137\ : Span4Mux_v
    port map (
            O => \N__22094\,
            I => \N__22091\
        );

    \I__5136\ : Span4Mux_v
    port map (
            O => \N__22091\,
            I => \N__22088\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__22088\,
            I => \this_sprites_ram.mem_out_bus1_0\
        );

    \I__5134\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22082\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__22082\,
            I => \N__22079\
        );

    \I__5132\ : Span12Mux_h
    port map (
            O => \N__22079\,
            I => \N__22076\
        );

    \I__5131\ : Odrv12
    port map (
            O => \N__22076\,
            I => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\
        );

    \I__5130\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22069\
        );

    \I__5129\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22066\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__22069\,
            I => \N__22063\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__22066\,
            I => \N__22060\
        );

    \I__5126\ : Odrv12
    port map (
            O => \N__22063\,
            I => \this_vga_signals.N_483\
        );

    \I__5125\ : Odrv4
    port map (
            O => \N__22060\,
            I => \this_vga_signals.N_483\
        );

    \I__5124\ : InMux
    port map (
            O => \N__22055\,
            I => \N__22049\
        );

    \I__5123\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22046\
        );

    \I__5122\ : InMux
    port map (
            O => \N__22053\,
            I => \N__22037\
        );

    \I__5121\ : InMux
    port map (
            O => \N__22052\,
            I => \N__22032\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__22049\,
            I => \N__22023\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__22046\,
            I => \N__22018\
        );

    \I__5118\ : InMux
    port map (
            O => \N__22045\,
            I => \N__22011\
        );

    \I__5117\ : InMux
    port map (
            O => \N__22044\,
            I => \N__22011\
        );

    \I__5116\ : InMux
    port map (
            O => \N__22043\,
            I => \N__22011\
        );

    \I__5115\ : InMux
    port map (
            O => \N__22042\,
            I => \N__22004\
        );

    \I__5114\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22004\
        );

    \I__5113\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22004\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__22037\,
            I => \N__22000\
        );

    \I__5111\ : InMux
    port map (
            O => \N__22036\,
            I => \N__21995\
        );

    \I__5110\ : InMux
    port map (
            O => \N__22035\,
            I => \N__21995\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__22032\,
            I => \N__21992\
        );

    \I__5108\ : InMux
    port map (
            O => \N__22031\,
            I => \N__21989\
        );

    \I__5107\ : InMux
    port map (
            O => \N__22030\,
            I => \N__21986\
        );

    \I__5106\ : InMux
    port map (
            O => \N__22029\,
            I => \N__21983\
        );

    \I__5105\ : InMux
    port map (
            O => \N__22028\,
            I => \N__21978\
        );

    \I__5104\ : InMux
    port map (
            O => \N__22027\,
            I => \N__21978\
        );

    \I__5103\ : InMux
    port map (
            O => \N__22026\,
            I => \N__21972\
        );

    \I__5102\ : Span4Mux_v
    port map (
            O => \N__22023\,
            I => \N__21969\
        );

    \I__5101\ : InMux
    port map (
            O => \N__22022\,
            I => \N__21966\
        );

    \I__5100\ : InMux
    port map (
            O => \N__22021\,
            I => \N__21963\
        );

    \I__5099\ : Span4Mux_v
    port map (
            O => \N__22018\,
            I => \N__21956\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__22011\,
            I => \N__21956\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__22004\,
            I => \N__21956\
        );

    \I__5096\ : InMux
    port map (
            O => \N__22003\,
            I => \N__21953\
        );

    \I__5095\ : Sp12to4
    port map (
            O => \N__22000\,
            I => \N__21948\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__21995\,
            I => \N__21948\
        );

    \I__5093\ : Span4Mux_v
    port map (
            O => \N__21992\,
            I => \N__21939\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__21989\,
            I => \N__21939\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__21986\,
            I => \N__21939\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__21983\,
            I => \N__21939\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__21978\,
            I => \N__21936\
        );

    \I__5088\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21929\
        );

    \I__5087\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21929\
        );

    \I__5086\ : InMux
    port map (
            O => \N__21975\,
            I => \N__21929\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__21972\,
            I => \N__21922\
        );

    \I__5084\ : Sp12to4
    port map (
            O => \N__21969\,
            I => \N__21922\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__21966\,
            I => \N__21922\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__21963\,
            I => \N__21917\
        );

    \I__5081\ : Span4Mux_h
    port map (
            O => \N__21956\,
            I => \N__21917\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__21953\,
            I => \N__21912\
        );

    \I__5079\ : Span12Mux_v
    port map (
            O => \N__21948\,
            I => \N__21912\
        );

    \I__5078\ : Span4Mux_h
    port map (
            O => \N__21939\,
            I => \N__21905\
        );

    \I__5077\ : Span4Mux_v
    port map (
            O => \N__21936\,
            I => \N__21905\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__21929\,
            I => \N__21905\
        );

    \I__5075\ : Span12Mux_h
    port map (
            O => \N__21922\,
            I => \N__21902\
        );

    \I__5074\ : Span4Mux_h
    port map (
            O => \N__21917\,
            I => \N__21899\
        );

    \I__5073\ : Odrv12
    port map (
            O => \N__21912\,
            I => \N_175_0\
        );

    \I__5072\ : Odrv4
    port map (
            O => \N__21905\,
            I => \N_175_0\
        );

    \I__5071\ : Odrv12
    port map (
            O => \N__21902\,
            I => \N_175_0\
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__21899\,
            I => \N_175_0\
        );

    \I__5069\ : CEMux
    port map (
            O => \N__21890\,
            I => \N__21887\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__21887\,
            I => \N__21883\
        );

    \I__5067\ : CEMux
    port map (
            O => \N__21886\,
            I => \N__21880\
        );

    \I__5066\ : Span4Mux_s2_v
    port map (
            O => \N__21883\,
            I => \N__21875\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__21880\,
            I => \N__21875\
        );

    \I__5064\ : Span4Mux_v
    port map (
            O => \N__21875\,
            I => \N__21872\
        );

    \I__5063\ : Span4Mux_v
    port map (
            O => \N__21872\,
            I => \N__21869\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__21869\,
            I => \this_sprites_ram.mem_WE_0\
        );

    \I__5061\ : CEMux
    port map (
            O => \N__21866\,
            I => \N__21862\
        );

    \I__5060\ : CEMux
    port map (
            O => \N__21865\,
            I => \N__21859\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__21862\,
            I => \N__21856\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__21859\,
            I => \N__21853\
        );

    \I__5057\ : Span4Mux_s3_v
    port map (
            O => \N__21856\,
            I => \N__21850\
        );

    \I__5056\ : Span4Mux_h
    port map (
            O => \N__21853\,
            I => \N__21847\
        );

    \I__5055\ : Span4Mux_v
    port map (
            O => \N__21850\,
            I => \N__21844\
        );

    \I__5054\ : Span4Mux_v
    port map (
            O => \N__21847\,
            I => \N__21841\
        );

    \I__5053\ : Odrv4
    port map (
            O => \N__21844\,
            I => \this_sprites_ram.mem_WE_14\
        );

    \I__5052\ : Odrv4
    port map (
            O => \N__21841\,
            I => \this_sprites_ram.mem_WE_14\
        );

    \I__5051\ : InMux
    port map (
            O => \N__21836\,
            I => \N__21833\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__21833\,
            I => \N__21830\
        );

    \I__5049\ : Span4Mux_v
    port map (
            O => \N__21830\,
            I => \N__21827\
        );

    \I__5048\ : Span4Mux_h
    port map (
            O => \N__21827\,
            I => \N__21824\
        );

    \I__5047\ : Sp12to4
    port map (
            O => \N__21824\,
            I => \N__21821\
        );

    \I__5046\ : Odrv12
    port map (
            O => \N__21821\,
            I => \M_this_vram_write_data_2\
        );

    \I__5045\ : InMux
    port map (
            O => \N__21818\,
            I => \N__21815\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__21815\,
            I => \N__21812\
        );

    \I__5043\ : Span4Mux_v
    port map (
            O => \N__21812\,
            I => \N__21809\
        );

    \I__5042\ : Span4Mux_h
    port map (
            O => \N__21809\,
            I => \N__21806\
        );

    \I__5041\ : Span4Mux_h
    port map (
            O => \N__21806\,
            I => \N__21803\
        );

    \I__5040\ : Odrv4
    port map (
            O => \N__21803\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0\
        );

    \I__5039\ : InMux
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__5037\ : Span4Mux_v
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__5036\ : Span4Mux_v
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__5035\ : Span4Mux_v
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__5034\ : Span4Mux_v
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__5033\ : Odrv4
    port map (
            O => \N__21782\,
            I => \this_sprites_ram.mem_out_bus6_2\
        );

    \I__5032\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__5030\ : Span4Mux_v
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__5029\ : Odrv4
    port map (
            O => \N__21770\,
            I => \this_sprites_ram.mem_out_bus2_2\
        );

    \I__5028\ : CascadeMux
    port map (
            O => \N__21767\,
            I => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0_cascade_\
        );

    \I__5027\ : CascadeMux
    port map (
            O => \N__21764\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\
        );

    \I__5026\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__21758\,
            I => \M_this_sprites_ram_read_data_2\
        );

    \I__5024\ : CascadeMux
    port map (
            O => \N__21755\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\
        );

    \I__5023\ : InMux
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__21749\,
            I => \N__21746\
        );

    \I__5021\ : Odrv12
    port map (
            O => \N__21746\,
            I => \M_this_sprites_ram_read_data_1\
        );

    \I__5020\ : InMux
    port map (
            O => \N__21743\,
            I => \N__21740\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__5018\ : Span4Mux_v
    port map (
            O => \N__21737\,
            I => \N__21734\
        );

    \I__5017\ : Span4Mux_v
    port map (
            O => \N__21734\,
            I => \N__21731\
        );

    \I__5016\ : Odrv4
    port map (
            O => \N__21731\,
            I => \this_sprites_ram.mem_out_bus5_1\
        );

    \I__5015\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21725\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__5013\ : Span4Mux_v
    port map (
            O => \N__21722\,
            I => \N__21719\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__21719\,
            I => \N__21716\
        );

    \I__5011\ : Span4Mux_v
    port map (
            O => \N__21716\,
            I => \N__21713\
        );

    \I__5010\ : Odrv4
    port map (
            O => \N__21713\,
            I => \this_sprites_ram.mem_out_bus1_1\
        );

    \I__5009\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21707\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__21707\,
            I => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\
        );

    \I__5007\ : InMux
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__21701\,
            I => \N__21698\
        );

    \I__5005\ : Span4Mux_h
    port map (
            O => \N__21698\,
            I => \N__21695\
        );

    \I__5004\ : Odrv4
    port map (
            O => \N__21695\,
            I => \this_sprites_ram.mem_out_bus4_0\
        );

    \I__5003\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21689\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__21689\,
            I => \N__21686\
        );

    \I__5001\ : Span4Mux_h
    port map (
            O => \N__21686\,
            I => \N__21683\
        );

    \I__5000\ : Span4Mux_v
    port map (
            O => \N__21683\,
            I => \N__21680\
        );

    \I__4999\ : Span4Mux_v
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__4998\ : Span4Mux_v
    port map (
            O => \N__21677\,
            I => \N__21674\
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__21674\,
            I => \this_sprites_ram.mem_out_bus0_0\
        );

    \I__4996\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21668\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__21668\,
            I => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0\
        );

    \I__4994\ : CascadeMux
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__4993\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21653\
        );

    \I__4992\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21653\
        );

    \I__4991\ : InMux
    port map (
            O => \N__21660\,
            I => \N__21653\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__21653\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__4989\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21646\
        );

    \I__4988\ : InMux
    port map (
            O => \N__21649\,
            I => \N__21643\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__21646\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__21643\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__21638\,
            I => \N__21630\
        );

    \I__4984\ : CascadeMux
    port map (
            O => \N__21637\,
            I => \N__21627\
        );

    \I__4983\ : CascadeMux
    port map (
            O => \N__21636\,
            I => \N__21622\
        );

    \I__4982\ : CascadeMux
    port map (
            O => \N__21635\,
            I => \N__21619\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__21634\,
            I => \N__21616\
        );

    \I__4980\ : CascadeMux
    port map (
            O => \N__21633\,
            I => \N__21613\
        );

    \I__4979\ : InMux
    port map (
            O => \N__21630\,
            I => \N__21609\
        );

    \I__4978\ : InMux
    port map (
            O => \N__21627\,
            I => \N__21606\
        );

    \I__4977\ : CascadeMux
    port map (
            O => \N__21626\,
            I => \N__21603\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__21625\,
            I => \N__21598\
        );

    \I__4975\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21595\
        );

    \I__4974\ : InMux
    port map (
            O => \N__21619\,
            I => \N__21592\
        );

    \I__4973\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21587\
        );

    \I__4972\ : InMux
    port map (
            O => \N__21613\,
            I => \N__21587\
        );

    \I__4971\ : CascadeMux
    port map (
            O => \N__21612\,
            I => \N__21584\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__21609\,
            I => \N__21580\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__21606\,
            I => \N__21577\
        );

    \I__4968\ : InMux
    port map (
            O => \N__21603\,
            I => \N__21572\
        );

    \I__4967\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21572\
        );

    \I__4966\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21567\
        );

    \I__4965\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21567\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__21595\,
            I => \N__21563\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__21592\,
            I => \N__21560\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__21587\,
            I => \N__21557\
        );

    \I__4961\ : InMux
    port map (
            O => \N__21584\,
            I => \N__21554\
        );

    \I__4960\ : InMux
    port map (
            O => \N__21583\,
            I => \N__21551\
        );

    \I__4959\ : Span4Mux_v
    port map (
            O => \N__21580\,
            I => \N__21542\
        );

    \I__4958\ : Span4Mux_h
    port map (
            O => \N__21577\,
            I => \N__21542\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__21572\,
            I => \N__21542\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__21567\,
            I => \N__21542\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__21566\,
            I => \N__21538\
        );

    \I__4954\ : Span4Mux_h
    port map (
            O => \N__21563\,
            I => \N__21535\
        );

    \I__4953\ : Span4Mux_v
    port map (
            O => \N__21560\,
            I => \N__21528\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__21557\,
            I => \N__21528\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__21554\,
            I => \N__21528\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__21551\,
            I => \N__21525\
        );

    \I__4949\ : Span4Mux_h
    port map (
            O => \N__21542\,
            I => \N__21522\
        );

    \I__4948\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21517\
        );

    \I__4947\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21517\
        );

    \I__4946\ : Odrv4
    port map (
            O => \N__21535\,
            I => \N_14_0\
        );

    \I__4945\ : Odrv4
    port map (
            O => \N__21528\,
            I => \N_14_0\
        );

    \I__4944\ : Odrv4
    port map (
            O => \N__21525\,
            I => \N_14_0\
        );

    \I__4943\ : Odrv4
    port map (
            O => \N__21522\,
            I => \N_14_0\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__21517\,
            I => \N_14_0\
        );

    \I__4941\ : CascadeMux
    port map (
            O => \N__21506\,
            I => \N__21503\
        );

    \I__4940\ : CascadeBuf
    port map (
            O => \N__21503\,
            I => \N__21500\
        );

    \I__4939\ : CascadeMux
    port map (
            O => \N__21500\,
            I => \N__21497\
        );

    \I__4938\ : CascadeBuf
    port map (
            O => \N__21497\,
            I => \N__21494\
        );

    \I__4937\ : CascadeMux
    port map (
            O => \N__21494\,
            I => \N__21491\
        );

    \I__4936\ : CascadeBuf
    port map (
            O => \N__21491\,
            I => \N__21488\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__21488\,
            I => \N__21485\
        );

    \I__4934\ : CascadeBuf
    port map (
            O => \N__21485\,
            I => \N__21482\
        );

    \I__4933\ : CascadeMux
    port map (
            O => \N__21482\,
            I => \N__21479\
        );

    \I__4932\ : CascadeBuf
    port map (
            O => \N__21479\,
            I => \N__21476\
        );

    \I__4931\ : CascadeMux
    port map (
            O => \N__21476\,
            I => \N__21473\
        );

    \I__4930\ : CascadeBuf
    port map (
            O => \N__21473\,
            I => \N__21470\
        );

    \I__4929\ : CascadeMux
    port map (
            O => \N__21470\,
            I => \N__21467\
        );

    \I__4928\ : CascadeBuf
    port map (
            O => \N__21467\,
            I => \N__21464\
        );

    \I__4927\ : CascadeMux
    port map (
            O => \N__21464\,
            I => \N__21461\
        );

    \I__4926\ : CascadeBuf
    port map (
            O => \N__21461\,
            I => \N__21458\
        );

    \I__4925\ : CascadeMux
    port map (
            O => \N__21458\,
            I => \N__21455\
        );

    \I__4924\ : CascadeBuf
    port map (
            O => \N__21455\,
            I => \N__21452\
        );

    \I__4923\ : CascadeMux
    port map (
            O => \N__21452\,
            I => \N__21449\
        );

    \I__4922\ : CascadeBuf
    port map (
            O => \N__21449\,
            I => \N__21446\
        );

    \I__4921\ : CascadeMux
    port map (
            O => \N__21446\,
            I => \N__21443\
        );

    \I__4920\ : CascadeBuf
    port map (
            O => \N__21443\,
            I => \N__21440\
        );

    \I__4919\ : CascadeMux
    port map (
            O => \N__21440\,
            I => \N__21437\
        );

    \I__4918\ : CascadeBuf
    port map (
            O => \N__21437\,
            I => \N__21434\
        );

    \I__4917\ : CascadeMux
    port map (
            O => \N__21434\,
            I => \N__21431\
        );

    \I__4916\ : CascadeBuf
    port map (
            O => \N__21431\,
            I => \N__21428\
        );

    \I__4915\ : CascadeMux
    port map (
            O => \N__21428\,
            I => \N__21425\
        );

    \I__4914\ : CascadeBuf
    port map (
            O => \N__21425\,
            I => \N__21422\
        );

    \I__4913\ : CascadeMux
    port map (
            O => \N__21422\,
            I => \N__21419\
        );

    \I__4912\ : CascadeBuf
    port map (
            O => \N__21419\,
            I => \N__21416\
        );

    \I__4911\ : CascadeMux
    port map (
            O => \N__21416\,
            I => \N__21413\
        );

    \I__4910\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21410\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__21410\,
            I => \N__21407\
        );

    \I__4908\ : Span4Mux_s1_v
    port map (
            O => \N__21407\,
            I => \N__21403\
        );

    \I__4907\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21400\
        );

    \I__4906\ : Sp12to4
    port map (
            O => \N__21403\,
            I => \N__21396\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__21400\,
            I => \N__21393\
        );

    \I__4904\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21390\
        );

    \I__4903\ : Span12Mux_h
    port map (
            O => \N__21396\,
            I => \N__21387\
        );

    \I__4902\ : Odrv12
    port map (
            O => \N__21393\,
            I => \M_this_internal_address_qZ0Z_5\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__21390\,
            I => \M_this_internal_address_qZ0Z_5\
        );

    \I__4900\ : Odrv12
    port map (
            O => \N__21387\,
            I => \M_this_internal_address_qZ0Z_5\
        );

    \I__4899\ : InMux
    port map (
            O => \N__21380\,
            I => \N__21377\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__21377\,
            I => \M_this_internal_address_q_3_ns_1_5\
        );

    \I__4897\ : CascadeMux
    port map (
            O => \N__21374\,
            I => \N__21371\
        );

    \I__4896\ : CascadeBuf
    port map (
            O => \N__21371\,
            I => \N__21368\
        );

    \I__4895\ : CascadeMux
    port map (
            O => \N__21368\,
            I => \N__21365\
        );

    \I__4894\ : CascadeBuf
    port map (
            O => \N__21365\,
            I => \N__21362\
        );

    \I__4893\ : CascadeMux
    port map (
            O => \N__21362\,
            I => \N__21359\
        );

    \I__4892\ : CascadeBuf
    port map (
            O => \N__21359\,
            I => \N__21356\
        );

    \I__4891\ : CascadeMux
    port map (
            O => \N__21356\,
            I => \N__21353\
        );

    \I__4890\ : CascadeBuf
    port map (
            O => \N__21353\,
            I => \N__21350\
        );

    \I__4889\ : CascadeMux
    port map (
            O => \N__21350\,
            I => \N__21347\
        );

    \I__4888\ : CascadeBuf
    port map (
            O => \N__21347\,
            I => \N__21344\
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__21344\,
            I => \N__21341\
        );

    \I__4886\ : CascadeBuf
    port map (
            O => \N__21341\,
            I => \N__21338\
        );

    \I__4885\ : CascadeMux
    port map (
            O => \N__21338\,
            I => \N__21335\
        );

    \I__4884\ : CascadeBuf
    port map (
            O => \N__21335\,
            I => \N__21332\
        );

    \I__4883\ : CascadeMux
    port map (
            O => \N__21332\,
            I => \N__21329\
        );

    \I__4882\ : CascadeBuf
    port map (
            O => \N__21329\,
            I => \N__21326\
        );

    \I__4881\ : CascadeMux
    port map (
            O => \N__21326\,
            I => \N__21323\
        );

    \I__4880\ : CascadeBuf
    port map (
            O => \N__21323\,
            I => \N__21320\
        );

    \I__4879\ : CascadeMux
    port map (
            O => \N__21320\,
            I => \N__21317\
        );

    \I__4878\ : CascadeBuf
    port map (
            O => \N__21317\,
            I => \N__21314\
        );

    \I__4877\ : CascadeMux
    port map (
            O => \N__21314\,
            I => \N__21311\
        );

    \I__4876\ : CascadeBuf
    port map (
            O => \N__21311\,
            I => \N__21308\
        );

    \I__4875\ : CascadeMux
    port map (
            O => \N__21308\,
            I => \N__21305\
        );

    \I__4874\ : CascadeBuf
    port map (
            O => \N__21305\,
            I => \N__21302\
        );

    \I__4873\ : CascadeMux
    port map (
            O => \N__21302\,
            I => \N__21299\
        );

    \I__4872\ : CascadeBuf
    port map (
            O => \N__21299\,
            I => \N__21296\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__21296\,
            I => \N__21293\
        );

    \I__4870\ : CascadeBuf
    port map (
            O => \N__21293\,
            I => \N__21290\
        );

    \I__4869\ : CascadeMux
    port map (
            O => \N__21290\,
            I => \N__21287\
        );

    \I__4868\ : CascadeBuf
    port map (
            O => \N__21287\,
            I => \N__21284\
        );

    \I__4867\ : CascadeMux
    port map (
            O => \N__21284\,
            I => \N__21281\
        );

    \I__4866\ : InMux
    port map (
            O => \N__21281\,
            I => \N__21276\
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__21280\,
            I => \N__21273\
        );

    \I__4864\ : InMux
    port map (
            O => \N__21279\,
            I => \N__21270\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__21276\,
            I => \N__21267\
        );

    \I__4862\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21264\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__21270\,
            I => \N__21261\
        );

    \I__4860\ : Span12Mux_h
    port map (
            O => \N__21267\,
            I => \N__21258\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__21264\,
            I => \M_this_internal_address_qZ0Z_6\
        );

    \I__4858\ : Odrv4
    port map (
            O => \N__21261\,
            I => \M_this_internal_address_qZ0Z_6\
        );

    \I__4857\ : Odrv12
    port map (
            O => \N__21258\,
            I => \M_this_internal_address_qZ0Z_6\
        );

    \I__4856\ : CascadeMux
    port map (
            O => \N__21251\,
            I => \N__21248\
        );

    \I__4855\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21245\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__21245\,
            I => \M_this_internal_address_q_3_ns_1_6\
        );

    \I__4853\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21239\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__21239\,
            I => \N__21236\
        );

    \I__4851\ : Odrv12
    port map (
            O => \N__21236\,
            I => \M_this_internal_address_q_3_ns_1_13\
        );

    \I__4850\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21226\
        );

    \I__4849\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21226\
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__21231\,
            I => \N__21220\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__21226\,
            I => \N__21216\
        );

    \I__4846\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21207\
        );

    \I__4845\ : InMux
    port map (
            O => \N__21224\,
            I => \N__21207\
        );

    \I__4844\ : InMux
    port map (
            O => \N__21223\,
            I => \N__21204\
        );

    \I__4843\ : InMux
    port map (
            O => \N__21220\,
            I => \N__21199\
        );

    \I__4842\ : InMux
    port map (
            O => \N__21219\,
            I => \N__21199\
        );

    \I__4841\ : Span4Mux_v
    port map (
            O => \N__21216\,
            I => \N__21193\
        );

    \I__4840\ : InMux
    port map (
            O => \N__21215\,
            I => \N__21190\
        );

    \I__4839\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21183\
        );

    \I__4838\ : InMux
    port map (
            O => \N__21213\,
            I => \N__21183\
        );

    \I__4837\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21183\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__21207\,
            I => \N__21178\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__21204\,
            I => \N__21178\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__21199\,
            I => \N__21175\
        );

    \I__4833\ : InMux
    port map (
            O => \N__21198\,
            I => \N__21172\
        );

    \I__4832\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21166\
        );

    \I__4831\ : InMux
    port map (
            O => \N__21196\,
            I => \N__21163\
        );

    \I__4830\ : Span4Mux_h
    port map (
            O => \N__21193\,
            I => \N__21160\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__21190\,
            I => \N__21155\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__21183\,
            I => \N__21155\
        );

    \I__4827\ : Span4Mux_h
    port map (
            O => \N__21178\,
            I => \N__21152\
        );

    \I__4826\ : Span4Mux_v
    port map (
            O => \N__21175\,
            I => \N__21147\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__21172\,
            I => \N__21147\
        );

    \I__4824\ : InMux
    port map (
            O => \N__21171\,
            I => \N__21142\
        );

    \I__4823\ : InMux
    port map (
            O => \N__21170\,
            I => \N__21142\
        );

    \I__4822\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21139\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__21166\,
            I => \N_355\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__21163\,
            I => \N_355\
        );

    \I__4819\ : Odrv4
    port map (
            O => \N__21160\,
            I => \N_355\
        );

    \I__4818\ : Odrv12
    port map (
            O => \N__21155\,
            I => \N_355\
        );

    \I__4817\ : Odrv4
    port map (
            O => \N__21152\,
            I => \N_355\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__21147\,
            I => \N_355\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__21142\,
            I => \N_355\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__21139\,
            I => \N_355\
        );

    \I__4813\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21119\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__21119\,
            I => \M_this_internal_address_q_3_ns_1_12\
        );

    \I__4811\ : InMux
    port map (
            O => \N__21116\,
            I => \N__21110\
        );

    \I__4810\ : InMux
    port map (
            O => \N__21115\,
            I => \N__21107\
        );

    \I__4809\ : InMux
    port map (
            O => \N__21114\,
            I => \N__21104\
        );

    \I__4808\ : InMux
    port map (
            O => \N__21113\,
            I => \N__21101\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__21110\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__21107\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__21104\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__21101\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__21092\,
            I => \N__21088\
        );

    \I__4802\ : CascadeMux
    port map (
            O => \N__21091\,
            I => \N__21085\
        );

    \I__4801\ : InMux
    port map (
            O => \N__21088\,
            I => \N__21082\
        );

    \I__4800\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21079\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__21082\,
            I => \N__21073\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__21079\,
            I => \N__21073\
        );

    \I__4797\ : InMux
    port map (
            O => \N__21078\,
            I => \N__21070\
        );

    \I__4796\ : Span4Mux_v
    port map (
            O => \N__21073\,
            I => \N__21067\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__21070\,
            I => \N__21064\
        );

    \I__4794\ : Sp12to4
    port map (
            O => \N__21067\,
            I => \N__21061\
        );

    \I__4793\ : Span4Mux_v
    port map (
            O => \N__21064\,
            I => \N__21058\
        );

    \I__4792\ : Span12Mux_h
    port map (
            O => \N__21061\,
            I => \N__21055\
        );

    \I__4791\ : Sp12to4
    port map (
            O => \N__21058\,
            I => \N__21052\
        );

    \I__4790\ : Odrv12
    port map (
            O => \N__21055\,
            I => port_data_c_5
        );

    \I__4789\ : Odrv12
    port map (
            O => \N__21052\,
            I => port_data_c_5
        );

    \I__4788\ : CascadeMux
    port map (
            O => \N__21047\,
            I => \N__21044\
        );

    \I__4787\ : InMux
    port map (
            O => \N__21044\,
            I => \N__21039\
        );

    \I__4786\ : CascadeMux
    port map (
            O => \N__21043\,
            I => \N__21036\
        );

    \I__4785\ : CascadeMux
    port map (
            O => \N__21042\,
            I => \N__21032\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__21039\,
            I => \N__21029\
        );

    \I__4783\ : InMux
    port map (
            O => \N__21036\,
            I => \N__21026\
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__21035\,
            I => \N__21023\
        );

    \I__4781\ : InMux
    port map (
            O => \N__21032\,
            I => \N__21020\
        );

    \I__4780\ : Span4Mux_v
    port map (
            O => \N__21029\,
            I => \N__21017\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__21026\,
            I => \N__21014\
        );

    \I__4778\ : InMux
    port map (
            O => \N__21023\,
            I => \N__21011\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__21020\,
            I => \N__21008\
        );

    \I__4776\ : Span4Mux_h
    port map (
            O => \N__21017\,
            I => \N__21001\
        );

    \I__4775\ : Span4Mux_v
    port map (
            O => \N__21014\,
            I => \N__21001\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__21011\,
            I => \N__21001\
        );

    \I__4773\ : Span4Mux_v
    port map (
            O => \N__21008\,
            I => \N__20998\
        );

    \I__4772\ : Span4Mux_h
    port map (
            O => \N__21001\,
            I => \N__20995\
        );

    \I__4771\ : Sp12to4
    port map (
            O => \N__20998\,
            I => \N__20992\
        );

    \I__4770\ : Span4Mux_v
    port map (
            O => \N__20995\,
            I => \N__20989\
        );

    \I__4769\ : Span12Mux_h
    port map (
            O => \N__20992\,
            I => \N__20986\
        );

    \I__4768\ : Span4Mux_v
    port map (
            O => \N__20989\,
            I => \N__20983\
        );

    \I__4767\ : Span12Mux_v
    port map (
            O => \N__20986\,
            I => \N__20980\
        );

    \I__4766\ : Span4Mux_v
    port map (
            O => \N__20983\,
            I => \N__20977\
        );

    \I__4765\ : Odrv12
    port map (
            O => \N__20980\,
            I => port_data_c_1
        );

    \I__4764\ : Odrv4
    port map (
            O => \N__20977\,
            I => port_data_c_1
        );

    \I__4763\ : InMux
    port map (
            O => \N__20972\,
            I => \N__20969\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__20969\,
            I => \N__20963\
        );

    \I__4761\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20960\
        );

    \I__4760\ : InMux
    port map (
            O => \N__20967\,
            I => \N__20957\
        );

    \I__4759\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20953\
        );

    \I__4758\ : Span4Mux_h
    port map (
            O => \N__20963\,
            I => \N__20949\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__20960\,
            I => \N__20946\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__20957\,
            I => \N__20943\
        );

    \I__4755\ : InMux
    port map (
            O => \N__20956\,
            I => \N__20940\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__20953\,
            I => \N__20935\
        );

    \I__4753\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20932\
        );

    \I__4752\ : Span4Mux_v
    port map (
            O => \N__20949\,
            I => \N__20927\
        );

    \I__4751\ : Span4Mux_h
    port map (
            O => \N__20946\,
            I => \N__20927\
        );

    \I__4750\ : Span4Mux_v
    port map (
            O => \N__20943\,
            I => \N__20922\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__20940\,
            I => \N__20922\
        );

    \I__4748\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20919\
        );

    \I__4747\ : InMux
    port map (
            O => \N__20938\,
            I => \N__20916\
        );

    \I__4746\ : Span12Mux_s11_h
    port map (
            O => \N__20935\,
            I => \N__20913\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__20932\,
            I => \N__20910\
        );

    \I__4744\ : Span4Mux_v
    port map (
            O => \N__20927\,
            I => \N__20907\
        );

    \I__4743\ : Span4Mux_v
    port map (
            O => \N__20922\,
            I => \N__20902\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__20919\,
            I => \N__20902\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__20916\,
            I => \N__20899\
        );

    \I__4740\ : Span12Mux_v
    port map (
            O => \N__20913\,
            I => \N__20894\
        );

    \I__4739\ : Span12Mux_s11_h
    port map (
            O => \N__20910\,
            I => \N__20894\
        );

    \I__4738\ : Span4Mux_v
    port map (
            O => \N__20907\,
            I => \N__20887\
        );

    \I__4737\ : Span4Mux_h
    port map (
            O => \N__20902\,
            I => \N__20887\
        );

    \I__4736\ : Span4Mux_h
    port map (
            O => \N__20899\,
            I => \N__20887\
        );

    \I__4735\ : Odrv12
    port map (
            O => \N__20894\,
            I => \M_this_sprites_ram_write_data_1\
        );

    \I__4734\ : Odrv4
    port map (
            O => \N__20887\,
            I => \M_this_sprites_ram_write_data_1\
        );

    \I__4733\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20878\
        );

    \I__4732\ : InMux
    port map (
            O => \N__20881\,
            I => \N__20875\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__20878\,
            I => \N__20870\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__20875\,
            I => \N__20867\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__20874\,
            I => \N__20864\
        );

    \I__4728\ : CascadeMux
    port map (
            O => \N__20873\,
            I => \N__20861\
        );

    \I__4727\ : Span12Mux_h
    port map (
            O => \N__20870\,
            I => \N__20858\
        );

    \I__4726\ : Span4Mux_v
    port map (
            O => \N__20867\,
            I => \N__20855\
        );

    \I__4725\ : InMux
    port map (
            O => \N__20864\,
            I => \N__20850\
        );

    \I__4724\ : InMux
    port map (
            O => \N__20861\,
            I => \N__20850\
        );

    \I__4723\ : Span12Mux_v
    port map (
            O => \N__20858\,
            I => \N__20847\
        );

    \I__4722\ : Sp12to4
    port map (
            O => \N__20855\,
            I => \N__20842\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__20850\,
            I => \N__20842\
        );

    \I__4720\ : Span12Mux_h
    port map (
            O => \N__20847\,
            I => \N__20839\
        );

    \I__4719\ : Span12Mux_h
    port map (
            O => \N__20842\,
            I => \N__20836\
        );

    \I__4718\ : Odrv12
    port map (
            O => \N__20839\,
            I => port_data_c_0
        );

    \I__4717\ : Odrv12
    port map (
            O => \N__20836\,
            I => port_data_c_0
        );

    \I__4716\ : CascadeMux
    port map (
            O => \N__20831\,
            I => \N__20828\
        );

    \I__4715\ : InMux
    port map (
            O => \N__20828\,
            I => \N__20824\
        );

    \I__4714\ : CascadeMux
    port map (
            O => \N__20827\,
            I => \N__20820\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__20824\,
            I => \N__20817\
        );

    \I__4712\ : InMux
    port map (
            O => \N__20823\,
            I => \N__20812\
        );

    \I__4711\ : InMux
    port map (
            O => \N__20820\,
            I => \N__20812\
        );

    \I__4710\ : Span4Mux_v
    port map (
            O => \N__20817\,
            I => \N__20809\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__20812\,
            I => \N__20806\
        );

    \I__4708\ : Span4Mux_v
    port map (
            O => \N__20809\,
            I => \N__20803\
        );

    \I__4707\ : Span12Mux_v
    port map (
            O => \N__20806\,
            I => \N__20800\
        );

    \I__4706\ : Sp12to4
    port map (
            O => \N__20803\,
            I => \N__20797\
        );

    \I__4705\ : Span12Mux_h
    port map (
            O => \N__20800\,
            I => \N__20794\
        );

    \I__4704\ : Odrv12
    port map (
            O => \N__20797\,
            I => port_data_c_4
        );

    \I__4703\ : Odrv12
    port map (
            O => \N__20794\,
            I => port_data_c_4
        );

    \I__4702\ : InMux
    port map (
            O => \N__20789\,
            I => \N__20786\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__20786\,
            I => \N__20782\
        );

    \I__4700\ : InMux
    port map (
            O => \N__20785\,
            I => \N__20779\
        );

    \I__4699\ : Span4Mux_h
    port map (
            O => \N__20782\,
            I => \N__20774\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__20779\,
            I => \N__20771\
        );

    \I__4697\ : InMux
    port map (
            O => \N__20778\,
            I => \N__20768\
        );

    \I__4696\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20764\
        );

    \I__4695\ : Span4Mux_v
    port map (
            O => \N__20774\,
            I => \N__20758\
        );

    \I__4694\ : Span4Mux_h
    port map (
            O => \N__20771\,
            I => \N__20758\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__20768\,
            I => \N__20755\
        );

    \I__4692\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20752\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__20764\,
            I => \N__20749\
        );

    \I__4690\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20746\
        );

    \I__4689\ : Span4Mux_v
    port map (
            O => \N__20758\,
            I => \N__20739\
        );

    \I__4688\ : Span4Mux_h
    port map (
            O => \N__20755\,
            I => \N__20739\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__20752\,
            I => \N__20736\
        );

    \I__4686\ : Span4Mux_v
    port map (
            O => \N__20749\,
            I => \N__20731\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__20746\,
            I => \N__20731\
        );

    \I__4684\ : InMux
    port map (
            O => \N__20745\,
            I => \N__20728\
        );

    \I__4683\ : InMux
    port map (
            O => \N__20744\,
            I => \N__20725\
        );

    \I__4682\ : Span4Mux_v
    port map (
            O => \N__20739\,
            I => \N__20720\
        );

    \I__4681\ : Span4Mux_h
    port map (
            O => \N__20736\,
            I => \N__20720\
        );

    \I__4680\ : Span4Mux_h
    port map (
            O => \N__20731\,
            I => \N__20717\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__20728\,
            I => \N__20714\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__20725\,
            I => \N__20711\
        );

    \I__4677\ : Span4Mux_v
    port map (
            O => \N__20720\,
            I => \N__20702\
        );

    \I__4676\ : Span4Mux_v
    port map (
            O => \N__20717\,
            I => \N__20702\
        );

    \I__4675\ : Span4Mux_h
    port map (
            O => \N__20714\,
            I => \N__20702\
        );

    \I__4674\ : Span4Mux_h
    port map (
            O => \N__20711\,
            I => \N__20702\
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__20702\,
            I => \M_this_sprites_ram_write_data_0\
        );

    \I__4672\ : InMux
    port map (
            O => \N__20699\,
            I => \N__20696\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__20696\,
            I => \N__20693\
        );

    \I__4670\ : Span4Mux_v
    port map (
            O => \N__20693\,
            I => \N__20690\
        );

    \I__4669\ : Sp12to4
    port map (
            O => \N__20690\,
            I => \N__20687\
        );

    \I__4668\ : Span12Mux_h
    port map (
            O => \N__20687\,
            I => \N__20684\
        );

    \I__4667\ : Span12Mux_v
    port map (
            O => \N__20684\,
            I => \N__20681\
        );

    \I__4666\ : Odrv12
    port map (
            O => \N__20681\,
            I => port_address_in_7
        );

    \I__4665\ : InMux
    port map (
            O => \N__20678\,
            I => \N__20675\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__20675\,
            I => \N__20672\
        );

    \I__4663\ : Sp12to4
    port map (
            O => \N__20672\,
            I => \N__20669\
        );

    \I__4662\ : Span12Mux_v
    port map (
            O => \N__20669\,
            I => \N__20666\
        );

    \I__4661\ : Span12Mux_h
    port map (
            O => \N__20666\,
            I => \N__20663\
        );

    \I__4660\ : Odrv12
    port map (
            O => \N__20663\,
            I => port_address_in_6
        );

    \I__4659\ : CascadeMux
    port map (
            O => \N__20660\,
            I => \N__20657\
        );

    \I__4658\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20654\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__20654\,
            I => \N__20651\
        );

    \I__4656\ : Span4Mux_v
    port map (
            O => \N__20651\,
            I => \N__20648\
        );

    \I__4655\ : Span4Mux_v
    port map (
            O => \N__20648\,
            I => \N__20645\
        );

    \I__4654\ : Sp12to4
    port map (
            O => \N__20645\,
            I => \N__20642\
        );

    \I__4653\ : Span12Mux_h
    port map (
            O => \N__20642\,
            I => \N__20638\
        );

    \I__4652\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20635\
        );

    \I__4651\ : Odrv12
    port map (
            O => \N__20638\,
            I => port_rw_in
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__20635\,
            I => port_rw_in
        );

    \I__4649\ : CascadeMux
    port map (
            O => \N__20630\,
            I => \N__20627\
        );

    \I__4648\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20622\
        );

    \I__4647\ : InMux
    port map (
            O => \N__20626\,
            I => \N__20619\
        );

    \I__4646\ : InMux
    port map (
            O => \N__20625\,
            I => \N__20616\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__20622\,
            I => \N__20611\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__20619\,
            I => \N__20611\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__20616\,
            I => \N__20608\
        );

    \I__4642\ : Span4Mux_h
    port map (
            O => \N__20611\,
            I => \N__20603\
        );

    \I__4641\ : Span4Mux_h
    port map (
            O => \N__20608\,
            I => \N__20603\
        );

    \I__4640\ : Odrv4
    port map (
            O => \N__20603\,
            I => \this_vga_signals.N_185_0\
        );

    \I__4639\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20597\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__20597\,
            I => \N__20594\
        );

    \I__4637\ : Odrv4
    port map (
            O => \N__20594\,
            I => \this_vga_signals.M_this_state_q_srsts_0_i_o4_4Z0Z_4\
        );

    \I__4636\ : CascadeMux
    port map (
            O => \N__20591\,
            I => \N__20586\
        );

    \I__4635\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20583\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__20589\,
            I => \N__20580\
        );

    \I__4633\ : InMux
    port map (
            O => \N__20586\,
            I => \N__20577\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__20583\,
            I => \N__20574\
        );

    \I__4631\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20571\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__20577\,
            I => \N__20568\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__20574\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__20571\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__4627\ : Odrv4
    port map (
            O => \N__20568\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__4626\ : CascadeMux
    port map (
            O => \N__20561\,
            I => \this_vga_signals.M_this_state_q_srsts_0_i_o4_4Z0Z_4_cascade_\
        );

    \I__4625\ : CascadeMux
    port map (
            O => \N__20558\,
            I => \this_vga_signals.N_490_cascade_\
        );

    \I__4624\ : CascadeMux
    port map (
            O => \N__20555\,
            I => \this_vga_signals.N_386_cascade_\
        );

    \I__4623\ : CascadeMux
    port map (
            O => \N__20552\,
            I => \this_vga_signals.N_387_cascade_\
        );

    \I__4622\ : CascadeMux
    port map (
            O => \N__20549\,
            I => \N__20546\
        );

    \I__4621\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20540\
        );

    \I__4620\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20537\
        );

    \I__4619\ : InMux
    port map (
            O => \N__20544\,
            I => \N__20532\
        );

    \I__4618\ : InMux
    port map (
            O => \N__20543\,
            I => \N__20532\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__20540\,
            I => \N__20529\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__20537\,
            I => \N__20524\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__20532\,
            I => \N__20524\
        );

    \I__4614\ : Span4Mux_v
    port map (
            O => \N__20529\,
            I => \N__20521\
        );

    \I__4613\ : Span4Mux_v
    port map (
            O => \N__20524\,
            I => \N__20518\
        );

    \I__4612\ : Sp12to4
    port map (
            O => \N__20521\,
            I => \N__20513\
        );

    \I__4611\ : Sp12to4
    port map (
            O => \N__20518\,
            I => \N__20513\
        );

    \I__4610\ : Span12Mux_h
    port map (
            O => \N__20513\,
            I => \N__20510\
        );

    \I__4609\ : Odrv12
    port map (
            O => \N__20510\,
            I => port_address_in_1
        );

    \I__4608\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20502\
        );

    \I__4607\ : InMux
    port map (
            O => \N__20506\,
            I => \N__20499\
        );

    \I__4606\ : InMux
    port map (
            O => \N__20505\,
            I => \N__20496\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__20502\,
            I => \N__20491\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__20499\,
            I => \N__20491\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__20496\,
            I => \N__20488\
        );

    \I__4602\ : Span4Mux_v
    port map (
            O => \N__20491\,
            I => \N__20482\
        );

    \I__4601\ : Span4Mux_v
    port map (
            O => \N__20488\,
            I => \N__20482\
        );

    \I__4600\ : InMux
    port map (
            O => \N__20487\,
            I => \N__20479\
        );

    \I__4599\ : Sp12to4
    port map (
            O => \N__20482\,
            I => \N__20476\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__20479\,
            I => \N__20473\
        );

    \I__4597\ : Span12Mux_h
    port map (
            O => \N__20476\,
            I => \N__20470\
        );

    \I__4596\ : Span12Mux_v
    port map (
            O => \N__20473\,
            I => \N__20467\
        );

    \I__4595\ : Odrv12
    port map (
            O => \N__20470\,
            I => port_address_in_0
        );

    \I__4594\ : Odrv12
    port map (
            O => \N__20467\,
            I => port_address_in_0
        );

    \I__4593\ : CascadeMux
    port map (
            O => \N__20462\,
            I => \this_vga_signals.N_391_cascade_\
        );

    \I__4592\ : InMux
    port map (
            O => \N__20459\,
            I => \N__20453\
        );

    \I__4591\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20453\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__20453\,
            I => \this_vga_signals.N_490\
        );

    \I__4589\ : InMux
    port map (
            O => \N__20450\,
            I => \N__20442\
        );

    \I__4588\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20439\
        );

    \I__4587\ : InMux
    port map (
            O => \N__20448\,
            I => \N__20436\
        );

    \I__4586\ : InMux
    port map (
            O => \N__20447\,
            I => \N__20433\
        );

    \I__4585\ : InMux
    port map (
            O => \N__20446\,
            I => \N__20428\
        );

    \I__4584\ : InMux
    port map (
            O => \N__20445\,
            I => \N__20428\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__20442\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__20439\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__20436\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__20433\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__20428\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__4578\ : InMux
    port map (
            O => \N__20417\,
            I => \N__20414\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__20411\,
            I => \M_this_internal_address_q_RNO_1Z0Z_5\
        );

    \I__4575\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20405\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__20405\,
            I => \N__20402\
        );

    \I__4573\ : Odrv4
    port map (
            O => \N__20402\,
            I => \M_this_internal_address_q_RNO_1Z0Z_6\
        );

    \I__4572\ : InMux
    port map (
            O => \N__20399\,
            I => \N__20396\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__20393\,
            I => \M_this_internal_address_q_RNO_1Z0Z_12\
        );

    \I__4569\ : InMux
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__20387\,
            I => \M_this_internal_address_q_3_ns_1_11\
        );

    \I__4567\ : InMux
    port map (
            O => \N__20384\,
            I => \N__20381\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__20381\,
            I => \M_this_internal_address_q_3_ns_1_4\
        );

    \I__4565\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20375\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__20375\,
            I => \N__20372\
        );

    \I__4563\ : Span4Mux_h
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__4562\ : Odrv4
    port map (
            O => \N__20369\,
            I => \M_this_internal_address_q_RNO_1Z0Z_4\
        );

    \I__4561\ : CascadeMux
    port map (
            O => \N__20366\,
            I => \N__20363\
        );

    \I__4560\ : CascadeBuf
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__4559\ : CascadeMux
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__4558\ : CascadeBuf
    port map (
            O => \N__20357\,
            I => \N__20354\
        );

    \I__4557\ : CascadeMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__4556\ : CascadeBuf
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__4555\ : CascadeMux
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__4554\ : CascadeBuf
    port map (
            O => \N__20345\,
            I => \N__20342\
        );

    \I__4553\ : CascadeMux
    port map (
            O => \N__20342\,
            I => \N__20339\
        );

    \I__4552\ : CascadeBuf
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__4551\ : CascadeMux
    port map (
            O => \N__20336\,
            I => \N__20333\
        );

    \I__4550\ : CascadeBuf
    port map (
            O => \N__20333\,
            I => \N__20330\
        );

    \I__4549\ : CascadeMux
    port map (
            O => \N__20330\,
            I => \N__20327\
        );

    \I__4548\ : CascadeBuf
    port map (
            O => \N__20327\,
            I => \N__20324\
        );

    \I__4547\ : CascadeMux
    port map (
            O => \N__20324\,
            I => \N__20321\
        );

    \I__4546\ : CascadeBuf
    port map (
            O => \N__20321\,
            I => \N__20318\
        );

    \I__4545\ : CascadeMux
    port map (
            O => \N__20318\,
            I => \N__20315\
        );

    \I__4544\ : CascadeBuf
    port map (
            O => \N__20315\,
            I => \N__20312\
        );

    \I__4543\ : CascadeMux
    port map (
            O => \N__20312\,
            I => \N__20309\
        );

    \I__4542\ : CascadeBuf
    port map (
            O => \N__20309\,
            I => \N__20306\
        );

    \I__4541\ : CascadeMux
    port map (
            O => \N__20306\,
            I => \N__20303\
        );

    \I__4540\ : CascadeBuf
    port map (
            O => \N__20303\,
            I => \N__20300\
        );

    \I__4539\ : CascadeMux
    port map (
            O => \N__20300\,
            I => \N__20297\
        );

    \I__4538\ : CascadeBuf
    port map (
            O => \N__20297\,
            I => \N__20294\
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__20294\,
            I => \N__20291\
        );

    \I__4536\ : CascadeBuf
    port map (
            O => \N__20291\,
            I => \N__20288\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__20288\,
            I => \N__20285\
        );

    \I__4534\ : CascadeBuf
    port map (
            O => \N__20285\,
            I => \N__20282\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__20282\,
            I => \N__20279\
        );

    \I__4532\ : CascadeBuf
    port map (
            O => \N__20279\,
            I => \N__20276\
        );

    \I__4531\ : CascadeMux
    port map (
            O => \N__20276\,
            I => \N__20273\
        );

    \I__4530\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20270\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__20270\,
            I => \N__20266\
        );

    \I__4528\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20263\
        );

    \I__4527\ : Span4Mux_v
    port map (
            O => \N__20266\,
            I => \N__20260\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__20263\,
            I => \N__20256\
        );

    \I__4525\ : Span4Mux_h
    port map (
            O => \N__20260\,
            I => \N__20253\
        );

    \I__4524\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20250\
        );

    \I__4523\ : Span4Mux_v
    port map (
            O => \N__20256\,
            I => \N__20245\
        );

    \I__4522\ : Span4Mux_v
    port map (
            O => \N__20253\,
            I => \N__20245\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__20250\,
            I => \M_this_internal_address_qZ0Z_4\
        );

    \I__4520\ : Odrv4
    port map (
            O => \N__20245\,
            I => \M_this_internal_address_qZ0Z_4\
        );

    \I__4519\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20237\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__20237\,
            I => \N__20234\
        );

    \I__4517\ : Span4Mux_h
    port map (
            O => \N__20234\,
            I => \N__20231\
        );

    \I__4516\ : Span4Mux_h
    port map (
            O => \N__20231\,
            I => \N__20228\
        );

    \I__4515\ : Span4Mux_h
    port map (
            O => \N__20228\,
            I => \N__20225\
        );

    \I__4514\ : Odrv4
    port map (
            O => \N__20225\,
            I => \M_this_vram_write_data_1\
        );

    \I__4513\ : IoInMux
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__20219\,
            I => \N__20215\
        );

    \I__4511\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20211\
        );

    \I__4510\ : Span4Mux_s3_h
    port map (
            O => \N__20215\,
            I => \N__20208\
        );

    \I__4509\ : InMux
    port map (
            O => \N__20214\,
            I => \N__20205\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__20211\,
            I => \N__20202\
        );

    \I__4507\ : Span4Mux_v
    port map (
            O => \N__20208\,
            I => \N__20199\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__20205\,
            I => \N__20196\
        );

    \I__4505\ : Span4Mux_v
    port map (
            O => \N__20202\,
            I => \N__20193\
        );

    \I__4504\ : Sp12to4
    port map (
            O => \N__20199\,
            I => \N__20189\
        );

    \I__4503\ : Span4Mux_v
    port map (
            O => \N__20196\,
            I => \N__20186\
        );

    \I__4502\ : Span4Mux_v
    port map (
            O => \N__20193\,
            I => \N__20183\
        );

    \I__4501\ : InMux
    port map (
            O => \N__20192\,
            I => \N__20180\
        );

    \I__4500\ : Span12Mux_h
    port map (
            O => \N__20189\,
            I => \N__20177\
        );

    \I__4499\ : Sp12to4
    port map (
            O => \N__20186\,
            I => \N__20174\
        );

    \I__4498\ : Span4Mux_h
    port map (
            O => \N__20183\,
            I => \N__20171\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__20180\,
            I => \N__20168\
        );

    \I__4496\ : Span12Mux_v
    port map (
            O => \N__20177\,
            I => \N__20162\
        );

    \I__4495\ : Span12Mux_h
    port map (
            O => \N__20174\,
            I => \N__20162\
        );

    \I__4494\ : Span4Mux_h
    port map (
            O => \N__20171\,
            I => \N__20157\
        );

    \I__4493\ : Span4Mux_v
    port map (
            O => \N__20168\,
            I => \N__20157\
        );

    \I__4492\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20154\
        );

    \I__4491\ : Odrv12
    port map (
            O => \N__20162\,
            I => \N_235_0\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__20157\,
            I => \N_235_0\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__20154\,
            I => \N_235_0\
        );

    \I__4488\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20144\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__20144\,
            I => \this_vga_signals.N_319\
        );

    \I__4486\ : CascadeMux
    port map (
            O => \N__20141\,
            I => \N__20137\
        );

    \I__4485\ : InMux
    port map (
            O => \N__20140\,
            I => \N__20134\
        );

    \I__4484\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20131\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__20134\,
            I => un19_i_i_i_a2
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__20131\,
            I => un19_i_i_i_a2
        );

    \I__4481\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20123\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__20123\,
            I => \M_this_internal_address_q_RNO_1Z0Z_11\
        );

    \I__4479\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__20117\,
            I => \M_this_internal_address_q_3_ns_1_0\
        );

    \I__4477\ : InMux
    port map (
            O => \N__20114\,
            I => \N__20111\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__20111\,
            I => \N__20108\
        );

    \I__4475\ : Odrv4
    port map (
            O => \N__20108\,
            I => \M_this_internal_address_q_RNO_1Z0Z_0\
        );

    \I__4474\ : CascadeMux
    port map (
            O => \N__20105\,
            I => \N__20102\
        );

    \I__4473\ : CascadeBuf
    port map (
            O => \N__20102\,
            I => \N__20099\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__20099\,
            I => \N__20096\
        );

    \I__4471\ : CascadeBuf
    port map (
            O => \N__20096\,
            I => \N__20093\
        );

    \I__4470\ : CascadeMux
    port map (
            O => \N__20093\,
            I => \N__20090\
        );

    \I__4469\ : CascadeBuf
    port map (
            O => \N__20090\,
            I => \N__20087\
        );

    \I__4468\ : CascadeMux
    port map (
            O => \N__20087\,
            I => \N__20084\
        );

    \I__4467\ : CascadeBuf
    port map (
            O => \N__20084\,
            I => \N__20081\
        );

    \I__4466\ : CascadeMux
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__4465\ : CascadeBuf
    port map (
            O => \N__20078\,
            I => \N__20075\
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__20075\,
            I => \N__20072\
        );

    \I__4463\ : CascadeBuf
    port map (
            O => \N__20072\,
            I => \N__20069\
        );

    \I__4462\ : CascadeMux
    port map (
            O => \N__20069\,
            I => \N__20066\
        );

    \I__4461\ : CascadeBuf
    port map (
            O => \N__20066\,
            I => \N__20063\
        );

    \I__4460\ : CascadeMux
    port map (
            O => \N__20063\,
            I => \N__20060\
        );

    \I__4459\ : CascadeBuf
    port map (
            O => \N__20060\,
            I => \N__20057\
        );

    \I__4458\ : CascadeMux
    port map (
            O => \N__20057\,
            I => \N__20054\
        );

    \I__4457\ : CascadeBuf
    port map (
            O => \N__20054\,
            I => \N__20051\
        );

    \I__4456\ : CascadeMux
    port map (
            O => \N__20051\,
            I => \N__20048\
        );

    \I__4455\ : CascadeBuf
    port map (
            O => \N__20048\,
            I => \N__20045\
        );

    \I__4454\ : CascadeMux
    port map (
            O => \N__20045\,
            I => \N__20042\
        );

    \I__4453\ : CascadeBuf
    port map (
            O => \N__20042\,
            I => \N__20039\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__20039\,
            I => \N__20036\
        );

    \I__4451\ : CascadeBuf
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__4449\ : CascadeBuf
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__4448\ : CascadeMux
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__4447\ : CascadeBuf
    port map (
            O => \N__20024\,
            I => \N__20021\
        );

    \I__4446\ : CascadeMux
    port map (
            O => \N__20021\,
            I => \N__20018\
        );

    \I__4445\ : CascadeBuf
    port map (
            O => \N__20018\,
            I => \N__20015\
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__20015\,
            I => \N__20012\
        );

    \I__4443\ : InMux
    port map (
            O => \N__20012\,
            I => \N__20008\
        );

    \I__4442\ : InMux
    port map (
            O => \N__20011\,
            I => \N__20005\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__20008\,
            I => \N__20001\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__20005\,
            I => \N__19998\
        );

    \I__4439\ : InMux
    port map (
            O => \N__20004\,
            I => \N__19995\
        );

    \I__4438\ : Span12Mux_s9_v
    port map (
            O => \N__20001\,
            I => \N__19992\
        );

    \I__4437\ : Odrv4
    port map (
            O => \N__19998\,
            I => \M_this_internal_address_qZ0Z_0\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__19995\,
            I => \M_this_internal_address_qZ0Z_0\
        );

    \I__4435\ : Odrv12
    port map (
            O => \N__19992\,
            I => \M_this_internal_address_qZ0Z_0\
        );

    \I__4434\ : InMux
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__19982\,
            I => \N__19979\
        );

    \I__4432\ : Odrv4
    port map (
            O => \N__19979\,
            I => \M_this_internal_address_q_3_ns_1_1\
        );

    \I__4431\ : InMux
    port map (
            O => \N__19976\,
            I => \N__19973\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__19973\,
            I => \N__19970\
        );

    \I__4429\ : Span4Mux_h
    port map (
            O => \N__19970\,
            I => \N__19967\
        );

    \I__4428\ : Odrv4
    port map (
            O => \N__19967\,
            I => \M_this_internal_address_q_RNO_1Z0Z_1\
        );

    \I__4427\ : CascadeMux
    port map (
            O => \N__19964\,
            I => \N__19961\
        );

    \I__4426\ : CascadeBuf
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__4425\ : CascadeMux
    port map (
            O => \N__19958\,
            I => \N__19955\
        );

    \I__4424\ : CascadeBuf
    port map (
            O => \N__19955\,
            I => \N__19952\
        );

    \I__4423\ : CascadeMux
    port map (
            O => \N__19952\,
            I => \N__19949\
        );

    \I__4422\ : CascadeBuf
    port map (
            O => \N__19949\,
            I => \N__19946\
        );

    \I__4421\ : CascadeMux
    port map (
            O => \N__19946\,
            I => \N__19943\
        );

    \I__4420\ : CascadeBuf
    port map (
            O => \N__19943\,
            I => \N__19940\
        );

    \I__4419\ : CascadeMux
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__4418\ : CascadeBuf
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__4417\ : CascadeMux
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__4416\ : CascadeBuf
    port map (
            O => \N__19931\,
            I => \N__19928\
        );

    \I__4415\ : CascadeMux
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__4414\ : CascadeBuf
    port map (
            O => \N__19925\,
            I => \N__19922\
        );

    \I__4413\ : CascadeMux
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__4412\ : CascadeBuf
    port map (
            O => \N__19919\,
            I => \N__19916\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__19916\,
            I => \N__19913\
        );

    \I__4410\ : CascadeBuf
    port map (
            O => \N__19913\,
            I => \N__19910\
        );

    \I__4409\ : CascadeMux
    port map (
            O => \N__19910\,
            I => \N__19907\
        );

    \I__4408\ : CascadeBuf
    port map (
            O => \N__19907\,
            I => \N__19904\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__19904\,
            I => \N__19901\
        );

    \I__4406\ : CascadeBuf
    port map (
            O => \N__19901\,
            I => \N__19898\
        );

    \I__4405\ : CascadeMux
    port map (
            O => \N__19898\,
            I => \N__19895\
        );

    \I__4404\ : CascadeBuf
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__4403\ : CascadeMux
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__4402\ : CascadeBuf
    port map (
            O => \N__19889\,
            I => \N__19886\
        );

    \I__4401\ : CascadeMux
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__4400\ : CascadeBuf
    port map (
            O => \N__19883\,
            I => \N__19880\
        );

    \I__4399\ : CascadeMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__4398\ : CascadeBuf
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__4397\ : CascadeMux
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__4396\ : InMux
    port map (
            O => \N__19871\,
            I => \N__19868\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__19868\,
            I => \N__19865\
        );

    \I__4394\ : Span4Mux_s2_v
    port map (
            O => \N__19865\,
            I => \N__19862\
        );

    \I__4393\ : Span4Mux_h
    port map (
            O => \N__19862\,
            I => \N__19857\
        );

    \I__4392\ : InMux
    port map (
            O => \N__19861\,
            I => \N__19854\
        );

    \I__4391\ : InMux
    port map (
            O => \N__19860\,
            I => \N__19851\
        );

    \I__4390\ : Span4Mux_h
    port map (
            O => \N__19857\,
            I => \N__19848\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__19854\,
            I => \N__19843\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__19851\,
            I => \N__19843\
        );

    \I__4387\ : Span4Mux_v
    port map (
            O => \N__19848\,
            I => \N__19840\
        );

    \I__4386\ : Odrv4
    port map (
            O => \N__19843\,
            I => \M_this_internal_address_qZ0Z_1\
        );

    \I__4385\ : Odrv4
    port map (
            O => \N__19840\,
            I => \M_this_internal_address_qZ0Z_1\
        );

    \I__4384\ : InMux
    port map (
            O => \N__19835\,
            I => \N__19832\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__19832\,
            I => \N_476\
        );

    \I__4382\ : InMux
    port map (
            O => \N__19829\,
            I => \N__19825\
        );

    \I__4381\ : InMux
    port map (
            O => \N__19828\,
            I => \N__19822\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__19825\,
            I => \N__19816\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__19822\,
            I => \N__19816\
        );

    \I__4378\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19813\
        );

    \I__4377\ : Span4Mux_h
    port map (
            O => \N__19816\,
            I => \N__19808\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__19813\,
            I => \N__19808\
        );

    \I__4375\ : Span4Mux_v
    port map (
            O => \N__19808\,
            I => \N__19805\
        );

    \I__4374\ : Odrv4
    port map (
            O => \N__19805\,
            I => \N_240\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__19802\,
            I => \N__19795\
        );

    \I__4372\ : InMux
    port map (
            O => \N__19801\,
            I => \N__19789\
        );

    \I__4371\ : InMux
    port map (
            O => \N__19800\,
            I => \N__19789\
        );

    \I__4370\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19786\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19798\,
            I => \N__19783\
        );

    \I__4368\ : InMux
    port map (
            O => \N__19795\,
            I => \N__19778\
        );

    \I__4367\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19778\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__19789\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__19786\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__19783\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__19778\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__19769\,
            I => \this_vga_signals.N_343_cascade_\
        );

    \I__4361\ : InMux
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__19763\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_c3_0
        );

    \I__4359\ : InMux
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__19757\,
            I => \N__19751\
        );

    \I__4357\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19746\
        );

    \I__4356\ : InMux
    port map (
            O => \N__19755\,
            I => \N__19746\
        );

    \I__4355\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19743\
        );

    \I__4354\ : Odrv4
    port map (
            O => \N__19751\,
            I => \this_ppu_sprites_N_2_1\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__19746\,
            I => \this_ppu_sprites_N_2_1\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__19743\,
            I => \this_ppu_sprites_N_2_1\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__19736\,
            I => \N__19733\
        );

    \I__4350\ : CascadeBuf
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__4348\ : CascadeBuf
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__4347\ : CascadeMux
    port map (
            O => \N__19724\,
            I => \N__19721\
        );

    \I__4346\ : CascadeBuf
    port map (
            O => \N__19721\,
            I => \N__19718\
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__4344\ : CascadeBuf
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__4342\ : CascadeBuf
    port map (
            O => \N__19709\,
            I => \N__19706\
        );

    \I__4341\ : CascadeMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__4340\ : CascadeBuf
    port map (
            O => \N__19703\,
            I => \N__19700\
        );

    \I__4339\ : CascadeMux
    port map (
            O => \N__19700\,
            I => \N__19697\
        );

    \I__4338\ : CascadeBuf
    port map (
            O => \N__19697\,
            I => \N__19694\
        );

    \I__4337\ : CascadeMux
    port map (
            O => \N__19694\,
            I => \N__19691\
        );

    \I__4336\ : CascadeBuf
    port map (
            O => \N__19691\,
            I => \N__19688\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__19688\,
            I => \N__19685\
        );

    \I__4334\ : CascadeBuf
    port map (
            O => \N__19685\,
            I => \N__19682\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__19682\,
            I => \N__19679\
        );

    \I__4332\ : CascadeBuf
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__4331\ : CascadeMux
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__4330\ : CascadeBuf
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__4329\ : CascadeMux
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__4328\ : CascadeBuf
    port map (
            O => \N__19667\,
            I => \N__19664\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__4326\ : CascadeBuf
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__4324\ : CascadeBuf
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__4323\ : CascadeMux
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__4322\ : CascadeBuf
    port map (
            O => \N__19649\,
            I => \N__19646\
        );

    \I__4321\ : CascadeMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__4320\ : InMux
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__4318\ : Span12Mux_s10_h
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__4317\ : Span12Mux_v
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__4316\ : Odrv12
    port map (
            O => \N__19631\,
            I => \N_134_0\
        );

    \I__4315\ : InMux
    port map (
            O => \N__19628\,
            I => \N__19625\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__19625\,
            I => \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_4\
        );

    \I__4313\ : CascadeMux
    port map (
            O => \N__19622\,
            I => \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_4_cascade_\
        );

    \I__4312\ : InMux
    port map (
            O => \N__19619\,
            I => \N__19616\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__19616\,
            I => \this_vga_signals.M_this_state_q_srsts_0_i_1Z0Z_4\
        );

    \I__4310\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__19610\,
            I => \this_vga_signals.M_this_state_q_srsts_0_i_0Z0Z_4\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__19607\,
            I => \N__19604\
        );

    \I__4307\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19601\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__19601\,
            I => \this_vga_signals.N_224_0\
        );

    \I__4305\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__19595\,
            I => \N__19591\
        );

    \I__4303\ : IoInMux
    port map (
            O => \N__19594\,
            I => \N__19588\
        );

    \I__4302\ : Span4Mux_v
    port map (
            O => \N__19591\,
            I => \N__19585\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__19588\,
            I => \N__19582\
        );

    \I__4300\ : Span4Mux_v
    port map (
            O => \N__19585\,
            I => \N__19579\
        );

    \I__4299\ : Span12Mux_s11_v
    port map (
            O => \N__19582\,
            I => \N__19576\
        );

    \I__4298\ : Odrv4
    port map (
            O => \N__19579\,
            I => \M_this_state_q_nss_0\
        );

    \I__4297\ : Odrv12
    port map (
            O => \N__19576\,
            I => \M_this_state_q_nss_0\
        );

    \I__4296\ : CascadeMux
    port map (
            O => \N__19571\,
            I => \N__19568\
        );

    \I__4295\ : InMux
    port map (
            O => \N__19568\,
            I => \N__19564\
        );

    \I__4294\ : InMux
    port map (
            O => \N__19567\,
            I => \N__19561\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__19564\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__19561\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__4291\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19552\
        );

    \I__4290\ : InMux
    port map (
            O => \N__19555\,
            I => \N__19549\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__19552\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__19549\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__4287\ : CascadeMux
    port map (
            O => \N__19544\,
            I => \N__19541\
        );

    \I__4286\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19537\
        );

    \I__4285\ : InMux
    port map (
            O => \N__19540\,
            I => \N__19534\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__19537\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__19534\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__4282\ : CascadeMux
    port map (
            O => \N__19529\,
            I => \N__19526\
        );

    \I__4281\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19522\
        );

    \I__4280\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19519\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__19522\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__19519\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__4277\ : CascadeMux
    port map (
            O => \N__19514\,
            I => \N__19510\
        );

    \I__4276\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19507\
        );

    \I__4275\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19504\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__19507\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__19504\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__4272\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19495\
        );

    \I__4271\ : InMux
    port map (
            O => \N__19498\,
            I => \N__19492\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__19495\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__19492\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__4268\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19483\
        );

    \I__4267\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19480\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__19483\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__19480\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__19475\,
            I => \N__19472\
        );

    \I__4263\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19468\
        );

    \I__4262\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19465\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__19468\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__19465\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__19460\,
            I => \N__19456\
        );

    \I__4258\ : CascadeMux
    port map (
            O => \N__19459\,
            I => \N__19453\
        );

    \I__4257\ : InMux
    port map (
            O => \N__19456\,
            I => \N__19450\
        );

    \I__4256\ : InMux
    port map (
            O => \N__19453\,
            I => \N__19447\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__19450\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__19447\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__4253\ : InMux
    port map (
            O => \N__19442\,
            I => \N__19438\
        );

    \I__4252\ : InMux
    port map (
            O => \N__19441\,
            I => \N__19435\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__19438\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__19435\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__4249\ : CascadeMux
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__4248\ : InMux
    port map (
            O => \N__19427\,
            I => \N__19423\
        );

    \I__4247\ : InMux
    port map (
            O => \N__19426\,
            I => \N__19420\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__19423\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__19420\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__4244\ : InMux
    port map (
            O => \N__19415\,
            I => \N__19411\
        );

    \I__4243\ : InMux
    port map (
            O => \N__19414\,
            I => \N__19408\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__19411\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__19408\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__4240\ : CascadeMux
    port map (
            O => \N__19403\,
            I => \N__19399\
        );

    \I__4239\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19396\
        );

    \I__4238\ : InMux
    port map (
            O => \N__19399\,
            I => \N__19393\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__19396\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__19393\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__4235\ : CascadeMux
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__4234\ : InMux
    port map (
            O => \N__19385\,
            I => \N__19381\
        );

    \I__4233\ : InMux
    port map (
            O => \N__19384\,
            I => \N__19378\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__19381\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__19378\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__4230\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__19370\,
            I => \M_this_state_q_srsts_0_a2_1_9_4\
        );

    \I__4228\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__19364\,
            I => \M_this_state_q_srsts_0_a2_1_7_4\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__19361\,
            I => \M_this_state_q_srsts_0_a2_1_8_4_cascade_\
        );

    \I__4225\ : InMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__19355\,
            I => \M_this_state_q_srsts_0_a2_1_6_4\
        );

    \I__4223\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19346\
        );

    \I__4222\ : InMux
    port map (
            O => \N__19351\,
            I => \N__19346\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__19346\,
            I => \N__19341\
        );

    \I__4220\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19336\
        );

    \I__4219\ : InMux
    port map (
            O => \N__19344\,
            I => \N__19336\
        );

    \I__4218\ : Sp12to4
    port map (
            O => \N__19341\,
            I => \N__19331\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__19336\,
            I => \N__19331\
        );

    \I__4216\ : Span12Mux_v
    port map (
            O => \N__19331\,
            I => \N__19328\
        );

    \I__4215\ : Odrv12
    port map (
            O => \N__19328\,
            I => rst_n_c
        );

    \I__4214\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19322\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__19322\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__4212\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__19316\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__19313\,
            I => \N__19310\
        );

    \I__4209\ : CascadeBuf
    port map (
            O => \N__19310\,
            I => \N__19307\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__19307\,
            I => \N__19304\
        );

    \I__4207\ : CascadeBuf
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__4206\ : CascadeMux
    port map (
            O => \N__19301\,
            I => \N__19298\
        );

    \I__4205\ : CascadeBuf
    port map (
            O => \N__19298\,
            I => \N__19295\
        );

    \I__4204\ : CascadeMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__4203\ : CascadeBuf
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__19289\,
            I => \N__19286\
        );

    \I__4201\ : CascadeBuf
    port map (
            O => \N__19286\,
            I => \N__19283\
        );

    \I__4200\ : CascadeMux
    port map (
            O => \N__19283\,
            I => \N__19280\
        );

    \I__4199\ : CascadeBuf
    port map (
            O => \N__19280\,
            I => \N__19277\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__4197\ : CascadeBuf
    port map (
            O => \N__19274\,
            I => \N__19271\
        );

    \I__4196\ : CascadeMux
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__4195\ : CascadeBuf
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__19265\,
            I => \N__19262\
        );

    \I__4193\ : CascadeBuf
    port map (
            O => \N__19262\,
            I => \N__19259\
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__19259\,
            I => \N__19256\
        );

    \I__4191\ : CascadeBuf
    port map (
            O => \N__19256\,
            I => \N__19253\
        );

    \I__4190\ : CascadeMux
    port map (
            O => \N__19253\,
            I => \N__19250\
        );

    \I__4189\ : CascadeBuf
    port map (
            O => \N__19250\,
            I => \N__19247\
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__19247\,
            I => \N__19244\
        );

    \I__4187\ : CascadeBuf
    port map (
            O => \N__19244\,
            I => \N__19241\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__19241\,
            I => \N__19238\
        );

    \I__4185\ : CascadeBuf
    port map (
            O => \N__19238\,
            I => \N__19235\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__4183\ : CascadeBuf
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__19229\,
            I => \N__19226\
        );

    \I__4181\ : CascadeBuf
    port map (
            O => \N__19226\,
            I => \N__19223\
        );

    \I__4180\ : CascadeMux
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__4179\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19217\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__19217\,
            I => \N__19212\
        );

    \I__4177\ : InMux
    port map (
            O => \N__19216\,
            I => \N__19209\
        );

    \I__4176\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19206\
        );

    \I__4175\ : Span12Mux_s11_v
    port map (
            O => \N__19212\,
            I => \N__19203\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__19209\,
            I => \M_this_internal_address_qZ0Z_8\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__19206\,
            I => \M_this_internal_address_qZ0Z_8\
        );

    \I__4172\ : Odrv12
    port map (
            O => \N__19203\,
            I => \M_this_internal_address_qZ0Z_8\
        );

    \I__4171\ : InMux
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__19193\,
            I => \M_this_internal_address_q_RNO_1Z0Z_8\
        );

    \I__4169\ : InMux
    port map (
            O => \N__19190\,
            I => \bfn_16_22_0_\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__4167\ : CascadeBuf
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__4166\ : CascadeMux
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__4165\ : CascadeBuf
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__4164\ : CascadeMux
    port map (
            O => \N__19175\,
            I => \N__19172\
        );

    \I__4163\ : CascadeBuf
    port map (
            O => \N__19172\,
            I => \N__19169\
        );

    \I__4162\ : CascadeMux
    port map (
            O => \N__19169\,
            I => \N__19166\
        );

    \I__4161\ : CascadeBuf
    port map (
            O => \N__19166\,
            I => \N__19163\
        );

    \I__4160\ : CascadeMux
    port map (
            O => \N__19163\,
            I => \N__19160\
        );

    \I__4159\ : CascadeBuf
    port map (
            O => \N__19160\,
            I => \N__19157\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__19157\,
            I => \N__19154\
        );

    \I__4157\ : CascadeBuf
    port map (
            O => \N__19154\,
            I => \N__19151\
        );

    \I__4156\ : CascadeMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__4155\ : CascadeBuf
    port map (
            O => \N__19148\,
            I => \N__19145\
        );

    \I__4154\ : CascadeMux
    port map (
            O => \N__19145\,
            I => \N__19142\
        );

    \I__4153\ : CascadeBuf
    port map (
            O => \N__19142\,
            I => \N__19139\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__4151\ : CascadeBuf
    port map (
            O => \N__19136\,
            I => \N__19133\
        );

    \I__4150\ : CascadeMux
    port map (
            O => \N__19133\,
            I => \N__19130\
        );

    \I__4149\ : CascadeBuf
    port map (
            O => \N__19130\,
            I => \N__19127\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__19127\,
            I => \N__19124\
        );

    \I__4147\ : CascadeBuf
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__4146\ : CascadeMux
    port map (
            O => \N__19121\,
            I => \N__19118\
        );

    \I__4145\ : CascadeBuf
    port map (
            O => \N__19118\,
            I => \N__19115\
        );

    \I__4144\ : CascadeMux
    port map (
            O => \N__19115\,
            I => \N__19112\
        );

    \I__4143\ : CascadeBuf
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__4142\ : CascadeMux
    port map (
            O => \N__19109\,
            I => \N__19106\
        );

    \I__4141\ : CascadeBuf
    port map (
            O => \N__19106\,
            I => \N__19103\
        );

    \I__4140\ : CascadeMux
    port map (
            O => \N__19103\,
            I => \N__19100\
        );

    \I__4139\ : CascadeBuf
    port map (
            O => \N__19100\,
            I => \N__19097\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__19097\,
            I => \N__19094\
        );

    \I__4137\ : InMux
    port map (
            O => \N__19094\,
            I => \N__19090\
        );

    \I__4136\ : CascadeMux
    port map (
            O => \N__19093\,
            I => \N__19087\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__19090\,
            I => \N__19083\
        );

    \I__4134\ : InMux
    port map (
            O => \N__19087\,
            I => \N__19080\
        );

    \I__4133\ : InMux
    port map (
            O => \N__19086\,
            I => \N__19077\
        );

    \I__4132\ : Span12Mux_h
    port map (
            O => \N__19083\,
            I => \N__19074\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__19080\,
            I => \M_this_internal_address_qZ0Z_9\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__19077\,
            I => \M_this_internal_address_qZ0Z_9\
        );

    \I__4129\ : Odrv12
    port map (
            O => \N__19074\,
            I => \M_this_internal_address_qZ0Z_9\
        );

    \I__4128\ : InMux
    port map (
            O => \N__19067\,
            I => \N__19064\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__19064\,
            I => \M_this_internal_address_q_RNO_1Z0Z_9\
        );

    \I__4126\ : InMux
    port map (
            O => \N__19061\,
            I => \un1_M_this_internal_address_q_cry_8\
        );

    \I__4125\ : CascadeMux
    port map (
            O => \N__19058\,
            I => \N__19055\
        );

    \I__4124\ : CascadeBuf
    port map (
            O => \N__19055\,
            I => \N__19052\
        );

    \I__4123\ : CascadeMux
    port map (
            O => \N__19052\,
            I => \N__19049\
        );

    \I__4122\ : CascadeBuf
    port map (
            O => \N__19049\,
            I => \N__19046\
        );

    \I__4121\ : CascadeMux
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__4120\ : CascadeBuf
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__4118\ : CascadeBuf
    port map (
            O => \N__19037\,
            I => \N__19034\
        );

    \I__4117\ : CascadeMux
    port map (
            O => \N__19034\,
            I => \N__19031\
        );

    \I__4116\ : CascadeBuf
    port map (
            O => \N__19031\,
            I => \N__19028\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__19028\,
            I => \N__19025\
        );

    \I__4114\ : CascadeBuf
    port map (
            O => \N__19025\,
            I => \N__19022\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__4112\ : CascadeBuf
    port map (
            O => \N__19019\,
            I => \N__19016\
        );

    \I__4111\ : CascadeMux
    port map (
            O => \N__19016\,
            I => \N__19013\
        );

    \I__4110\ : CascadeBuf
    port map (
            O => \N__19013\,
            I => \N__19010\
        );

    \I__4109\ : CascadeMux
    port map (
            O => \N__19010\,
            I => \N__19007\
        );

    \I__4108\ : CascadeBuf
    port map (
            O => \N__19007\,
            I => \N__19004\
        );

    \I__4107\ : CascadeMux
    port map (
            O => \N__19004\,
            I => \N__19001\
        );

    \I__4106\ : CascadeBuf
    port map (
            O => \N__19001\,
            I => \N__18998\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__18998\,
            I => \N__18995\
        );

    \I__4104\ : CascadeBuf
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__18992\,
            I => \N__18989\
        );

    \I__4102\ : CascadeBuf
    port map (
            O => \N__18989\,
            I => \N__18986\
        );

    \I__4101\ : CascadeMux
    port map (
            O => \N__18986\,
            I => \N__18983\
        );

    \I__4100\ : CascadeBuf
    port map (
            O => \N__18983\,
            I => \N__18980\
        );

    \I__4099\ : CascadeMux
    port map (
            O => \N__18980\,
            I => \N__18977\
        );

    \I__4098\ : CascadeBuf
    port map (
            O => \N__18977\,
            I => \N__18974\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__18974\,
            I => \N__18971\
        );

    \I__4096\ : CascadeBuf
    port map (
            O => \N__18971\,
            I => \N__18968\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__18968\,
            I => \N__18965\
        );

    \I__4094\ : InMux
    port map (
            O => \N__18965\,
            I => \N__18962\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__18962\,
            I => \N__18959\
        );

    \I__4092\ : Span4Mux_s3_v
    port map (
            O => \N__18959\,
            I => \N__18955\
        );

    \I__4091\ : InMux
    port map (
            O => \N__18958\,
            I => \N__18952\
        );

    \I__4090\ : Sp12to4
    port map (
            O => \N__18955\,
            I => \N__18948\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__18952\,
            I => \N__18945\
        );

    \I__4088\ : InMux
    port map (
            O => \N__18951\,
            I => \N__18942\
        );

    \I__4087\ : Span12Mux_h
    port map (
            O => \N__18948\,
            I => \N__18939\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__18945\,
            I => \M_this_internal_address_qZ0Z_10\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__18942\,
            I => \M_this_internal_address_qZ0Z_10\
        );

    \I__4084\ : Odrv12
    port map (
            O => \N__18939\,
            I => \M_this_internal_address_qZ0Z_10\
        );

    \I__4083\ : InMux
    port map (
            O => \N__18932\,
            I => \N__18929\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__18929\,
            I => \N__18926\
        );

    \I__4081\ : Odrv4
    port map (
            O => \N__18926\,
            I => \M_this_internal_address_q_RNO_1Z0Z_10\
        );

    \I__4080\ : InMux
    port map (
            O => \N__18923\,
            I => \un1_M_this_internal_address_q_cry_9\
        );

    \I__4079\ : InMux
    port map (
            O => \N__18920\,
            I => \un1_M_this_internal_address_q_cry_10\
        );

    \I__4078\ : InMux
    port map (
            O => \N__18917\,
            I => \un1_M_this_internal_address_q_cry_11\
        );

    \I__4077\ : InMux
    port map (
            O => \N__18914\,
            I => \un1_M_this_internal_address_q_cry_12\
        );

    \I__4076\ : InMux
    port map (
            O => \N__18911\,
            I => \N__18908\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__18908\,
            I => \N__18905\
        );

    \I__4074\ : Span4Mux_h
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__18902\,
            I => \M_this_internal_address_q_RNO_1Z0Z_13\
        );

    \I__4072\ : CascadeMux
    port map (
            O => \N__18899\,
            I => \N__18896\
        );

    \I__4071\ : CascadeBuf
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__4070\ : CascadeMux
    port map (
            O => \N__18893\,
            I => \N__18890\
        );

    \I__4069\ : CascadeBuf
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__4068\ : CascadeMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__4067\ : CascadeBuf
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__4066\ : CascadeMux
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__4065\ : CascadeBuf
    port map (
            O => \N__18878\,
            I => \N__18875\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__4063\ : CascadeBuf
    port map (
            O => \N__18872\,
            I => \N__18869\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__4061\ : CascadeBuf
    port map (
            O => \N__18866\,
            I => \N__18863\
        );

    \I__4060\ : CascadeMux
    port map (
            O => \N__18863\,
            I => \N__18860\
        );

    \I__4059\ : CascadeBuf
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__18857\,
            I => \N__18854\
        );

    \I__4057\ : CascadeBuf
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__4056\ : CascadeMux
    port map (
            O => \N__18851\,
            I => \N__18848\
        );

    \I__4055\ : CascadeBuf
    port map (
            O => \N__18848\,
            I => \N__18845\
        );

    \I__4054\ : CascadeMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__4053\ : CascadeBuf
    port map (
            O => \N__18842\,
            I => \N__18839\
        );

    \I__4052\ : CascadeMux
    port map (
            O => \N__18839\,
            I => \N__18836\
        );

    \I__4051\ : CascadeBuf
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__4050\ : CascadeMux
    port map (
            O => \N__18833\,
            I => \N__18830\
        );

    \I__4049\ : CascadeBuf
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__4047\ : CascadeBuf
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__4046\ : CascadeMux
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__4045\ : CascadeBuf
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__4044\ : CascadeMux
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__4043\ : CascadeBuf
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__18809\,
            I => \N__18805\
        );

    \I__4041\ : InMux
    port map (
            O => \N__18808\,
            I => \N__18802\
        );

    \I__4040\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18798\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__18802\,
            I => \N__18795\
        );

    \I__4038\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18792\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__18798\,
            I => \N__18789\
        );

    \I__4036\ : Span4Mux_v
    port map (
            O => \N__18795\,
            I => \N__18784\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__18792\,
            I => \N__18784\
        );

    \I__4034\ : Span12Mux_h
    port map (
            O => \N__18789\,
            I => \N__18781\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__18784\,
            I => \M_this_internal_address_qZ0Z_7\
        );

    \I__4032\ : Odrv12
    port map (
            O => \N__18781\,
            I => \M_this_internal_address_qZ0Z_7\
        );

    \I__4031\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18773\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__18773\,
            I => \N__18770\
        );

    \I__4029\ : Odrv4
    port map (
            O => \N__18770\,
            I => \M_this_internal_address_q_3_ns_1_7\
        );

    \I__4028\ : IoInMux
    port map (
            O => \N__18767\,
            I => \N__18763\
        );

    \I__4027\ : IoInMux
    port map (
            O => \N__18766\,
            I => \N__18760\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__18763\,
            I => \N__18753\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__18760\,
            I => \N__18753\
        );

    \I__4024\ : IoInMux
    port map (
            O => \N__18759\,
            I => \N__18750\
        );

    \I__4023\ : IoInMux
    port map (
            O => \N__18758\,
            I => \N__18745\
        );

    \I__4022\ : IoSpan4Mux
    port map (
            O => \N__18753\,
            I => \N__18742\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__18750\,
            I => \N__18736\
        );

    \I__4020\ : IoInMux
    port map (
            O => \N__18749\,
            I => \N__18733\
        );

    \I__4019\ : IoInMux
    port map (
            O => \N__18748\,
            I => \N__18730\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__18745\,
            I => \N__18726\
        );

    \I__4017\ : IoSpan4Mux
    port map (
            O => \N__18742\,
            I => \N__18723\
        );

    \I__4016\ : IoInMux
    port map (
            O => \N__18741\,
            I => \N__18720\
        );

    \I__4015\ : IoInMux
    port map (
            O => \N__18740\,
            I => \N__18717\
        );

    \I__4014\ : IoInMux
    port map (
            O => \N__18739\,
            I => \N__18711\
        );

    \I__4013\ : IoSpan4Mux
    port map (
            O => \N__18736\,
            I => \N__18704\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__18733\,
            I => \N__18704\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__18730\,
            I => \N__18704\
        );

    \I__4010\ : IoInMux
    port map (
            O => \N__18729\,
            I => \N__18701\
        );

    \I__4009\ : IoSpan4Mux
    port map (
            O => \N__18726\,
            I => \N__18698\
        );

    \I__4008\ : IoSpan4Mux
    port map (
            O => \N__18723\,
            I => \N__18691\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__18720\,
            I => \N__18691\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__18717\,
            I => \N__18691\
        );

    \I__4005\ : IoInMux
    port map (
            O => \N__18716\,
            I => \N__18688\
        );

    \I__4004\ : IoInMux
    port map (
            O => \N__18715\,
            I => \N__18685\
        );

    \I__4003\ : IoInMux
    port map (
            O => \N__18714\,
            I => \N__18682\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__18711\,
            I => \N__18679\
        );

    \I__4001\ : IoSpan4Mux
    port map (
            O => \N__18704\,
            I => \N__18674\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__18701\,
            I => \N__18674\
        );

    \I__3999\ : Span4Mux_s3_h
    port map (
            O => \N__18698\,
            I => \N__18670\
        );

    \I__3998\ : IoSpan4Mux
    port map (
            O => \N__18691\,
            I => \N__18663\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__18688\,
            I => \N__18663\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__18685\,
            I => \N__18663\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__18682\,
            I => \N__18660\
        );

    \I__3994\ : Span4Mux_s3_h
    port map (
            O => \N__18679\,
            I => \N__18657\
        );

    \I__3993\ : IoSpan4Mux
    port map (
            O => \N__18674\,
            I => \N__18654\
        );

    \I__3992\ : IoInMux
    port map (
            O => \N__18673\,
            I => \N__18650\
        );

    \I__3991\ : Span4Mux_v
    port map (
            O => \N__18670\,
            I => \N__18643\
        );

    \I__3990\ : IoSpan4Mux
    port map (
            O => \N__18663\,
            I => \N__18643\
        );

    \I__3989\ : IoSpan4Mux
    port map (
            O => \N__18660\,
            I => \N__18643\
        );

    \I__3988\ : Sp12to4
    port map (
            O => \N__18657\,
            I => \N__18639\
        );

    \I__3987\ : Span4Mux_s1_v
    port map (
            O => \N__18654\,
            I => \N__18635\
        );

    \I__3986\ : IoInMux
    port map (
            O => \N__18653\,
            I => \N__18632\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__18650\,
            I => \N__18629\
        );

    \I__3984\ : Span4Mux_s3_h
    port map (
            O => \N__18643\,
            I => \N__18626\
        );

    \I__3983\ : IoInMux
    port map (
            O => \N__18642\,
            I => \N__18623\
        );

    \I__3982\ : Span12Mux_s9_v
    port map (
            O => \N__18639\,
            I => \N__18620\
        );

    \I__3981\ : IoInMux
    port map (
            O => \N__18638\,
            I => \N__18617\
        );

    \I__3980\ : Sp12to4
    port map (
            O => \N__18635\,
            I => \N__18612\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__18632\,
            I => \N__18612\
        );

    \I__3978\ : Span4Mux_s2_v
    port map (
            O => \N__18629\,
            I => \N__18609\
        );

    \I__3977\ : Span4Mux_h
    port map (
            O => \N__18626\,
            I => \N__18606\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__18623\,
            I => \N__18603\
        );

    \I__3975\ : Span12Mux_h
    port map (
            O => \N__18620\,
            I => \N__18598\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__18617\,
            I => \N__18598\
        );

    \I__3973\ : Span12Mux_s9_v
    port map (
            O => \N__18612\,
            I => \N__18595\
        );

    \I__3972\ : Span4Mux_v
    port map (
            O => \N__18609\,
            I => \N__18592\
        );

    \I__3971\ : Sp12to4
    port map (
            O => \N__18606\,
            I => \N__18585\
        );

    \I__3970\ : Span12Mux_s4_h
    port map (
            O => \N__18603\,
            I => \N__18585\
        );

    \I__3969\ : Span12Mux_s9_v
    port map (
            O => \N__18598\,
            I => \N__18585\
        );

    \I__3968\ : Odrv12
    port map (
            O => \N__18595\,
            I => \N_235_0_i\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__18592\,
            I => \N_235_0_i\
        );

    \I__3966\ : Odrv12
    port map (
            O => \N__18585\,
            I => \N_235_0_i\
        );

    \I__3965\ : InMux
    port map (
            O => \N__18578\,
            I => \un1_M_this_internal_address_q_cry_0\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__18575\,
            I => \N__18572\
        );

    \I__3963\ : CascadeBuf
    port map (
            O => \N__18572\,
            I => \N__18569\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__18569\,
            I => \N__18566\
        );

    \I__3961\ : CascadeBuf
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__3960\ : CascadeMux
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__3959\ : CascadeBuf
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__3957\ : CascadeBuf
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__3955\ : CascadeBuf
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__3954\ : CascadeMux
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__3953\ : CascadeBuf
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__3952\ : CascadeMux
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__3951\ : CascadeBuf
    port map (
            O => \N__18536\,
            I => \N__18533\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__3949\ : CascadeBuf
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__3948\ : CascadeMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__3947\ : CascadeBuf
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__3946\ : CascadeMux
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__3945\ : CascadeBuf
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__3944\ : CascadeMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__3943\ : CascadeBuf
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__3942\ : CascadeMux
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__3941\ : CascadeBuf
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__3939\ : CascadeBuf
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__3938\ : CascadeMux
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__3937\ : CascadeBuf
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__3936\ : CascadeMux
    port map (
            O => \N__18491\,
            I => \N__18488\
        );

    \I__3935\ : CascadeBuf
    port map (
            O => \N__18488\,
            I => \N__18485\
        );

    \I__3934\ : CascadeMux
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__3933\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__3931\ : Span4Mux_h
    port map (
            O => \N__18476\,
            I => \N__18473\
        );

    \I__3930\ : Sp12to4
    port map (
            O => \N__18473\,
            I => \N__18468\
        );

    \I__3929\ : InMux
    port map (
            O => \N__18472\,
            I => \N__18465\
        );

    \I__3928\ : InMux
    port map (
            O => \N__18471\,
            I => \N__18462\
        );

    \I__3927\ : Span12Mux_s11_v
    port map (
            O => \N__18468\,
            I => \N__18459\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__18465\,
            I => \M_this_internal_address_qZ0Z_2\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__18462\,
            I => \M_this_internal_address_qZ0Z_2\
        );

    \I__3924\ : Odrv12
    port map (
            O => \N__18459\,
            I => \M_this_internal_address_qZ0Z_2\
        );

    \I__3923\ : InMux
    port map (
            O => \N__18452\,
            I => \N__18449\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__18449\,
            I => \M_this_internal_address_q_RNO_1Z0Z_2\
        );

    \I__3921\ : InMux
    port map (
            O => \N__18446\,
            I => \un1_M_this_internal_address_q_cry_1\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__3919\ : CascadeBuf
    port map (
            O => \N__18440\,
            I => \N__18437\
        );

    \I__3918\ : CascadeMux
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__3917\ : CascadeBuf
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__3916\ : CascadeMux
    port map (
            O => \N__18431\,
            I => \N__18428\
        );

    \I__3915\ : CascadeBuf
    port map (
            O => \N__18428\,
            I => \N__18425\
        );

    \I__3914\ : CascadeMux
    port map (
            O => \N__18425\,
            I => \N__18422\
        );

    \I__3913\ : CascadeBuf
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__3911\ : CascadeBuf
    port map (
            O => \N__18416\,
            I => \N__18413\
        );

    \I__3910\ : CascadeMux
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__3909\ : CascadeBuf
    port map (
            O => \N__18410\,
            I => \N__18407\
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__18407\,
            I => \N__18404\
        );

    \I__3907\ : CascadeBuf
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__3906\ : CascadeMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__3905\ : CascadeBuf
    port map (
            O => \N__18398\,
            I => \N__18395\
        );

    \I__3904\ : CascadeMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__3903\ : CascadeBuf
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__3901\ : CascadeBuf
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__3900\ : CascadeMux
    port map (
            O => \N__18383\,
            I => \N__18380\
        );

    \I__3899\ : CascadeBuf
    port map (
            O => \N__18380\,
            I => \N__18377\
        );

    \I__3898\ : CascadeMux
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__3897\ : CascadeBuf
    port map (
            O => \N__18374\,
            I => \N__18371\
        );

    \I__3896\ : CascadeMux
    port map (
            O => \N__18371\,
            I => \N__18368\
        );

    \I__3895\ : CascadeBuf
    port map (
            O => \N__18368\,
            I => \N__18365\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__18365\,
            I => \N__18362\
        );

    \I__3893\ : CascadeBuf
    port map (
            O => \N__18362\,
            I => \N__18359\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__18359\,
            I => \N__18356\
        );

    \I__3891\ : CascadeBuf
    port map (
            O => \N__18356\,
            I => \N__18353\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__18353\,
            I => \N__18350\
        );

    \I__3889\ : InMux
    port map (
            O => \N__18350\,
            I => \N__18347\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__18347\,
            I => \N__18343\
        );

    \I__3887\ : InMux
    port map (
            O => \N__18346\,
            I => \N__18339\
        );

    \I__3886\ : Sp12to4
    port map (
            O => \N__18343\,
            I => \N__18336\
        );

    \I__3885\ : InMux
    port map (
            O => \N__18342\,
            I => \N__18333\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__18339\,
            I => \N__18328\
        );

    \I__3883\ : Span12Mux_s11_v
    port map (
            O => \N__18336\,
            I => \N__18328\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__18333\,
            I => \M_this_internal_address_qZ0Z_3\
        );

    \I__3881\ : Odrv12
    port map (
            O => \N__18328\,
            I => \M_this_internal_address_qZ0Z_3\
        );

    \I__3880\ : InMux
    port map (
            O => \N__18323\,
            I => \N__18320\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__18320\,
            I => \M_this_internal_address_q_RNO_1Z0Z_3\
        );

    \I__3878\ : InMux
    port map (
            O => \N__18317\,
            I => \un1_M_this_internal_address_q_cry_2\
        );

    \I__3877\ : InMux
    port map (
            O => \N__18314\,
            I => \un1_M_this_internal_address_q_cry_3\
        );

    \I__3876\ : InMux
    port map (
            O => \N__18311\,
            I => \un1_M_this_internal_address_q_cry_4\
        );

    \I__3875\ : InMux
    port map (
            O => \N__18308\,
            I => \un1_M_this_internal_address_q_cry_5\
        );

    \I__3874\ : InMux
    port map (
            O => \N__18305\,
            I => \N__18302\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__18302\,
            I => \N__18299\
        );

    \I__3872\ : Span4Mux_h
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__18296\,
            I => \M_this_internal_address_q_RNO_1Z0Z_7\
        );

    \I__3870\ : InMux
    port map (
            O => \N__18293\,
            I => \un1_M_this_internal_address_q_cry_6\
        );

    \I__3869\ : CascadeMux
    port map (
            O => \N__18290\,
            I => \this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_c3_0_cascade_\
        );

    \I__3868\ : InMux
    port map (
            O => \N__18287\,
            I => \N__18282\
        );

    \I__3867\ : InMux
    port map (
            O => \N__18286\,
            I => \N__18277\
        );

    \I__3866\ : InMux
    port map (
            O => \N__18285\,
            I => \N__18277\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__18282\,
            I => if_generate_plus_mult1_un89_sum_axbxc3
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__18277\,
            I => if_generate_plus_mult1_un89_sum_axbxc3
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__18272\,
            I => \this_ppu.sprites_N_7_0_cascade_\
        );

    \I__3862\ : InMux
    port map (
            O => \N__18269\,
            I => \N__18265\
        );

    \I__3861\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18262\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__18265\,
            I => \this_ppu.un5_sprites_addr_1_c2\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__18262\,
            I => \this_ppu.un5_sprites_addr_1_c2\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__18257\,
            I => \this_ppu.sprites_m7Z0Z_0_cascade_\
        );

    \I__3857\ : InMux
    port map (
            O => \N__18254\,
            I => \N__18251\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__18251\,
            I => \N__18241\
        );

    \I__3855\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18232\
        );

    \I__3854\ : InMux
    port map (
            O => \N__18249\,
            I => \N__18232\
        );

    \I__3853\ : InMux
    port map (
            O => \N__18248\,
            I => \N__18232\
        );

    \I__3852\ : InMux
    port map (
            O => \N__18247\,
            I => \N__18232\
        );

    \I__3851\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18229\
        );

    \I__3850\ : InMux
    port map (
            O => \N__18245\,
            I => \N__18224\
        );

    \I__3849\ : InMux
    port map (
            O => \N__18244\,
            I => \N__18224\
        );

    \I__3848\ : Odrv4
    port map (
            O => \N__18241\,
            I => if_generate_plus_mult1_un68_sum_axbxc3_ns
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__18232\,
            I => if_generate_plus_mult1_un68_sum_axbxc3_ns
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__18229\,
            I => if_generate_plus_mult1_un68_sum_axbxc3_ns
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__18224\,
            I => if_generate_plus_mult1_un68_sum_axbxc3_ns
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__18215\,
            I => \N__18212\
        );

    \I__3843\ : CascadeBuf
    port map (
            O => \N__18212\,
            I => \N__18209\
        );

    \I__3842\ : CascadeMux
    port map (
            O => \N__18209\,
            I => \N__18206\
        );

    \I__3841\ : CascadeBuf
    port map (
            O => \N__18206\,
            I => \N__18203\
        );

    \I__3840\ : CascadeMux
    port map (
            O => \N__18203\,
            I => \N__18200\
        );

    \I__3839\ : CascadeBuf
    port map (
            O => \N__18200\,
            I => \N__18197\
        );

    \I__3838\ : CascadeMux
    port map (
            O => \N__18197\,
            I => \N__18194\
        );

    \I__3837\ : CascadeBuf
    port map (
            O => \N__18194\,
            I => \N__18191\
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__18191\,
            I => \N__18188\
        );

    \I__3835\ : CascadeBuf
    port map (
            O => \N__18188\,
            I => \N__18185\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__18185\,
            I => \N__18182\
        );

    \I__3833\ : CascadeBuf
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__18179\,
            I => \N__18176\
        );

    \I__3831\ : CascadeBuf
    port map (
            O => \N__18176\,
            I => \N__18173\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__3829\ : CascadeBuf
    port map (
            O => \N__18170\,
            I => \N__18167\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__3827\ : CascadeBuf
    port map (
            O => \N__18164\,
            I => \N__18161\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__18161\,
            I => \N__18158\
        );

    \I__3825\ : CascadeBuf
    port map (
            O => \N__18158\,
            I => \N__18155\
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__3823\ : CascadeBuf
    port map (
            O => \N__18152\,
            I => \N__18149\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__18149\,
            I => \N__18146\
        );

    \I__3821\ : CascadeBuf
    port map (
            O => \N__18146\,
            I => \N__18143\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__18143\,
            I => \N__18140\
        );

    \I__3819\ : CascadeBuf
    port map (
            O => \N__18140\,
            I => \N__18137\
        );

    \I__3818\ : CascadeMux
    port map (
            O => \N__18137\,
            I => \N__18134\
        );

    \I__3817\ : CascadeBuf
    port map (
            O => \N__18134\,
            I => \N__18131\
        );

    \I__3816\ : CascadeMux
    port map (
            O => \N__18131\,
            I => \N__18128\
        );

    \I__3815\ : CascadeBuf
    port map (
            O => \N__18128\,
            I => \N__18125\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__18125\,
            I => \N__18122\
        );

    \I__3813\ : InMux
    port map (
            O => \N__18122\,
            I => \N__18119\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__18119\,
            I => \N__18116\
        );

    \I__3811\ : Span12Mux_s10_h
    port map (
            O => \N__18116\,
            I => \N__18113\
        );

    \I__3810\ : Span12Mux_v
    port map (
            O => \N__18113\,
            I => \N__18110\
        );

    \I__3809\ : Odrv12
    port map (
            O => \N__18110\,
            I => \N_140_i\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__18107\,
            I => \N__18102\
        );

    \I__3807\ : InMux
    port map (
            O => \N__18106\,
            I => \N__18094\
        );

    \I__3806\ : InMux
    port map (
            O => \N__18105\,
            I => \N__18090\
        );

    \I__3805\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18087\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__18101\,
            I => \N__18084\
        );

    \I__3803\ : InMux
    port map (
            O => \N__18100\,
            I => \N__18079\
        );

    \I__3802\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18076\
        );

    \I__3801\ : InMux
    port map (
            O => \N__18098\,
            I => \N__18071\
        );

    \I__3800\ : InMux
    port map (
            O => \N__18097\,
            I => \N__18071\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__18094\,
            I => \N__18068\
        );

    \I__3798\ : CascadeMux
    port map (
            O => \N__18093\,
            I => \N__18063\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__18090\,
            I => \N__18057\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__18087\,
            I => \N__18057\
        );

    \I__3795\ : InMux
    port map (
            O => \N__18084\,
            I => \N__18054\
        );

    \I__3794\ : InMux
    port map (
            O => \N__18083\,
            I => \N__18049\
        );

    \I__3793\ : InMux
    port map (
            O => \N__18082\,
            I => \N__18049\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__18079\,
            I => \N__18046\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__18076\,
            I => \N__18041\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__18071\,
            I => \N__18041\
        );

    \I__3789\ : Span12Mux_v
    port map (
            O => \N__18068\,
            I => \N__18038\
        );

    \I__3788\ : InMux
    port map (
            O => \N__18067\,
            I => \N__18035\
        );

    \I__3787\ : InMux
    port map (
            O => \N__18066\,
            I => \N__18032\
        );

    \I__3786\ : InMux
    port map (
            O => \N__18063\,
            I => \N__18027\
        );

    \I__3785\ : InMux
    port map (
            O => \N__18062\,
            I => \N__18027\
        );

    \I__3784\ : Span4Mux_v
    port map (
            O => \N__18057\,
            I => \N__18024\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__18054\,
            I => \N__18021\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__18049\,
            I => \N__18018\
        );

    \I__3781\ : Span4Mux_v
    port map (
            O => \N__18046\,
            I => \N__18013\
        );

    \I__3780\ : Span4Mux_h
    port map (
            O => \N__18041\,
            I => \N__18013\
        );

    \I__3779\ : Odrv12
    port map (
            O => \N__18038\,
            I => \this_vga_signals_M_hcounter_q_2\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__18035\,
            I => \this_vga_signals_M_hcounter_q_2\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__18032\,
            I => \this_vga_signals_M_hcounter_q_2\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__18027\,
            I => \this_vga_signals_M_hcounter_q_2\
        );

    \I__3775\ : Odrv4
    port map (
            O => \N__18024\,
            I => \this_vga_signals_M_hcounter_q_2\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__18021\,
            I => \this_vga_signals_M_hcounter_q_2\
        );

    \I__3773\ : Odrv12
    port map (
            O => \N__18018\,
            I => \this_vga_signals_M_hcounter_q_2\
        );

    \I__3772\ : Odrv4
    port map (
            O => \N__18013\,
            I => \this_vga_signals_M_hcounter_q_2\
        );

    \I__3771\ : InMux
    port map (
            O => \N__17996\,
            I => \N__17989\
        );

    \I__3770\ : InMux
    port map (
            O => \N__17995\,
            I => \N__17989\
        );

    \I__3769\ : InMux
    port map (
            O => \N__17994\,
            I => \N__17986\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__17989\,
            I => \N__17983\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__17986\,
            I => \N__17980\
        );

    \I__3766\ : Span4Mux_v
    port map (
            O => \N__17983\,
            I => \N__17974\
        );

    \I__3765\ : Span4Mux_h
    port map (
            O => \N__17980\,
            I => \N__17974\
        );

    \I__3764\ : InMux
    port map (
            O => \N__17979\,
            I => \N__17971\
        );

    \I__3763\ : Odrv4
    port map (
            O => \N__17974\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__17971\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1
        );

    \I__3761\ : InMux
    port map (
            O => \N__17966\,
            I => \N__17962\
        );

    \I__3760\ : InMux
    port map (
            O => \N__17965\,
            I => \N__17959\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__17962\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__17959\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3
        );

    \I__3757\ : InMux
    port map (
            O => \N__17954\,
            I => \N__17946\
        );

    \I__3756\ : InMux
    port map (
            O => \N__17953\,
            I => \N__17946\
        );

    \I__3755\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17941\
        );

    \I__3754\ : InMux
    port map (
            O => \N__17951\,
            I => \N__17941\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__17946\,
            I => if_generate_plus_mult1_un75_sum_axbxc3
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__17941\,
            I => if_generate_plus_mult1_un75_sum_axbxc3
        );

    \I__3751\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17930\
        );

    \I__3750\ : InMux
    port map (
            O => \N__17935\,
            I => \N__17920\
        );

    \I__3749\ : InMux
    port map (
            O => \N__17934\,
            I => \N__17920\
        );

    \I__3748\ : InMux
    port map (
            O => \N__17933\,
            I => \N__17920\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__17930\,
            I => \N__17917\
        );

    \I__3746\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17910\
        );

    \I__3745\ : InMux
    port map (
            O => \N__17928\,
            I => \N__17910\
        );

    \I__3744\ : InMux
    port map (
            O => \N__17927\,
            I => \N__17910\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__17920\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__17917\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__17910\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0
        );

    \I__3740\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17898\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__17902\,
            I => \N__17893\
        );

    \I__3738\ : InMux
    port map (
            O => \N__17901\,
            I => \N__17890\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__17898\,
            I => \N__17885\
        );

    \I__3736\ : InMux
    port map (
            O => \N__17897\,
            I => \N__17882\
        );

    \I__3735\ : InMux
    port map (
            O => \N__17896\,
            I => \N__17878\
        );

    \I__3734\ : InMux
    port map (
            O => \N__17893\,
            I => \N__17875\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__17890\,
            I => \N__17872\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__17889\,
            I => \N__17866\
        );

    \I__3731\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17862\
        );

    \I__3730\ : Span4Mux_h
    port map (
            O => \N__17885\,
            I => \N__17859\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__17882\,
            I => \N__17856\
        );

    \I__3728\ : InMux
    port map (
            O => \N__17881\,
            I => \N__17853\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__17878\,
            I => \N__17848\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__17875\,
            I => \N__17848\
        );

    \I__3725\ : Span4Mux_h
    port map (
            O => \N__17872\,
            I => \N__17845\
        );

    \I__3724\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17842\
        );

    \I__3723\ : InMux
    port map (
            O => \N__17870\,
            I => \N__17839\
        );

    \I__3722\ : InMux
    port map (
            O => \N__17869\,
            I => \N__17832\
        );

    \I__3721\ : InMux
    port map (
            O => \N__17866\,
            I => \N__17832\
        );

    \I__3720\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17832\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__17862\,
            I => \N__17829\
        );

    \I__3718\ : Span4Mux_v
    port map (
            O => \N__17859\,
            I => \N__17820\
        );

    \I__3717\ : Span4Mux_h
    port map (
            O => \N__17856\,
            I => \N__17820\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__17853\,
            I => \N__17820\
        );

    \I__3715\ : Span4Mux_h
    port map (
            O => \N__17848\,
            I => \N__17820\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__17845\,
            I => \this_vga_signals_M_hcounter_q_1\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__17842\,
            I => \this_vga_signals_M_hcounter_q_1\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__17839\,
            I => \this_vga_signals_M_hcounter_q_1\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__17832\,
            I => \this_vga_signals_M_hcounter_q_1\
        );

    \I__3710\ : Odrv12
    port map (
            O => \N__17829\,
            I => \this_vga_signals_M_hcounter_q_1\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__17820\,
            I => \this_vga_signals_M_hcounter_q_1\
        );

    \I__3708\ : CascadeMux
    port map (
            O => \N__17807\,
            I => \N__17804\
        );

    \I__3707\ : InMux
    port map (
            O => \N__17804\,
            I => \N__17796\
        );

    \I__3706\ : InMux
    port map (
            O => \N__17803\,
            I => \N__17792\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__17802\,
            I => \N__17789\
        );

    \I__3704\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17785\
        );

    \I__3703\ : CascadeMux
    port map (
            O => \N__17800\,
            I => \N__17782\
        );

    \I__3702\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17779\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__17796\,
            I => \N__17776\
        );

    \I__3700\ : CascadeMux
    port map (
            O => \N__17795\,
            I => \N__17770\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__17792\,
            I => \N__17767\
        );

    \I__3698\ : InMux
    port map (
            O => \N__17789\,
            I => \N__17762\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17788\,
            I => \N__17762\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__17785\,
            I => \N__17759\
        );

    \I__3695\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17756\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__17779\,
            I => \N__17751\
        );

    \I__3693\ : Span4Mux_v
    port map (
            O => \N__17776\,
            I => \N__17751\
        );

    \I__3692\ : InMux
    port map (
            O => \N__17775\,
            I => \N__17746\
        );

    \I__3691\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17746\
        );

    \I__3690\ : InMux
    port map (
            O => \N__17773\,
            I => \N__17743\
        );

    \I__3689\ : InMux
    port map (
            O => \N__17770\,
            I => \N__17740\
        );

    \I__3688\ : Span4Mux_h
    port map (
            O => \N__17767\,
            I => \N__17735\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__17762\,
            I => \N__17735\
        );

    \I__3686\ : Span4Mux_v
    port map (
            O => \N__17759\,
            I => \N__17728\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__17756\,
            I => \N__17728\
        );

    \I__3684\ : Span4Mux_h
    port map (
            O => \N__17751\,
            I => \N__17728\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__17746\,
            I => \this_vga_signals_M_hcounter_q_0\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__17743\,
            I => \this_vga_signals_M_hcounter_q_0\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__17740\,
            I => \this_vga_signals_M_hcounter_q_0\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__17735\,
            I => \this_vga_signals_M_hcounter_q_0\
        );

    \I__3679\ : Odrv4
    port map (
            O => \N__17728\,
            I => \this_vga_signals_M_hcounter_q_0\
        );

    \I__3678\ : CascadeMux
    port map (
            O => \N__17717\,
            I => \this_ppu.sprites_mZ0Z1_cascade_\
        );

    \I__3677\ : InMux
    port map (
            O => \N__17714\,
            I => \N__17709\
        );

    \I__3676\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17704\
        );

    \I__3675\ : InMux
    port map (
            O => \N__17712\,
            I => \N__17704\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__17709\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axb1
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__17704\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axb1
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__17699\,
            I => \M_this_internal_address_q_3_ns_1_10_cascade_\
        );

    \I__3671\ : SRMux
    port map (
            O => \N__17696\,
            I => \N__17692\
        );

    \I__3670\ : SRMux
    port map (
            O => \N__17695\,
            I => \N__17689\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__17692\,
            I => \N__17686\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__17689\,
            I => \N__17683\
        );

    \I__3667\ : Span4Mux_h
    port map (
            O => \N__17686\,
            I => \N__17680\
        );

    \I__3666\ : Odrv4
    port map (
            O => \N__17683\,
            I => \M_this_state_q_RNI20CEZ0Z_0\
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__17680\,
            I => \M_this_state_q_RNI20CEZ0Z_0\
        );

    \I__3664\ : SRMux
    port map (
            O => \N__17675\,
            I => \N__17668\
        );

    \I__3663\ : SRMux
    port map (
            O => \N__17674\,
            I => \N__17665\
        );

    \I__3662\ : SRMux
    port map (
            O => \N__17673\,
            I => \N__17662\
        );

    \I__3661\ : SRMux
    port map (
            O => \N__17672\,
            I => \N__17655\
        );

    \I__3660\ : SRMux
    port map (
            O => \N__17671\,
            I => \N__17652\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__17668\,
            I => \N__17649\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__17665\,
            I => \N__17644\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__17662\,
            I => \N__17644\
        );

    \I__3656\ : SRMux
    port map (
            O => \N__17661\,
            I => \N__17641\
        );

    \I__3655\ : SRMux
    port map (
            O => \N__17660\,
            I => \N__17638\
        );

    \I__3654\ : SRMux
    port map (
            O => \N__17659\,
            I => \N__17632\
        );

    \I__3653\ : SRMux
    port map (
            O => \N__17658\,
            I => \N__17626\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__17655\,
            I => \N__17623\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__17652\,
            I => \N__17620\
        );

    \I__3650\ : Span4Mux_h
    port map (
            O => \N__17649\,
            I => \N__17611\
        );

    \I__3649\ : Span4Mux_s3_v
    port map (
            O => \N__17644\,
            I => \N__17611\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__17641\,
            I => \N__17611\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__17638\,
            I => \N__17611\
        );

    \I__3646\ : SRMux
    port map (
            O => \N__17637\,
            I => \N__17608\
        );

    \I__3645\ : SRMux
    port map (
            O => \N__17636\,
            I => \N__17605\
        );

    \I__3644\ : SRMux
    port map (
            O => \N__17635\,
            I => \N__17599\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__17632\,
            I => \N__17595\
        );

    \I__3642\ : SRMux
    port map (
            O => \N__17631\,
            I => \N__17592\
        );

    \I__3641\ : SRMux
    port map (
            O => \N__17630\,
            I => \N__17586\
        );

    \I__3640\ : SRMux
    port map (
            O => \N__17629\,
            I => \N__17581\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__17626\,
            I => \N__17578\
        );

    \I__3638\ : Span4Mux_v
    port map (
            O => \N__17623\,
            I => \N__17567\
        );

    \I__3637\ : Span4Mux_h
    port map (
            O => \N__17620\,
            I => \N__17567\
        );

    \I__3636\ : Span4Mux_v
    port map (
            O => \N__17611\,
            I => \N__17567\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__17608\,
            I => \N__17567\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__17605\,
            I => \N__17567\
        );

    \I__3633\ : SRMux
    port map (
            O => \N__17604\,
            I => \N__17564\
        );

    \I__3632\ : SRMux
    port map (
            O => \N__17603\,
            I => \N__17561\
        );

    \I__3631\ : IoInMux
    port map (
            O => \N__17602\,
            I => \N__17556\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__17599\,
            I => \N__17553\
        );

    \I__3629\ : SRMux
    port map (
            O => \N__17598\,
            I => \N__17550\
        );

    \I__3628\ : Span4Mux_v
    port map (
            O => \N__17595\,
            I => \N__17544\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__17592\,
            I => \N__17544\
        );

    \I__3626\ : SRMux
    port map (
            O => \N__17591\,
            I => \N__17541\
        );

    \I__3625\ : SRMux
    port map (
            O => \N__17590\,
            I => \N__17537\
        );

    \I__3624\ : SRMux
    port map (
            O => \N__17589\,
            I => \N__17534\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__17586\,
            I => \N__17530\
        );

    \I__3622\ : SRMux
    port map (
            O => \N__17585\,
            I => \N__17527\
        );

    \I__3621\ : SRMux
    port map (
            O => \N__17584\,
            I => \N__17524\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__17581\,
            I => \N__17519\
        );

    \I__3619\ : Span4Mux_h
    port map (
            O => \N__17578\,
            I => \N__17510\
        );

    \I__3618\ : Span4Mux_v
    port map (
            O => \N__17567\,
            I => \N__17510\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__17564\,
            I => \N__17510\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__17561\,
            I => \N__17510\
        );

    \I__3615\ : SRMux
    port map (
            O => \N__17560\,
            I => \N__17507\
        );

    \I__3614\ : SRMux
    port map (
            O => \N__17559\,
            I => \N__17504\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__17556\,
            I => \N__17499\
        );

    \I__3612\ : Span4Mux_v
    port map (
            O => \N__17553\,
            I => \N__17496\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__17550\,
            I => \N__17493\
        );

    \I__3610\ : SRMux
    port map (
            O => \N__17549\,
            I => \N__17489\
        );

    \I__3609\ : Span4Mux_v
    port map (
            O => \N__17544\,
            I => \N__17484\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__17541\,
            I => \N__17484\
        );

    \I__3607\ : SRMux
    port map (
            O => \N__17540\,
            I => \N__17481\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__17537\,
            I => \N__17478\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__17534\,
            I => \N__17475\
        );

    \I__3604\ : SRMux
    port map (
            O => \N__17533\,
            I => \N__17472\
        );

    \I__3603\ : Span4Mux_h
    port map (
            O => \N__17530\,
            I => \N__17465\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__17527\,
            I => \N__17465\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__17524\,
            I => \N__17465\
        );

    \I__3600\ : SRMux
    port map (
            O => \N__17523\,
            I => \N__17462\
        );

    \I__3599\ : SRMux
    port map (
            O => \N__17522\,
            I => \N__17459\
        );

    \I__3598\ : Span4Mux_h
    port map (
            O => \N__17519\,
            I => \N__17449\
        );

    \I__3597\ : Span4Mux_v
    port map (
            O => \N__17510\,
            I => \N__17449\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__17507\,
            I => \N__17449\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__17504\,
            I => \N__17449\
        );

    \I__3594\ : SRMux
    port map (
            O => \N__17503\,
            I => \N__17446\
        );

    \I__3593\ : SRMux
    port map (
            O => \N__17502\,
            I => \N__17443\
        );

    \I__3592\ : IoSpan4Mux
    port map (
            O => \N__17499\,
            I => \N__17440\
        );

    \I__3591\ : Span4Mux_v
    port map (
            O => \N__17496\,
            I => \N__17435\
        );

    \I__3590\ : Span4Mux_v
    port map (
            O => \N__17493\,
            I => \N__17435\
        );

    \I__3589\ : SRMux
    port map (
            O => \N__17492\,
            I => \N__17431\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__17489\,
            I => \N__17428\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__17484\,
            I => \N__17423\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__17481\,
            I => \N__17423\
        );

    \I__3585\ : Span4Mux_v
    port map (
            O => \N__17478\,
            I => \N__17416\
        );

    \I__3584\ : Span4Mux_h
    port map (
            O => \N__17475\,
            I => \N__17416\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__17472\,
            I => \N__17416\
        );

    \I__3582\ : Span4Mux_v
    port map (
            O => \N__17465\,
            I => \N__17409\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__17462\,
            I => \N__17409\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__17459\,
            I => \N__17409\
        );

    \I__3579\ : SRMux
    port map (
            O => \N__17458\,
            I => \N__17406\
        );

    \I__3578\ : Span4Mux_v
    port map (
            O => \N__17449\,
            I => \N__17399\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__17446\,
            I => \N__17399\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__17443\,
            I => \N__17399\
        );

    \I__3575\ : Span4Mux_s3_h
    port map (
            O => \N__17440\,
            I => \N__17396\
        );

    \I__3574\ : Span4Mux_h
    port map (
            O => \N__17435\,
            I => \N__17393\
        );

    \I__3573\ : InMux
    port map (
            O => \N__17434\,
            I => \N__17390\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__17431\,
            I => \N__17387\
        );

    \I__3571\ : Span4Mux_h
    port map (
            O => \N__17428\,
            I => \N__17384\
        );

    \I__3570\ : Span4Mux_v
    port map (
            O => \N__17423\,
            I => \N__17379\
        );

    \I__3569\ : Span4Mux_v
    port map (
            O => \N__17416\,
            I => \N__17379\
        );

    \I__3568\ : Span4Mux_v
    port map (
            O => \N__17409\,
            I => \N__17372\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__17406\,
            I => \N__17372\
        );

    \I__3566\ : Span4Mux_v
    port map (
            O => \N__17399\,
            I => \N__17372\
        );

    \I__3565\ : Span4Mux_h
    port map (
            O => \N__17396\,
            I => \N__17369\
        );

    \I__3564\ : Span4Mux_v
    port map (
            O => \N__17393\,
            I => \N__17364\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__17390\,
            I => \N__17364\
        );

    \I__3562\ : Span12Mux_s11_v
    port map (
            O => \N__17387\,
            I => \N__17361\
        );

    \I__3561\ : Span4Mux_v
    port map (
            O => \N__17384\,
            I => \N__17354\
        );

    \I__3560\ : Span4Mux_h
    port map (
            O => \N__17379\,
            I => \N__17354\
        );

    \I__3559\ : Span4Mux_h
    port map (
            O => \N__17372\,
            I => \N__17354\
        );

    \I__3558\ : Span4Mux_h
    port map (
            O => \N__17369\,
            I => \N__17349\
        );

    \I__3557\ : Span4Mux_v
    port map (
            O => \N__17364\,
            I => \N__17349\
        );

    \I__3556\ : Span12Mux_v
    port map (
            O => \N__17361\,
            I => \N__17343\
        );

    \I__3555\ : Span4Mux_h
    port map (
            O => \N__17354\,
            I => \N__17340\
        );

    \I__3554\ : Span4Mux_v
    port map (
            O => \N__17349\,
            I => \N__17337\
        );

    \I__3553\ : InMux
    port map (
            O => \N__17348\,
            I => \N__17334\
        );

    \I__3552\ : InMux
    port map (
            O => \N__17347\,
            I => \N__17329\
        );

    \I__3551\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17329\
        );

    \I__3550\ : Odrv12
    port map (
            O => \N__17343\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3549\ : Odrv4
    port map (
            O => \N__17340\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3548\ : Odrv4
    port map (
            O => \N__17337\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__17334\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__17329\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3545\ : InMux
    port map (
            O => \N__17318\,
            I => \bfn_15_25_0_\
        );

    \I__3544\ : InMux
    port map (
            O => \N__17315\,
            I => \N__17312\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__17312\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__17309\,
            I => \N__17306\
        );

    \I__3541\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17303\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__17303\,
            I => \N__17299\
        );

    \I__3539\ : CascadeMux
    port map (
            O => \N__17302\,
            I => \N__17296\
        );

    \I__3538\ : Span4Mux_h
    port map (
            O => \N__17299\,
            I => \N__17293\
        );

    \I__3537\ : InMux
    port map (
            O => \N__17296\,
            I => \N__17290\
        );

    \I__3536\ : Span4Mux_v
    port map (
            O => \N__17293\,
            I => \N__17287\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__17290\,
            I => \N__17284\
        );

    \I__3534\ : Span4Mux_v
    port map (
            O => \N__17287\,
            I => \N__17281\
        );

    \I__3533\ : Span4Mux_h
    port map (
            O => \N__17284\,
            I => \N__17278\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__17281\,
            I => \N_13_0\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__17278\,
            I => \N_13_0\
        );

    \I__3530\ : InMux
    port map (
            O => \N__17273\,
            I => \N__17267\
        );

    \I__3529\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17267\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__17267\,
            I => \M_this_vga_signals_address_5\
        );

    \I__3527\ : InMux
    port map (
            O => \N__17264\,
            I => \N__17260\
        );

    \I__3526\ : InMux
    port map (
            O => \N__17263\,
            I => \N__17257\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__17260\,
            I => \this_ppu.un5_sprites_addr_1_c4\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__17257\,
            I => \this_ppu.un5_sprites_addr_1_c4\
        );

    \I__3523\ : InMux
    port map (
            O => \N__17252\,
            I => \un1_M_this_data_count_q_cry_3\
        );

    \I__3522\ : InMux
    port map (
            O => \N__17249\,
            I => \un1_M_this_data_count_q_cry_4\
        );

    \I__3521\ : InMux
    port map (
            O => \N__17246\,
            I => \un1_M_this_data_count_q_cry_5\
        );

    \I__3520\ : InMux
    port map (
            O => \N__17243\,
            I => \un1_M_this_data_count_q_cry_6\
        );

    \I__3519\ : InMux
    port map (
            O => \N__17240\,
            I => \bfn_15_24_0_\
        );

    \I__3518\ : InMux
    port map (
            O => \N__17237\,
            I => \un1_M_this_data_count_q_cry_8\
        );

    \I__3517\ : InMux
    port map (
            O => \N__17234\,
            I => \un1_M_this_data_count_q_cry_9\
        );

    \I__3516\ : InMux
    port map (
            O => \N__17231\,
            I => \un1_M_this_data_count_q_cry_10\
        );

    \I__3515\ : InMux
    port map (
            O => \N__17228\,
            I => \un1_M_this_data_count_q_cry_11\
        );

    \I__3514\ : InMux
    port map (
            O => \N__17225\,
            I => \N__17222\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__17222\,
            I => \M_this_internal_address_q_3_ns_1_9\
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__17219\,
            I => \M_this_internal_address_q_3_ns_1_3_cascade_\
        );

    \I__3511\ : InMux
    port map (
            O => \N__17216\,
            I => \N__17213\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__17213\,
            I => \M_this_internal_address_q_3_ns_1_8\
        );

    \I__3509\ : InMux
    port map (
            O => \N__17210\,
            I => \un1_M_this_data_count_q_cry_0\
        );

    \I__3508\ : InMux
    port map (
            O => \N__17207\,
            I => \un1_M_this_data_count_q_cry_1\
        );

    \I__3507\ : InMux
    port map (
            O => \N__17204\,
            I => \un1_M_this_data_count_q_cry_2\
        );

    \I__3506\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17195\
        );

    \I__3505\ : InMux
    port map (
            O => \N__17200\,
            I => \N__17195\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__17195\,
            I => \N__17191\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__17194\,
            I => \N__17187\
        );

    \I__3502\ : Span4Mux_h
    port map (
            O => \N__17191\,
            I => \N__17184\
        );

    \I__3501\ : InMux
    port map (
            O => \N__17190\,
            I => \N__17179\
        );

    \I__3500\ : InMux
    port map (
            O => \N__17187\,
            I => \N__17179\
        );

    \I__3499\ : Odrv4
    port map (
            O => \N__17184\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_c3
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__17179\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_c3
        );

    \I__3497\ : InMux
    port map (
            O => \N__17174\,
            I => \N__17165\
        );

    \I__3496\ : InMux
    port map (
            O => \N__17173\,
            I => \N__17165\
        );

    \I__3495\ : InMux
    port map (
            O => \N__17172\,
            I => \N__17160\
        );

    \I__3494\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17160\
        );

    \I__3493\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17157\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__17165\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__17160\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__17157\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0
        );

    \I__3489\ : InMux
    port map (
            O => \N__17150\,
            I => \N__17133\
        );

    \I__3488\ : InMux
    port map (
            O => \N__17149\,
            I => \N__17133\
        );

    \I__3487\ : InMux
    port map (
            O => \N__17148\,
            I => \N__17133\
        );

    \I__3486\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17128\
        );

    \I__3485\ : InMux
    port map (
            O => \N__17146\,
            I => \N__17128\
        );

    \I__3484\ : InMux
    port map (
            O => \N__17145\,
            I => \N__17123\
        );

    \I__3483\ : InMux
    port map (
            O => \N__17144\,
            I => \N__17123\
        );

    \I__3482\ : InMux
    port map (
            O => \N__17143\,
            I => \N__17120\
        );

    \I__3481\ : InMux
    port map (
            O => \N__17142\,
            I => \N__17111\
        );

    \I__3480\ : InMux
    port map (
            O => \N__17141\,
            I => \N__17111\
        );

    \I__3479\ : InMux
    port map (
            O => \N__17140\,
            I => \N__17111\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__17133\,
            I => \N__17108\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__17128\,
            I => \N__17103\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__17123\,
            I => \N__17103\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__17120\,
            I => \N__17100\
        );

    \I__3474\ : InMux
    port map (
            O => \N__17119\,
            I => \N__17095\
        );

    \I__3473\ : InMux
    port map (
            O => \N__17118\,
            I => \N__17095\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__17111\,
            I => \N__17092\
        );

    \I__3471\ : Span4Mux_v
    port map (
            O => \N__17108\,
            I => \N__17087\
        );

    \I__3470\ : Span4Mux_h
    port map (
            O => \N__17103\,
            I => \N__17087\
        );

    \I__3469\ : Span12Mux_v
    port map (
            O => \N__17100\,
            I => \N__17083\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__17095\,
            I => \N__17080\
        );

    \I__3467\ : Span4Mux_h
    port map (
            O => \N__17092\,
            I => \N__17077\
        );

    \I__3466\ : Span4Mux_h
    port map (
            O => \N__17087\,
            I => \N__17074\
        );

    \I__3465\ : InMux
    port map (
            O => \N__17086\,
            I => \N__17071\
        );

    \I__3464\ : Span12Mux_h
    port map (
            O => \N__17083\,
            I => \N__17068\
        );

    \I__3463\ : Odrv12
    port map (
            O => \N__17080\,
            I => \this_vga_signals.GZ0Z_210\
        );

    \I__3462\ : Odrv4
    port map (
            O => \N__17077\,
            I => \this_vga_signals.GZ0Z_210\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__17074\,
            I => \this_vga_signals.GZ0Z_210\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__17071\,
            I => \this_vga_signals.GZ0Z_210\
        );

    \I__3459\ : Odrv12
    port map (
            O => \N__17068\,
            I => \this_vga_signals.GZ0Z_210\
        );

    \I__3458\ : SRMux
    port map (
            O => \N__17057\,
            I => \N__17051\
        );

    \I__3457\ : SRMux
    port map (
            O => \N__17056\,
            I => \N__17048\
        );

    \I__3456\ : SRMux
    port map (
            O => \N__17055\,
            I => \N__17045\
        );

    \I__3455\ : SRMux
    port map (
            O => \N__17054\,
            I => \N__17042\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__17051\,
            I => \N__17039\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__17048\,
            I => \N__17036\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__17045\,
            I => \N__17033\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__17042\,
            I => \N__17030\
        );

    \I__3450\ : Span4Mux_v
    port map (
            O => \N__17039\,
            I => \N__17026\
        );

    \I__3449\ : Span4Mux_h
    port map (
            O => \N__17036\,
            I => \N__17021\
        );

    \I__3448\ : Span4Mux_v
    port map (
            O => \N__17033\,
            I => \N__17021\
        );

    \I__3447\ : Span4Mux_v
    port map (
            O => \N__17030\,
            I => \N__17018\
        );

    \I__3446\ : InMux
    port map (
            O => \N__17029\,
            I => \N__17015\
        );

    \I__3445\ : Odrv4
    port map (
            O => \N__17026\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI4UBI1Z0Z_9\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__17021\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI4UBI1Z0Z_9\
        );

    \I__3443\ : Odrv4
    port map (
            O => \N__17018\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI4UBI1Z0Z_9\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__17015\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI4UBI1Z0Z_9\
        );

    \I__3441\ : InMux
    port map (
            O => \N__17006\,
            I => \N__17003\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__17003\,
            I => \N__16997\
        );

    \I__3439\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16993\
        );

    \I__3438\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16989\
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__17000\,
            I => \N__16983\
        );

    \I__3436\ : Span4Mux_v
    port map (
            O => \N__16997\,
            I => \N__16980\
        );

    \I__3435\ : InMux
    port map (
            O => \N__16996\,
            I => \N__16977\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__16993\,
            I => \N__16974\
        );

    \I__3433\ : InMux
    port map (
            O => \N__16992\,
            I => \N__16971\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__16989\,
            I => \N__16968\
        );

    \I__3431\ : InMux
    port map (
            O => \N__16988\,
            I => \N__16964\
        );

    \I__3430\ : InMux
    port map (
            O => \N__16987\,
            I => \N__16961\
        );

    \I__3429\ : InMux
    port map (
            O => \N__16986\,
            I => \N__16956\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16983\,
            I => \N__16956\
        );

    \I__3427\ : Span4Mux_h
    port map (
            O => \N__16980\,
            I => \N__16948\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__16977\,
            I => \N__16948\
        );

    \I__3425\ : Span4Mux_v
    port map (
            O => \N__16974\,
            I => \N__16948\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__16971\,
            I => \N__16943\
        );

    \I__3423\ : Span4Mux_v
    port map (
            O => \N__16968\,
            I => \N__16943\
        );

    \I__3422\ : InMux
    port map (
            O => \N__16967\,
            I => \N__16940\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__16964\,
            I => \N__16935\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__16961\,
            I => \N__16935\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__16956\,
            I => \N__16932\
        );

    \I__3418\ : InMux
    port map (
            O => \N__16955\,
            I => \N__16929\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__16948\,
            I => \this_vga_signals_M_hcounter_q_3\
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__16943\,
            I => \this_vga_signals_M_hcounter_q_3\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__16940\,
            I => \this_vga_signals_M_hcounter_q_3\
        );

    \I__3414\ : Odrv4
    port map (
            O => \N__16935\,
            I => \this_vga_signals_M_hcounter_q_3\
        );

    \I__3413\ : Odrv12
    port map (
            O => \N__16932\,
            I => \this_vga_signals_M_hcounter_q_3\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__16929\,
            I => \this_vga_signals_M_hcounter_q_3\
        );

    \I__3411\ : InMux
    port map (
            O => \N__16916\,
            I => \N__16913\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__16913\,
            I => \this_vga_signals.if_N_9_1\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16907\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__16907\,
            I => \this_ppu.sprites_m1_0_xZ0Z1\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__16904\,
            I => \this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3_cascade_\
        );

    \I__3406\ : InMux
    port map (
            O => \N__16901\,
            I => \N__16898\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__16898\,
            I => \this_ppu.sprites_m1_0_xZ0Z0\
        );

    \I__3404\ : InMux
    port map (
            O => \N__16895\,
            I => \N__16892\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__16892\,
            I => \M_this_internal_address_q_3_ns_1_2\
        );

    \I__3402\ : InMux
    port map (
            O => \N__16889\,
            I => \N__16884\
        );

    \I__3401\ : InMux
    port map (
            O => \N__16888\,
            I => \N__16879\
        );

    \I__3400\ : InMux
    port map (
            O => \N__16887\,
            I => \N__16879\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__16884\,
            I => \this_pixel_clk.M_counter_qZ0Z_0\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__16879\,
            I => \this_pixel_clk.M_counter_qZ0Z_0\
        );

    \I__3397\ : InMux
    port map (
            O => \N__16874\,
            I => \N__16871\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__16871\,
            I => \N__16864\
        );

    \I__3395\ : InMux
    port map (
            O => \N__16870\,
            I => \N__16861\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__16869\,
            I => \N__16857\
        );

    \I__3393\ : CascadeMux
    port map (
            O => \N__16868\,
            I => \N__16854\
        );

    \I__3392\ : InMux
    port map (
            O => \N__16867\,
            I => \N__16850\
        );

    \I__3391\ : Span4Mux_h
    port map (
            O => \N__16864\,
            I => \N__16845\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__16861\,
            I => \N__16845\
        );

    \I__3389\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16842\
        );

    \I__3388\ : InMux
    port map (
            O => \N__16857\,
            I => \N__16835\
        );

    \I__3387\ : InMux
    port map (
            O => \N__16854\,
            I => \N__16835\
        );

    \I__3386\ : InMux
    port map (
            O => \N__16853\,
            I => \N__16835\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__16850\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__3384\ : Odrv4
    port map (
            O => \N__16845\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__16842\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__16835\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__3381\ : CascadeMux
    port map (
            O => \N__16826\,
            I => \if_generate_plus_mult1_un75_sum_axbxc3_cascade_\
        );

    \I__3380\ : CascadeMux
    port map (
            O => \N__16823\,
            I => \this_ppu.un5_sprites_addr_1_c2_cascade_\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__16820\,
            I => \N__16817\
        );

    \I__3378\ : InMux
    port map (
            O => \N__16817\,
            I => \N__16812\
        );

    \I__3377\ : InMux
    port map (
            O => \N__16816\,
            I => \N__16809\
        );

    \I__3376\ : InMux
    port map (
            O => \N__16815\,
            I => \N__16806\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__16812\,
            I => \N__16803\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__16809\,
            I => \N__16800\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__16806\,
            I => \this_ppu.N_4_0_1\
        );

    \I__3372\ : Odrv4
    port map (
            O => \N__16803\,
            I => \this_ppu.N_4_0_1\
        );

    \I__3371\ : Odrv4
    port map (
            O => \N__16800\,
            I => \this_ppu.N_4_0_1\
        );

    \I__3370\ : InMux
    port map (
            O => \N__16793\,
            I => \N__16790\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__16790\,
            I => \this_ppu.sprites_addr_1_i_7_tz_0_9\
        );

    \I__3368\ : InMux
    port map (
            O => \N__16787\,
            I => \N__16784\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__16784\,
            I => \N__16781\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__16781\,
            I => \this_ppu.sprites_addr_1_i_a7Z0Z_9\
        );

    \I__3365\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16775\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__16775\,
            I => \N__16770\
        );

    \I__3363\ : InMux
    port map (
            O => \N__16774\,
            I => \N__16765\
        );

    \I__3362\ : InMux
    port map (
            O => \N__16773\,
            I => \N__16765\
        );

    \I__3361\ : Span4Mux_h
    port map (
            O => \N__16770\,
            I => \N__16759\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__16765\,
            I => \N__16756\
        );

    \I__3359\ : InMux
    port map (
            O => \N__16764\,
            I => \N__16753\
        );

    \I__3358\ : InMux
    port map (
            O => \N__16763\,
            I => \N__16748\
        );

    \I__3357\ : InMux
    port map (
            O => \N__16762\,
            I => \N__16748\
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__16759\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__16756\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__16753\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__16748\,
            I => this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__16739\,
            I => \N__16736\
        );

    \I__3351\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16733\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__16733\,
            I => \this_ppu.un5_sprites_addr1_4\
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__16730\,
            I => \this_vga_signals.if_N_8_i_0_cascade_\
        );

    \I__3348\ : InMux
    port map (
            O => \N__16727\,
            I => \N__16722\
        );

    \I__3347\ : InMux
    port map (
            O => \N__16726\,
            I => \N__16717\
        );

    \I__3346\ : InMux
    port map (
            O => \N__16725\,
            I => \N__16717\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__16722\,
            I => \this_vga_signals.mult1_un68_sum_axb1_1\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__16717\,
            I => \this_vga_signals.mult1_un68_sum_axb1_1\
        );

    \I__3343\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16709\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__16709\,
            I => \M_counter_q_RNIFKS8_0\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__16706\,
            I => \M_counter_q_RNIFKS8_0_cascade_\
        );

    \I__3340\ : InMux
    port map (
            O => \N__16703\,
            I => \N__16691\
        );

    \I__3339\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16691\
        );

    \I__3338\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16691\
        );

    \I__3337\ : InMux
    port map (
            O => \N__16700\,
            I => \N__16691\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__16691\,
            I => \this_pixel_clk_M_counter_q_i_1\
        );

    \I__3335\ : InMux
    port map (
            O => \N__16688\,
            I => \N__16685\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__16685\,
            I => \this_vga_signals.N_455\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__16682\,
            I => \N__16679\
        );

    \I__3332\ : InMux
    port map (
            O => \N__16679\,
            I => \N__16675\
        );

    \I__3331\ : InMux
    port map (
            O => \N__16678\,
            I => \N__16672\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__16675\,
            I => \N__16669\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__16672\,
            I => \N__16666\
        );

    \I__3328\ : Span4Mux_h
    port map (
            O => \N__16669\,
            I => \N__16663\
        );

    \I__3327\ : Span4Mux_h
    port map (
            O => \N__16666\,
            I => \N__16656\
        );

    \I__3326\ : Span4Mux_h
    port map (
            O => \N__16663\,
            I => \N__16656\
        );

    \I__3325\ : InMux
    port map (
            O => \N__16662\,
            I => \N__16651\
        );

    \I__3324\ : InMux
    port map (
            O => \N__16661\,
            I => \N__16651\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__16656\,
            I => \this_vga_signals.N_459\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__16651\,
            I => \this_vga_signals.N_459\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__16646\,
            I => \this_vga_signals.GZ0Z_210_cascade_\
        );

    \I__3320\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16634\
        );

    \I__3319\ : InMux
    port map (
            O => \N__16642\,
            I => \N__16631\
        );

    \I__3318\ : InMux
    port map (
            O => \N__16641\,
            I => \N__16627\
        );

    \I__3317\ : InMux
    port map (
            O => \N__16640\,
            I => \N__16624\
        );

    \I__3316\ : InMux
    port map (
            O => \N__16639\,
            I => \N__16621\
        );

    \I__3315\ : InMux
    port map (
            O => \N__16638\,
            I => \N__16616\
        );

    \I__3314\ : InMux
    port map (
            O => \N__16637\,
            I => \N__16616\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__16634\,
            I => \N__16608\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__16631\,
            I => \N__16605\
        );

    \I__3311\ : InMux
    port map (
            O => \N__16630\,
            I => \N__16602\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__16627\,
            I => \N__16599\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__16624\,
            I => \N__16592\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__16621\,
            I => \N__16592\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__16616\,
            I => \N__16592\
        );

    \I__3306\ : CascadeMux
    port map (
            O => \N__16615\,
            I => \N__16589\
        );

    \I__3305\ : CascadeMux
    port map (
            O => \N__16614\,
            I => \N__16585\
        );

    \I__3304\ : InMux
    port map (
            O => \N__16613\,
            I => \N__16582\
        );

    \I__3303\ : InMux
    port map (
            O => \N__16612\,
            I => \N__16578\
        );

    \I__3302\ : InMux
    port map (
            O => \N__16611\,
            I => \N__16575\
        );

    \I__3301\ : Span4Mux_v
    port map (
            O => \N__16608\,
            I => \N__16572\
        );

    \I__3300\ : Span12Mux_s9_h
    port map (
            O => \N__16605\,
            I => \N__16569\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__16602\,
            I => \N__16562\
        );

    \I__3298\ : Span4Mux_h
    port map (
            O => \N__16599\,
            I => \N__16562\
        );

    \I__3297\ : Span4Mux_v
    port map (
            O => \N__16592\,
            I => \N__16562\
        );

    \I__3296\ : InMux
    port map (
            O => \N__16589\,
            I => \N__16555\
        );

    \I__3295\ : InMux
    port map (
            O => \N__16588\,
            I => \N__16555\
        );

    \I__3294\ : InMux
    port map (
            O => \N__16585\,
            I => \N__16555\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__16582\,
            I => \N__16552\
        );

    \I__3292\ : InMux
    port map (
            O => \N__16581\,
            I => \N__16549\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__16578\,
            I => \N__16544\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__16575\,
            I => \N__16544\
        );

    \I__3289\ : Odrv4
    port map (
            O => \N__16572\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3288\ : Odrv12
    port map (
            O => \N__16569\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3287\ : Odrv4
    port map (
            O => \N__16562\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__16555\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3285\ : Odrv4
    port map (
            O => \N__16552\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__16549\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__16544\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3282\ : IoInMux
    port map (
            O => \N__16529\,
            I => \N__16526\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__3280\ : IoSpan4Mux
    port map (
            O => \N__16523\,
            I => \N__16520\
        );

    \I__3279\ : Span4Mux_s0_h
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__3278\ : Sp12to4
    port map (
            O => \N__16517\,
            I => \N__16514\
        );

    \I__3277\ : Span12Mux_s8_h
    port map (
            O => \N__16514\,
            I => \N__16511\
        );

    \I__3276\ : Odrv12
    port map (
            O => \N__16511\,
            I => \this_vga_signals.M_vcounter_q_esr_RNIIRV75Z0Z_9\
        );

    \I__3275\ : InMux
    port map (
            O => \N__16508\,
            I => \N__16505\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__3273\ : Odrv4
    port map (
            O => \N__16502\,
            I => \this_ppu.sprites_addr_1_i_2_1Z0Z_9\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__16499\,
            I => \this_ppu.sprites_addr_1_i_0_0Z0Z_9_cascade_\
        );

    \I__3271\ : InMux
    port map (
            O => \N__16496\,
            I => \N__16493\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__16493\,
            I => \N__16490\
        );

    \I__3269\ : Span4Mux_h
    port map (
            O => \N__16490\,
            I => \N__16487\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__16487\,
            I => \this_ppu.sprites_addr_1_i_a0_2Z0Z_9\
        );

    \I__3267\ : CascadeMux
    port map (
            O => \N__16484\,
            I => \this_ppu.sprites_addr_1_i_0_2Z0Z_9_cascade_\
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__16481\,
            I => \N__16478\
        );

    \I__3265\ : CascadeBuf
    port map (
            O => \N__16478\,
            I => \N__16475\
        );

    \I__3264\ : CascadeMux
    port map (
            O => \N__16475\,
            I => \N__16472\
        );

    \I__3263\ : CascadeBuf
    port map (
            O => \N__16472\,
            I => \N__16469\
        );

    \I__3262\ : CascadeMux
    port map (
            O => \N__16469\,
            I => \N__16466\
        );

    \I__3261\ : CascadeBuf
    port map (
            O => \N__16466\,
            I => \N__16463\
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__16463\,
            I => \N__16460\
        );

    \I__3259\ : CascadeBuf
    port map (
            O => \N__16460\,
            I => \N__16457\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__16457\,
            I => \N__16454\
        );

    \I__3257\ : CascadeBuf
    port map (
            O => \N__16454\,
            I => \N__16451\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__16451\,
            I => \N__16448\
        );

    \I__3255\ : CascadeBuf
    port map (
            O => \N__16448\,
            I => \N__16445\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__16445\,
            I => \N__16442\
        );

    \I__3253\ : CascadeBuf
    port map (
            O => \N__16442\,
            I => \N__16439\
        );

    \I__3252\ : CascadeMux
    port map (
            O => \N__16439\,
            I => \N__16436\
        );

    \I__3251\ : CascadeBuf
    port map (
            O => \N__16436\,
            I => \N__16433\
        );

    \I__3250\ : CascadeMux
    port map (
            O => \N__16433\,
            I => \N__16430\
        );

    \I__3249\ : CascadeBuf
    port map (
            O => \N__16430\,
            I => \N__16427\
        );

    \I__3248\ : CascadeMux
    port map (
            O => \N__16427\,
            I => \N__16424\
        );

    \I__3247\ : CascadeBuf
    port map (
            O => \N__16424\,
            I => \N__16421\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__16421\,
            I => \N__16418\
        );

    \I__3245\ : CascadeBuf
    port map (
            O => \N__16418\,
            I => \N__16415\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__16415\,
            I => \N__16412\
        );

    \I__3243\ : CascadeBuf
    port map (
            O => \N__16412\,
            I => \N__16409\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__16409\,
            I => \N__16406\
        );

    \I__3241\ : CascadeBuf
    port map (
            O => \N__16406\,
            I => \N__16403\
        );

    \I__3240\ : CascadeMux
    port map (
            O => \N__16403\,
            I => \N__16400\
        );

    \I__3239\ : CascadeBuf
    port map (
            O => \N__16400\,
            I => \N__16397\
        );

    \I__3238\ : CascadeMux
    port map (
            O => \N__16397\,
            I => \N__16394\
        );

    \I__3237\ : CascadeBuf
    port map (
            O => \N__16394\,
            I => \N__16391\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__16391\,
            I => \N__16388\
        );

    \I__3235\ : InMux
    port map (
            O => \N__16388\,
            I => \N__16385\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__16385\,
            I => \N__16382\
        );

    \I__3233\ : Span12Mux_h
    port map (
            O => \N__16382\,
            I => \N__16379\
        );

    \I__3232\ : Span12Mux_v
    port map (
            O => \N__16379\,
            I => \N__16376\
        );

    \I__3231\ : Odrv12
    port map (
            O => \N__16376\,
            I => \N_138_0\
        );

    \I__3230\ : InMux
    port map (
            O => \N__16373\,
            I => \N__16370\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__16370\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_0_1\
        );

    \I__3228\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16364\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__16364\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_x0\
        );

    \I__3226\ : InMux
    port map (
            O => \N__16361\,
            I => \N__16358\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__16358\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_x1\
        );

    \I__3224\ : InMux
    port map (
            O => \N__16355\,
            I => \N__16352\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__16352\,
            I => \this_vga_signals.mult1_un75_sum_ac0_1\
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__16349\,
            I => \if_generate_plus_mult1_un68_sum_axbxc3_ns_cascade_\
        );

    \I__3221\ : CascadeMux
    port map (
            O => \N__16346\,
            I => \this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_cascade_\
        );

    \I__3220\ : InMux
    port map (
            O => \N__16343\,
            I => \N__16339\
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__16342\,
            I => \N__16335\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__16339\,
            I => \N__16332\
        );

    \I__3217\ : InMux
    port map (
            O => \N__16338\,
            I => \N__16329\
        );

    \I__3216\ : InMux
    port map (
            O => \N__16335\,
            I => \N__16326\
        );

    \I__3215\ : Span4Mux_h
    port map (
            O => \N__16332\,
            I => \N__16323\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__16329\,
            I => \N__16320\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__16326\,
            I => \N__16311\
        );

    \I__3212\ : Span4Mux_v
    port map (
            O => \N__16323\,
            I => \N__16304\
        );

    \I__3211\ : Span4Mux_h
    port map (
            O => \N__16320\,
            I => \N__16304\
        );

    \I__3210\ : InMux
    port map (
            O => \N__16319\,
            I => \N__16301\
        );

    \I__3209\ : InMux
    port map (
            O => \N__16318\,
            I => \N__16292\
        );

    \I__3208\ : InMux
    port map (
            O => \N__16317\,
            I => \N__16292\
        );

    \I__3207\ : InMux
    port map (
            O => \N__16316\,
            I => \N__16292\
        );

    \I__3206\ : InMux
    port map (
            O => \N__16315\,
            I => \N__16292\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__16314\,
            I => \N__16287\
        );

    \I__3204\ : Span4Mux_v
    port map (
            O => \N__16311\,
            I => \N__16281\
        );

    \I__3203\ : InMux
    port map (
            O => \N__16310\,
            I => \N__16278\
        );

    \I__3202\ : InMux
    port map (
            O => \N__16309\,
            I => \N__16275\
        );

    \I__3201\ : Span4Mux_h
    port map (
            O => \N__16304\,
            I => \N__16268\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__16301\,
            I => \N__16268\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__16292\,
            I => \N__16268\
        );

    \I__3198\ : InMux
    port map (
            O => \N__16291\,
            I => \N__16257\
        );

    \I__3197\ : InMux
    port map (
            O => \N__16290\,
            I => \N__16257\
        );

    \I__3196\ : InMux
    port map (
            O => \N__16287\,
            I => \N__16257\
        );

    \I__3195\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16257\
        );

    \I__3194\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16257\
        );

    \I__3193\ : InMux
    port map (
            O => \N__16284\,
            I => \N__16254\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__16281\,
            I => \this_vga_signals_M_hcounter_q_5\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__16278\,
            I => \this_vga_signals_M_hcounter_q_5\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__16275\,
            I => \this_vga_signals_M_hcounter_q_5\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__16268\,
            I => \this_vga_signals_M_hcounter_q_5\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__16257\,
            I => \this_vga_signals_M_hcounter_q_5\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__16254\,
            I => \this_vga_signals_M_hcounter_q_5\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__16241\,
            I => \N__16237\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__16240\,
            I => \N__16234\
        );

    \I__3184\ : InMux
    port map (
            O => \N__16237\,
            I => \N__16230\
        );

    \I__3183\ : InMux
    port map (
            O => \N__16234\,
            I => \N__16225\
        );

    \I__3182\ : InMux
    port map (
            O => \N__16233\,
            I => \N__16225\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__16230\,
            I => \this_vga_signals.mult1_un54_sum_axb1_0\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__16225\,
            I => \this_vga_signals.mult1_un54_sum_axb1_0\
        );

    \I__3179\ : InMux
    port map (
            O => \N__16220\,
            I => \N__16217\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__16217\,
            I => \N__16211\
        );

    \I__3177\ : InMux
    port map (
            O => \N__16216\,
            I => \N__16208\
        );

    \I__3176\ : InMux
    port map (
            O => \N__16215\,
            I => \N__16199\
        );

    \I__3175\ : InMux
    port map (
            O => \N__16214\,
            I => \N__16194\
        );

    \I__3174\ : Span4Mux_h
    port map (
            O => \N__16211\,
            I => \N__16191\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__16208\,
            I => \N__16188\
        );

    \I__3172\ : InMux
    port map (
            O => \N__16207\,
            I => \N__16185\
        );

    \I__3171\ : InMux
    port map (
            O => \N__16206\,
            I => \N__16182\
        );

    \I__3170\ : InMux
    port map (
            O => \N__16205\,
            I => \N__16179\
        );

    \I__3169\ : InMux
    port map (
            O => \N__16204\,
            I => \N__16172\
        );

    \I__3168\ : InMux
    port map (
            O => \N__16203\,
            I => \N__16172\
        );

    \I__3167\ : InMux
    port map (
            O => \N__16202\,
            I => \N__16172\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__16199\,
            I => \N__16164\
        );

    \I__3165\ : InMux
    port map (
            O => \N__16198\,
            I => \N__16161\
        );

    \I__3164\ : InMux
    port map (
            O => \N__16197\,
            I => \N__16158\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__16194\,
            I => \N__16155\
        );

    \I__3162\ : Span4Mux_h
    port map (
            O => \N__16191\,
            I => \N__16148\
        );

    \I__3161\ : Span4Mux_h
    port map (
            O => \N__16188\,
            I => \N__16148\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__16185\,
            I => \N__16148\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__16182\,
            I => \N__16141\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__16179\,
            I => \N__16141\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__16172\,
            I => \N__16141\
        );

    \I__3156\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16130\
        );

    \I__3155\ : InMux
    port map (
            O => \N__16170\,
            I => \N__16130\
        );

    \I__3154\ : InMux
    port map (
            O => \N__16169\,
            I => \N__16130\
        );

    \I__3153\ : InMux
    port map (
            O => \N__16168\,
            I => \N__16130\
        );

    \I__3152\ : InMux
    port map (
            O => \N__16167\,
            I => \N__16130\
        );

    \I__3151\ : Odrv4
    port map (
            O => \N__16164\,
            I => \this_vga_signals_M_hcounter_q_4\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__16161\,
            I => \this_vga_signals_M_hcounter_q_4\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__16158\,
            I => \this_vga_signals_M_hcounter_q_4\
        );

    \I__3148\ : Odrv12
    port map (
            O => \N__16155\,
            I => \this_vga_signals_M_hcounter_q_4\
        );

    \I__3147\ : Odrv4
    port map (
            O => \N__16148\,
            I => \this_vga_signals_M_hcounter_q_4\
        );

    \I__3146\ : Odrv4
    port map (
            O => \N__16141\,
            I => \this_vga_signals_M_hcounter_q_4\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__16130\,
            I => \this_vga_signals_M_hcounter_q_4\
        );

    \I__3144\ : InMux
    port map (
            O => \N__16115\,
            I => \this_vga_signals.un1_M_hcounter_d_1_cry_2\
        );

    \I__3143\ : InMux
    port map (
            O => \N__16112\,
            I => \this_vga_signals.un1_M_hcounter_d_1_cry_3\
        );

    \I__3142\ : InMux
    port map (
            O => \N__16109\,
            I => \this_vga_signals.un1_M_hcounter_d_1_cry_4\
        );

    \I__3141\ : InMux
    port map (
            O => \N__16106\,
            I => \this_vga_signals.un1_M_hcounter_d_1_cry_5\
        );

    \I__3140\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16097\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__16102\,
            I => \N__16094\
        );

    \I__3138\ : InMux
    port map (
            O => \N__16101\,
            I => \N__16089\
        );

    \I__3137\ : InMux
    port map (
            O => \N__16100\,
            I => \N__16086\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__16097\,
            I => \N__16082\
        );

    \I__3135\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16077\
        );

    \I__3134\ : InMux
    port map (
            O => \N__16093\,
            I => \N__16077\
        );

    \I__3133\ : InMux
    port map (
            O => \N__16092\,
            I => \N__16074\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__16089\,
            I => \N__16069\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__16086\,
            I => \N__16069\
        );

    \I__3130\ : InMux
    port map (
            O => \N__16085\,
            I => \N__16066\
        );

    \I__3129\ : Span4Mux_v
    port map (
            O => \N__16082\,
            I => \N__16057\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__16077\,
            I => \N__16057\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__16074\,
            I => \N__16053\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__16069\,
            I => \N__16048\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__16066\,
            I => \N__16048\
        );

    \I__3124\ : InMux
    port map (
            O => \N__16065\,
            I => \N__16045\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__16064\,
            I => \N__16042\
        );

    \I__3122\ : CascadeMux
    port map (
            O => \N__16063\,
            I => \N__16039\
        );

    \I__3121\ : InMux
    port map (
            O => \N__16062\,
            I => \N__16036\
        );

    \I__3120\ : Span4Mux_h
    port map (
            O => \N__16057\,
            I => \N__16033\
        );

    \I__3119\ : InMux
    port map (
            O => \N__16056\,
            I => \N__16030\
        );

    \I__3118\ : Span4Mux_v
    port map (
            O => \N__16053\,
            I => \N__16023\
        );

    \I__3117\ : Span4Mux_h
    port map (
            O => \N__16048\,
            I => \N__16023\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__16045\,
            I => \N__16023\
        );

    \I__3115\ : InMux
    port map (
            O => \N__16042\,
            I => \N__16018\
        );

    \I__3114\ : InMux
    port map (
            O => \N__16039\,
            I => \N__16018\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__16036\,
            I => \this_vga_signals_M_hcounter_q_7\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__16033\,
            I => \this_vga_signals_M_hcounter_q_7\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__16030\,
            I => \this_vga_signals_M_hcounter_q_7\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__16023\,
            I => \this_vga_signals_M_hcounter_q_7\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__16018\,
            I => \this_vga_signals_M_hcounter_q_7\
        );

    \I__3108\ : InMux
    port map (
            O => \N__16007\,
            I => \this_vga_signals.un1_M_hcounter_d_1_cry_6\
        );

    \I__3107\ : CascadeMux
    port map (
            O => \N__16004\,
            I => \N__15999\
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__16003\,
            I => \N__15996\
        );

    \I__3105\ : InMux
    port map (
            O => \N__16002\,
            I => \N__15993\
        );

    \I__3104\ : InMux
    port map (
            O => \N__15999\,
            I => \N__15988\
        );

    \I__3103\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15985\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__15993\,
            I => \N__15980\
        );

    \I__3101\ : InMux
    port map (
            O => \N__15992\,
            I => \N__15977\
        );

    \I__3100\ : InMux
    port map (
            O => \N__15991\,
            I => \N__15973\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__15988\,
            I => \N__15968\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__15985\,
            I => \N__15968\
        );

    \I__3097\ : InMux
    port map (
            O => \N__15984\,
            I => \N__15965\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__15983\,
            I => \N__15962\
        );

    \I__3095\ : Span4Mux_v
    port map (
            O => \N__15980\,
            I => \N__15954\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__15977\,
            I => \N__15954\
        );

    \I__3093\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15951\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__15973\,
            I => \N__15948\
        );

    \I__3091\ : Span4Mux_v
    port map (
            O => \N__15968\,
            I => \N__15943\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__15965\,
            I => \N__15943\
        );

    \I__3089\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15940\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15935\
        );

    \I__3087\ : InMux
    port map (
            O => \N__15960\,
            I => \N__15932\
        );

    \I__3086\ : InMux
    port map (
            O => \N__15959\,
            I => \N__15929\
        );

    \I__3085\ : Span4Mux_h
    port map (
            O => \N__15954\,
            I => \N__15924\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__15951\,
            I => \N__15924\
        );

    \I__3083\ : Span4Mux_v
    port map (
            O => \N__15948\,
            I => \N__15917\
        );

    \I__3082\ : Span4Mux_h
    port map (
            O => \N__15943\,
            I => \N__15917\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__15940\,
            I => \N__15917\
        );

    \I__3080\ : InMux
    port map (
            O => \N__15939\,
            I => \N__15914\
        );

    \I__3079\ : InMux
    port map (
            O => \N__15938\,
            I => \N__15911\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__15935\,
            I => \this_vga_signals_M_hcounter_q_8\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__15932\,
            I => \this_vga_signals_M_hcounter_q_8\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__15929\,
            I => \this_vga_signals_M_hcounter_q_8\
        );

    \I__3075\ : Odrv4
    port map (
            O => \N__15924\,
            I => \this_vga_signals_M_hcounter_q_8\
        );

    \I__3074\ : Odrv4
    port map (
            O => \N__15917\,
            I => \this_vga_signals_M_hcounter_q_8\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__15914\,
            I => \this_vga_signals_M_hcounter_q_8\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__15911\,
            I => \this_vga_signals_M_hcounter_q_8\
        );

    \I__3071\ : InMux
    port map (
            O => \N__15896\,
            I => \this_vga_signals.un1_M_hcounter_d_1_cry_7\
        );

    \I__3070\ : InMux
    port map (
            O => \N__15893\,
            I => \bfn_14_18_0_\
        );

    \I__3069\ : InMux
    port map (
            O => \N__15890\,
            I => \N__15885\
        );

    \I__3068\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15882\
        );

    \I__3067\ : InMux
    port map (
            O => \N__15888\,
            I => \N__15879\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__15885\,
            I => \N__15870\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__15882\,
            I => \N__15870\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__15879\,
            I => \N__15867\
        );

    \I__3063\ : InMux
    port map (
            O => \N__15878\,
            I => \N__15864\
        );

    \I__3062\ : InMux
    port map (
            O => \N__15877\,
            I => \N__15860\
        );

    \I__3061\ : InMux
    port map (
            O => \N__15876\,
            I => \N__15857\
        );

    \I__3060\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15854\
        );

    \I__3059\ : Span4Mux_v
    port map (
            O => \N__15870\,
            I => \N__15847\
        );

    \I__3058\ : Span4Mux_v
    port map (
            O => \N__15867\,
            I => \N__15847\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__15864\,
            I => \N__15847\
        );

    \I__3056\ : InMux
    port map (
            O => \N__15863\,
            I => \N__15841\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__15860\,
            I => \N__15838\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__15857\,
            I => \N__15833\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__15854\,
            I => \N__15833\
        );

    \I__3052\ : Span4Mux_h
    port map (
            O => \N__15847\,
            I => \N__15830\
        );

    \I__3051\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15827\
        );

    \I__3050\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15824\
        );

    \I__3049\ : InMux
    port map (
            O => \N__15844\,
            I => \N__15821\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__15841\,
            I => \this_vga_signals_M_hcounter_q_9\
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__15838\,
            I => \this_vga_signals_M_hcounter_q_9\
        );

    \I__3046\ : Odrv4
    port map (
            O => \N__15833\,
            I => \this_vga_signals_M_hcounter_q_9\
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__15830\,
            I => \this_vga_signals_M_hcounter_q_9\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__15827\,
            I => \this_vga_signals_M_hcounter_q_9\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__15824\,
            I => \this_vga_signals_M_hcounter_q_9\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__15821\,
            I => \this_vga_signals_M_hcounter_q_9\
        );

    \I__3041\ : InMux
    port map (
            O => \N__15806\,
            I => \N__15802\
        );

    \I__3040\ : InMux
    port map (
            O => \N__15805\,
            I => \N__15799\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__15802\,
            I => \this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUFZ0\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__15799\,
            I => \this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUFZ0\
        );

    \I__3037\ : InMux
    port map (
            O => \N__15794\,
            I => \N__15785\
        );

    \I__3036\ : InMux
    port map (
            O => \N__15793\,
            I => \N__15785\
        );

    \I__3035\ : InMux
    port map (
            O => \N__15792\,
            I => \N__15782\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__15791\,
            I => \N__15778\
        );

    \I__3033\ : InMux
    port map (
            O => \N__15790\,
            I => \N__15775\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__15785\,
            I => \N__15769\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__15782\,
            I => \N__15769\
        );

    \I__3030\ : InMux
    port map (
            O => \N__15781\,
            I => \N__15760\
        );

    \I__3029\ : InMux
    port map (
            O => \N__15778\,
            I => \N__15760\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__15775\,
            I => \N__15757\
        );

    \I__3027\ : InMux
    port map (
            O => \N__15774\,
            I => \N__15754\
        );

    \I__3026\ : Span4Mux_v
    port map (
            O => \N__15769\,
            I => \N__15751\
        );

    \I__3025\ : InMux
    port map (
            O => \N__15768\,
            I => \N__15748\
        );

    \I__3024\ : CascadeMux
    port map (
            O => \N__15767\,
            I => \N__15745\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__15766\,
            I => \N__15742\
        );

    \I__3022\ : InMux
    port map (
            O => \N__15765\,
            I => \N__15739\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__15760\,
            I => \N__15736\
        );

    \I__3020\ : Span4Mux_v
    port map (
            O => \N__15757\,
            I => \N__15731\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__15754\,
            I => \N__15731\
        );

    \I__3018\ : Span4Mux_h
    port map (
            O => \N__15751\,
            I => \N__15726\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__15748\,
            I => \N__15726\
        );

    \I__3016\ : InMux
    port map (
            O => \N__15745\,
            I => \N__15723\
        );

    \I__3015\ : InMux
    port map (
            O => \N__15742\,
            I => \N__15720\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__15739\,
            I => \this_vga_signals_M_hcounter_q_6\
        );

    \I__3013\ : Odrv4
    port map (
            O => \N__15736\,
            I => \this_vga_signals_M_hcounter_q_6\
        );

    \I__3012\ : Odrv4
    port map (
            O => \N__15731\,
            I => \this_vga_signals_M_hcounter_q_6\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__15726\,
            I => \this_vga_signals_M_hcounter_q_6\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__15723\,
            I => \this_vga_signals_M_hcounter_q_6\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__15720\,
            I => \this_vga_signals_M_hcounter_q_6\
        );

    \I__3008\ : CEMux
    port map (
            O => \N__15707\,
            I => \N__15703\
        );

    \I__3007\ : CEMux
    port map (
            O => \N__15706\,
            I => \N__15700\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__15703\,
            I => \N__15697\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__15700\,
            I => \N__15694\
        );

    \I__3004\ : Span4Mux_h
    port map (
            O => \N__15697\,
            I => \N__15691\
        );

    \I__3003\ : Odrv4
    port map (
            O => \N__15694\,
            I => \this_vga_signals.N_517_0\
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__15691\,
            I => \this_vga_signals.N_517_0\
        );

    \I__3001\ : InMux
    port map (
            O => \N__15686\,
            I => \N__15682\
        );

    \I__3000\ : InMux
    port map (
            O => \N__15685\,
            I => \N__15679\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__15682\,
            I => \this_vga_signals.mult1_un61_sum_axbxc1\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__15679\,
            I => \this_vga_signals.mult1_un61_sum_axbxc1\
        );

    \I__2997\ : InMux
    port map (
            O => \N__15674\,
            I => \N__15671\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__15671\,
            I => \N__15668\
        );

    \I__2995\ : Odrv12
    port map (
            O => \N__15668\,
            I => \this_vga_signals.N_3\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__15665\,
            I => \N__15662\
        );

    \I__2993\ : InMux
    port map (
            O => \N__15662\,
            I => \N__15658\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__15661\,
            I => \N__15654\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__15658\,
            I => \N__15651\
        );

    \I__2990\ : InMux
    port map (
            O => \N__15657\,
            I => \N__15646\
        );

    \I__2989\ : InMux
    port map (
            O => \N__15654\,
            I => \N__15646\
        );

    \I__2988\ : Span4Mux_h
    port map (
            O => \N__15651\,
            I => \N__15643\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__15646\,
            I => \N__15640\
        );

    \I__2986\ : Sp12to4
    port map (
            O => \N__15643\,
            I => \N__15636\
        );

    \I__2985\ : Span4Mux_h
    port map (
            O => \N__15640\,
            I => \N__15633\
        );

    \I__2984\ : InMux
    port map (
            O => \N__15639\,
            I => \N__15630\
        );

    \I__2983\ : Odrv12
    port map (
            O => \N__15636\,
            I => \this_vga_signals.mult1_un68_sum_s_3\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__15633\,
            I => \this_vga_signals.mult1_un68_sum_s_3\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__15630\,
            I => \this_vga_signals.mult1_un68_sum_s_3\
        );

    \I__2980\ : ClkMux
    port map (
            O => \N__15623\,
            I => \N__15617\
        );

    \I__2979\ : ClkMux
    port map (
            O => \N__15622\,
            I => \N__15614\
        );

    \I__2978\ : ClkMux
    port map (
            O => \N__15621\,
            I => \N__15610\
        );

    \I__2977\ : ClkMux
    port map (
            O => \N__15620\,
            I => \N__15606\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__15617\,
            I => \N__15601\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__15614\,
            I => \N__15601\
        );

    \I__2974\ : ClkMux
    port map (
            O => \N__15613\,
            I => \N__15598\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__15610\,
            I => \N__15595\
        );

    \I__2972\ : ClkMux
    port map (
            O => \N__15609\,
            I => \N__15592\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__15606\,
            I => \N__15589\
        );

    \I__2970\ : IoSpan4Mux
    port map (
            O => \N__15601\,
            I => \N__15586\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__15598\,
            I => \N__15583\
        );

    \I__2968\ : Span4Mux_s2_h
    port map (
            O => \N__15595\,
            I => \N__15580\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__15592\,
            I => \N__15577\
        );

    \I__2966\ : Span4Mux_s2_h
    port map (
            O => \N__15589\,
            I => \N__15574\
        );

    \I__2965\ : IoSpan4Mux
    port map (
            O => \N__15586\,
            I => \N__15569\
        );

    \I__2964\ : IoSpan4Mux
    port map (
            O => \N__15583\,
            I => \N__15569\
        );

    \I__2963\ : Span4Mux_v
    port map (
            O => \N__15580\,
            I => \N__15566\
        );

    \I__2962\ : Span4Mux_s2_h
    port map (
            O => \N__15577\,
            I => \N__15563\
        );

    \I__2961\ : Sp12to4
    port map (
            O => \N__15574\,
            I => \N__15560\
        );

    \I__2960\ : Span4Mux_s1_h
    port map (
            O => \N__15569\,
            I => \N__15557\
        );

    \I__2959\ : Sp12to4
    port map (
            O => \N__15566\,
            I => \N__15552\
        );

    \I__2958\ : Sp12to4
    port map (
            O => \N__15563\,
            I => \N__15552\
        );

    \I__2957\ : Span12Mux_v
    port map (
            O => \N__15560\,
            I => \N__15545\
        );

    \I__2956\ : Sp12to4
    port map (
            O => \N__15557\,
            I => \N__15545\
        );

    \I__2955\ : Span12Mux_v
    port map (
            O => \N__15552\,
            I => \N__15545\
        );

    \I__2954\ : Odrv12
    port map (
            O => \N__15545\,
            I => \M_this_vga_signals_pixel_clk_0\
        );

    \I__2953\ : InMux
    port map (
            O => \N__15542\,
            I => \N__15539\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__15539\,
            I => \N__15534\
        );

    \I__2951\ : InMux
    port map (
            O => \N__15538\,
            I => \N__15529\
        );

    \I__2950\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15529\
        );

    \I__2949\ : Odrv12
    port map (
            O => \N__15534\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__15529\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__2947\ : CEMux
    port map (
            O => \N__15524\,
            I => \N__15503\
        );

    \I__2946\ : CEMux
    port map (
            O => \N__15523\,
            I => \N__15503\
        );

    \I__2945\ : CEMux
    port map (
            O => \N__15522\,
            I => \N__15503\
        );

    \I__2944\ : CEMux
    port map (
            O => \N__15521\,
            I => \N__15503\
        );

    \I__2943\ : CEMux
    port map (
            O => \N__15520\,
            I => \N__15503\
        );

    \I__2942\ : CEMux
    port map (
            O => \N__15519\,
            I => \N__15503\
        );

    \I__2941\ : CEMux
    port map (
            O => \N__15518\,
            I => \N__15503\
        );

    \I__2940\ : GlobalMux
    port map (
            O => \N__15503\,
            I => \N__15500\
        );

    \I__2939\ : gio2CtrlBuf
    port map (
            O => \N__15500\,
            I => \this_vga_signals.N_517_1_g\
        );

    \I__2938\ : InMux
    port map (
            O => \N__15497\,
            I => \N__15494\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__15494\,
            I => \N__15483\
        );

    \I__2936\ : SRMux
    port map (
            O => \N__15493\,
            I => \N__15464\
        );

    \I__2935\ : SRMux
    port map (
            O => \N__15492\,
            I => \N__15464\
        );

    \I__2934\ : SRMux
    port map (
            O => \N__15491\,
            I => \N__15464\
        );

    \I__2933\ : SRMux
    port map (
            O => \N__15490\,
            I => \N__15464\
        );

    \I__2932\ : SRMux
    port map (
            O => \N__15489\,
            I => \N__15464\
        );

    \I__2931\ : SRMux
    port map (
            O => \N__15488\,
            I => \N__15464\
        );

    \I__2930\ : SRMux
    port map (
            O => \N__15487\,
            I => \N__15464\
        );

    \I__2929\ : SRMux
    port map (
            O => \N__15486\,
            I => \N__15464\
        );

    \I__2928\ : Glb2LocalMux
    port map (
            O => \N__15483\,
            I => \N__15464\
        );

    \I__2927\ : GlobalMux
    port map (
            O => \N__15464\,
            I => \N__15461\
        );

    \I__2926\ : gio2CtrlBuf
    port map (
            O => \N__15461\,
            I => \this_vga_signals.N_684_g\
        );

    \I__2925\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15455\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__15455\,
            I => \this_vga_signals.N_272_0\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__15452\,
            I => \N__15443\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__15451\,
            I => \N__15437\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__15450\,
            I => \N__15434\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__15449\,
            I => \N__15419\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__15448\,
            I => \N__15416\
        );

    \I__2918\ : CascadeMux
    port map (
            O => \N__15447\,
            I => \N__15411\
        );

    \I__2917\ : InMux
    port map (
            O => \N__15446\,
            I => \N__15408\
        );

    \I__2916\ : InMux
    port map (
            O => \N__15443\,
            I => \N__15403\
        );

    \I__2915\ : InMux
    port map (
            O => \N__15442\,
            I => \N__15403\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__15441\,
            I => \N__15399\
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__15440\,
            I => \N__15394\
        );

    \I__2912\ : InMux
    port map (
            O => \N__15437\,
            I => \N__15389\
        );

    \I__2911\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15389\
        );

    \I__2910\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15384\
        );

    \I__2909\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15384\
        );

    \I__2908\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15381\
        );

    \I__2907\ : InMux
    port map (
            O => \N__15430\,
            I => \N__15376\
        );

    \I__2906\ : InMux
    port map (
            O => \N__15429\,
            I => \N__15376\
        );

    \I__2905\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15373\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__15427\,
            I => \N__15370\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__15426\,
            I => \N__15366\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__15425\,
            I => \N__15363\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__15424\,
            I => \N__15359\
        );

    \I__2900\ : InMux
    port map (
            O => \N__15423\,
            I => \N__15355\
        );

    \I__2899\ : InMux
    port map (
            O => \N__15422\,
            I => \N__15352\
        );

    \I__2898\ : InMux
    port map (
            O => \N__15419\,
            I => \N__15349\
        );

    \I__2897\ : InMux
    port map (
            O => \N__15416\,
            I => \N__15340\
        );

    \I__2896\ : InMux
    port map (
            O => \N__15415\,
            I => \N__15340\
        );

    \I__2895\ : InMux
    port map (
            O => \N__15414\,
            I => \N__15340\
        );

    \I__2894\ : InMux
    port map (
            O => \N__15411\,
            I => \N__15340\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__15408\,
            I => \N__15334\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__15403\,
            I => \N__15334\
        );

    \I__2891\ : InMux
    port map (
            O => \N__15402\,
            I => \N__15329\
        );

    \I__2890\ : InMux
    port map (
            O => \N__15399\,
            I => \N__15329\
        );

    \I__2889\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15326\
        );

    \I__2888\ : InMux
    port map (
            O => \N__15397\,
            I => \N__15323\
        );

    \I__2887\ : InMux
    port map (
            O => \N__15394\,
            I => \N__15320\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__15389\,
            I => \N__15315\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__15384\,
            I => \N__15315\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__15381\,
            I => \N__15308\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__15376\,
            I => \N__15308\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__15373\,
            I => \N__15308\
        );

    \I__2881\ : InMux
    port map (
            O => \N__15370\,
            I => \N__15301\
        );

    \I__2880\ : InMux
    port map (
            O => \N__15369\,
            I => \N__15301\
        );

    \I__2879\ : InMux
    port map (
            O => \N__15366\,
            I => \N__15301\
        );

    \I__2878\ : InMux
    port map (
            O => \N__15363\,
            I => \N__15296\
        );

    \I__2877\ : InMux
    port map (
            O => \N__15362\,
            I => \N__15296\
        );

    \I__2876\ : InMux
    port map (
            O => \N__15359\,
            I => \N__15293\
        );

    \I__2875\ : InMux
    port map (
            O => \N__15358\,
            I => \N__15290\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__15355\,
            I => \N__15285\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__15352\,
            I => \N__15285\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__15349\,
            I => \N__15280\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__15340\,
            I => \N__15280\
        );

    \I__2870\ : InMux
    port map (
            O => \N__15339\,
            I => \N__15277\
        );

    \I__2869\ : Span4Mux_h
    port map (
            O => \N__15334\,
            I => \N__15272\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__15329\,
            I => \N__15272\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__15326\,
            I => \N__15265\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__15323\,
            I => \N__15265\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__15320\,
            I => \N__15265\
        );

    \I__2864\ : Span4Mux_v
    port map (
            O => \N__15315\,
            I => \N__15261\
        );

    \I__2863\ : Span4Mux_h
    port map (
            O => \N__15308\,
            I => \N__15256\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__15301\,
            I => \N__15256\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__15296\,
            I => \N__15251\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__15293\,
            I => \N__15251\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__15290\,
            I => \N__15244\
        );

    \I__2858\ : Span4Mux_v
    port map (
            O => \N__15285\,
            I => \N__15244\
        );

    \I__2857\ : Span4Mux_v
    port map (
            O => \N__15280\,
            I => \N__15244\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__15277\,
            I => \N__15237\
        );

    \I__2855\ : Span4Mux_v
    port map (
            O => \N__15272\,
            I => \N__15237\
        );

    \I__2854\ : Span4Mux_h
    port map (
            O => \N__15265\,
            I => \N__15237\
        );

    \I__2853\ : InMux
    port map (
            O => \N__15264\,
            I => \N__15233\
        );

    \I__2852\ : Span4Mux_h
    port map (
            O => \N__15261\,
            I => \N__15228\
        );

    \I__2851\ : Span4Mux_v
    port map (
            O => \N__15256\,
            I => \N__15228\
        );

    \I__2850\ : Span4Mux_h
    port map (
            O => \N__15251\,
            I => \N__15225\
        );

    \I__2849\ : Span4Mux_h
    port map (
            O => \N__15244\,
            I => \N__15222\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__15237\,
            I => \N__15219\
        );

    \I__2847\ : InMux
    port map (
            O => \N__15236\,
            I => \N__15216\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__15233\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__2845\ : Odrv4
    port map (
            O => \N__15228\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__15225\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__2843\ : Odrv4
    port map (
            O => \N__15222\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__15219\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__15216\,
            I => \this_vga_signals_M_vcounter_q_4\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__15203\,
            I => \N__15198\
        );

    \I__2839\ : InMux
    port map (
            O => \N__15202\,
            I => \N__15195\
        );

    \I__2838\ : InMux
    port map (
            O => \N__15201\,
            I => \N__15192\
        );

    \I__2837\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15188\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__15195\,
            I => \N__15185\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__15192\,
            I => \N__15182\
        );

    \I__2834\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15179\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__15188\,
            I => \N__15176\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__15185\,
            I => \N__15173\
        );

    \I__2831\ : Span4Mux_h
    port map (
            O => \N__15182\,
            I => \N__15170\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__15179\,
            I => \N__15167\
        );

    \I__2829\ : Span4Mux_h
    port map (
            O => \N__15176\,
            I => \N__15164\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__15173\,
            I => \N_475\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__15170\,
            I => \N_475\
        );

    \I__2826\ : Odrv4
    port map (
            O => \N__15167\,
            I => \N_475\
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__15164\,
            I => \N_475\
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__15155\,
            I => \N__15147\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__15154\,
            I => \N__15144\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__15153\,
            I => \N__15138\
        );

    \I__2821\ : InMux
    port map (
            O => \N__15152\,
            I => \N__15132\
        );

    \I__2820\ : InMux
    port map (
            O => \N__15151\,
            I => \N__15129\
        );

    \I__2819\ : InMux
    port map (
            O => \N__15150\,
            I => \N__15122\
        );

    \I__2818\ : InMux
    port map (
            O => \N__15147\,
            I => \N__15119\
        );

    \I__2817\ : InMux
    port map (
            O => \N__15144\,
            I => \N__15110\
        );

    \I__2816\ : InMux
    port map (
            O => \N__15143\,
            I => \N__15110\
        );

    \I__2815\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15110\
        );

    \I__2814\ : InMux
    port map (
            O => \N__15141\,
            I => \N__15110\
        );

    \I__2813\ : InMux
    port map (
            O => \N__15138\,
            I => \N__15107\
        );

    \I__2812\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15101\
        );

    \I__2811\ : InMux
    port map (
            O => \N__15136\,
            I => \N__15098\
        );

    \I__2810\ : InMux
    port map (
            O => \N__15135\,
            I => \N__15095\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__15132\,
            I => \N__15087\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__15129\,
            I => \N__15087\
        );

    \I__2807\ : InMux
    port map (
            O => \N__15128\,
            I => \N__15084\
        );

    \I__2806\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15080\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__15126\,
            I => \N__15077\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__15125\,
            I => \N__15074\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__15122\,
            I => \N__15071\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__15119\,
            I => \N__15068\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__15110\,
            I => \N__15065\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__15107\,
            I => \N__15060\
        );

    \I__2799\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15053\
        );

    \I__2798\ : InMux
    port map (
            O => \N__15105\,
            I => \N__15053\
        );

    \I__2797\ : InMux
    port map (
            O => \N__15104\,
            I => \N__15053\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__15101\,
            I => \N__15050\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__15098\,
            I => \N__15045\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__15095\,
            I => \N__15045\
        );

    \I__2793\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15041\
        );

    \I__2792\ : InMux
    port map (
            O => \N__15093\,
            I => \N__15038\
        );

    \I__2791\ : InMux
    port map (
            O => \N__15092\,
            I => \N__15035\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__15087\,
            I => \N__15030\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__15084\,
            I => \N__15030\
        );

    \I__2788\ : InMux
    port map (
            O => \N__15083\,
            I => \N__15026\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__15080\,
            I => \N__15023\
        );

    \I__2786\ : InMux
    port map (
            O => \N__15077\,
            I => \N__15018\
        );

    \I__2785\ : InMux
    port map (
            O => \N__15074\,
            I => \N__15018\
        );

    \I__2784\ : Span4Mux_v
    port map (
            O => \N__15071\,
            I => \N__15011\
        );

    \I__2783\ : Span4Mux_v
    port map (
            O => \N__15068\,
            I => \N__15011\
        );

    \I__2782\ : Span4Mux_v
    port map (
            O => \N__15065\,
            I => \N__15011\
        );

    \I__2781\ : InMux
    port map (
            O => \N__15064\,
            I => \N__15006\
        );

    \I__2780\ : InMux
    port map (
            O => \N__15063\,
            I => \N__15006\
        );

    \I__2779\ : Span4Mux_h
    port map (
            O => \N__15060\,
            I => \N__14997\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__15053\,
            I => \N__14997\
        );

    \I__2777\ : Span4Mux_v
    port map (
            O => \N__15050\,
            I => \N__14997\
        );

    \I__2776\ : Span4Mux_h
    port map (
            O => \N__15045\,
            I => \N__14997\
        );

    \I__2775\ : InMux
    port map (
            O => \N__15044\,
            I => \N__14994\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__15041\,
            I => \N__14989\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__15038\,
            I => \N__14989\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__15035\,
            I => \N__14986\
        );

    \I__2771\ : Span4Mux_v
    port map (
            O => \N__15030\,
            I => \N__14983\
        );

    \I__2770\ : InMux
    port map (
            O => \N__15029\,
            I => \N__14980\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__15026\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__2768\ : Odrv4
    port map (
            O => \N__15023\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__15018\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__2766\ : Odrv4
    port map (
            O => \N__15011\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__15006\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__14997\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__14994\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__2762\ : Odrv12
    port map (
            O => \N__14989\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__2761\ : Odrv12
    port map (
            O => \N__14986\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__2760\ : Odrv4
    port map (
            O => \N__14983\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__14980\,
            I => \this_vga_signals_M_vcounter_q_5\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14957\,
            I => \N__14954\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__14954\,
            I => \N__14951\
        );

    \I__2756\ : Span4Mux_v
    port map (
            O => \N__14951\,
            I => \N__14948\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__14948\,
            I => \this_vga_signals.N_404_0\
        );

    \I__2754\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14941\
        );

    \I__2753\ : InMux
    port map (
            O => \N__14944\,
            I => \N__14938\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__14941\,
            I => \N_204_0\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__14938\,
            I => \N_204_0\
        );

    \I__2750\ : InMux
    port map (
            O => \N__14933\,
            I => \this_vga_signals.un1_M_hcounter_d_1_cry_1\
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__14930\,
            I => \this_vga_signals.mult1_un54_sum_axb1_0_cascade_\
        );

    \I__2748\ : InMux
    port map (
            O => \N__14927\,
            I => \N__14924\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__14924\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_x1\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__14921\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_\
        );

    \I__2745\ : InMux
    port map (
            O => \N__14918\,
            I => \N__14915\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__14915\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_1\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__14912\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_cascade_\
        );

    \I__2742\ : InMux
    port map (
            O => \N__14909\,
            I => \N__14904\
        );

    \I__2741\ : InMux
    port map (
            O => \N__14908\,
            I => \N__14899\
        );

    \I__2740\ : InMux
    port map (
            O => \N__14907\,
            I => \N__14899\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__14904\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_1\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__14899\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_1\
        );

    \I__2737\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14891\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__14891\,
            I => \N__14887\
        );

    \I__2735\ : InMux
    port map (
            O => \N__14890\,
            I => \N__14884\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__14887\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__14884\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\
        );

    \I__2732\ : CascadeMux
    port map (
            O => \N__14879\,
            I => \N__14876\
        );

    \I__2731\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14873\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__14873\,
            I => \N__14870\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__14870\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\
        );

    \I__2728\ : InMux
    port map (
            O => \N__14867\,
            I => \N__14864\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__14864\,
            I => \N__14859\
        );

    \I__2726\ : InMux
    port map (
            O => \N__14863\,
            I => \N__14854\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14862\,
            I => \N__14854\
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__14859\,
            I => \this_vga_signals.N_336_0\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__14854\,
            I => \this_vga_signals.N_336_0\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__14849\,
            I => \this_vga_signals.N_336_0_cascade_\
        );

    \I__2721\ : InMux
    port map (
            O => \N__14846\,
            I => \N__14840\
        );

    \I__2720\ : InMux
    port map (
            O => \N__14845\,
            I => \N__14833\
        );

    \I__2719\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14833\
        );

    \I__2718\ : InMux
    port map (
            O => \N__14843\,
            I => \N__14833\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__14840\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_6\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__14833\,
            I => \this_vga_signals.M_hcounter_q_fastZ0Z_6\
        );

    \I__2715\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14825\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__14825\,
            I => \this_vga_signals.N_287\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__14822\,
            I => \this_vga_signals.N_287_cascade_\
        );

    \I__2712\ : InMux
    port map (
            O => \N__14819\,
            I => \N__14816\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__14816\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2_1_0\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__14813\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_\
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__14810\,
            I => \this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3_cascade_\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__14807\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_1_cascade_\
        );

    \I__2707\ : InMux
    port map (
            O => \N__14804\,
            I => \N__14794\
        );

    \I__2706\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14794\
        );

    \I__2705\ : InMux
    port map (
            O => \N__14802\,
            I => \N__14794\
        );

    \I__2704\ : InMux
    port map (
            O => \N__14801\,
            I => \N__14791\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__14794\,
            I => \this_vga_signals.SUM_7_i_1_0\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__14791\,
            I => \this_vga_signals.SUM_7_i_1_0\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__14786\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\
        );

    \I__2700\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14780\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__14780\,
            I => \G_504\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__14777\,
            I => \N__14774\
        );

    \I__2697\ : InMux
    port map (
            O => \N__14774\,
            I => \N__14771\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__14771\,
            I => \N__14768\
        );

    \I__2695\ : Span4Mux_v
    port map (
            O => \N__14768\,
            I => \N__14765\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__14765\,
            I => \this_vga_signals.mult1_un68_sum_cry_1_s\
        );

    \I__2693\ : InMux
    port map (
            O => \N__14762\,
            I => \N__14759\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__14759\,
            I => \G_503\
        );

    \I__2691\ : InMux
    port map (
            O => \N__14756\,
            I => \N__14753\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__14753\,
            I => \N__14750\
        );

    \I__2689\ : Odrv4
    port map (
            O => \N__14750\,
            I => \this_vga_signals.mult1_un75_sum_axb_3\
        );

    \I__2688\ : InMux
    port map (
            O => \N__14747\,
            I => \this_vga_signals.mult1_un75_sum_cry_2\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__14744\,
            I => \this_ppu.M_m12_0_o2_381Z0Z_4_cascade_\
        );

    \I__2686\ : InMux
    port map (
            O => \N__14741\,
            I => \N__14737\
        );

    \I__2685\ : InMux
    port map (
            O => \N__14740\,
            I => \N__14734\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__14737\,
            I => \N__14731\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__14734\,
            I => \N_275\
        );

    \I__2682\ : Odrv4
    port map (
            O => \N__14731\,
            I => \N_275\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__14726\,
            I => \this_ppu.M_m12_0_o2_381_5_cascade_\
        );

    \I__2680\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14720\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__14720\,
            I => \N__14717\
        );

    \I__2678\ : Span4Mux_h
    port map (
            O => \N__14717\,
            I => \N__14712\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14716\,
            I => \N__14709\
        );

    \I__2676\ : InMux
    port map (
            O => \N__14715\,
            I => \N__14706\
        );

    \I__2675\ : Odrv4
    port map (
            O => \N__14712\,
            I => \N_190_0\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__14709\,
            I => \N_190_0\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__14706\,
            I => \N_190_0\
        );

    \I__2672\ : InMux
    port map (
            O => \N__14699\,
            I => \N__14696\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__14696\,
            I => \N__14693\
        );

    \I__2670\ : Span4Mux_h
    port map (
            O => \N__14693\,
            I => \N__14690\
        );

    \I__2669\ : Odrv4
    port map (
            O => \N__14690\,
            I => \this_ppu.M_m12_0_o2_381_8\
        );

    \I__2668\ : InMux
    port map (
            O => \N__14687\,
            I => \N__14682\
        );

    \I__2667\ : InMux
    port map (
            O => \N__14686\,
            I => \N__14677\
        );

    \I__2666\ : InMux
    port map (
            O => \N__14685\,
            I => \N__14677\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__14682\,
            I => \M_this_delay_clk_out_0\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__14677\,
            I => \M_this_delay_clk_out_0\
        );

    \I__2663\ : InMux
    port map (
            O => \N__14672\,
            I => \N__14665\
        );

    \I__2662\ : InMux
    port map (
            O => \N__14671\,
            I => \N__14665\
        );

    \I__2661\ : InMux
    port map (
            O => \N__14670\,
            I => \N__14662\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__14665\,
            I => \N__14657\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__14662\,
            I => \N__14657\
        );

    \I__2658\ : Span4Mux_v
    port map (
            O => \N__14657\,
            I => \N__14654\
        );

    \I__2657\ : Span4Mux_h
    port map (
            O => \N__14654\,
            I => \N__14651\
        );

    \I__2656\ : Span4Mux_h
    port map (
            O => \N__14651\,
            I => \N__14648\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__14648\,
            I => port_enb_c
        );

    \I__2654\ : InMux
    port map (
            O => \N__14645\,
            I => \N__14642\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__14642\,
            I => \N__14638\
        );

    \I__2652\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14635\
        );

    \I__2651\ : Odrv4
    port map (
            O => \N__14638\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__14635\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__2649\ : InMux
    port map (
            O => \N__14630\,
            I => \N__14627\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__14627\,
            I => \this_vga_signals.mult1_un61_sum_i_0\
        );

    \I__2647\ : InMux
    port map (
            O => \N__14624\,
            I => \N__14620\
        );

    \I__2646\ : InMux
    port map (
            O => \N__14623\,
            I => \N__14617\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__14620\,
            I => \N__14614\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__14617\,
            I => \N__14611\
        );

    \I__2643\ : Span4Mux_h
    port map (
            O => \N__14614\,
            I => \N__14608\
        );

    \I__2642\ : Span4Mux_h
    port map (
            O => \N__14611\,
            I => \N__14605\
        );

    \I__2641\ : Span4Mux_v
    port map (
            O => \N__14608\,
            I => \N__14602\
        );

    \I__2640\ : Odrv4
    port map (
            O => \N__14605\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1_0\
        );

    \I__2639\ : Odrv4
    port map (
            O => \N__14602\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1_0\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__14597\,
            I => \N__14594\
        );

    \I__2637\ : InMux
    port map (
            O => \N__14594\,
            I => \N__14591\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__14591\,
            I => \N__14588\
        );

    \I__2635\ : Span12Mux_h
    port map (
            O => \N__14588\,
            I => \N__14585\
        );

    \I__2634\ : Odrv12
    port map (
            O => \N__14585\,
            I => \N_90_0\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__14582\,
            I => \N__14569\
        );

    \I__2632\ : CascadeMux
    port map (
            O => \N__14581\,
            I => \N__14566\
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__14580\,
            I => \N__14558\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__14579\,
            I => \N__14552\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__14578\,
            I => \N__14548\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__14577\,
            I => \N__14545\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__14576\,
            I => \N__14542\
        );

    \I__2626\ : InMux
    port map (
            O => \N__14575\,
            I => \N__14535\
        );

    \I__2625\ : InMux
    port map (
            O => \N__14574\,
            I => \N__14535\
        );

    \I__2624\ : InMux
    port map (
            O => \N__14573\,
            I => \N__14532\
        );

    \I__2623\ : InMux
    port map (
            O => \N__14572\,
            I => \N__14526\
        );

    \I__2622\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14526\
        );

    \I__2621\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14519\
        );

    \I__2620\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14519\
        );

    \I__2619\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14519\
        );

    \I__2618\ : InMux
    port map (
            O => \N__14563\,
            I => \N__14514\
        );

    \I__2617\ : InMux
    port map (
            O => \N__14562\,
            I => \N__14514\
        );

    \I__2616\ : CascadeMux
    port map (
            O => \N__14561\,
            I => \N__14509\
        );

    \I__2615\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14506\
        );

    \I__2614\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14499\
        );

    \I__2613\ : InMux
    port map (
            O => \N__14556\,
            I => \N__14499\
        );

    \I__2612\ : InMux
    port map (
            O => \N__14555\,
            I => \N__14499\
        );

    \I__2611\ : InMux
    port map (
            O => \N__14552\,
            I => \N__14495\
        );

    \I__2610\ : InMux
    port map (
            O => \N__14551\,
            I => \N__14488\
        );

    \I__2609\ : InMux
    port map (
            O => \N__14548\,
            I => \N__14488\
        );

    \I__2608\ : InMux
    port map (
            O => \N__14545\,
            I => \N__14488\
        );

    \I__2607\ : InMux
    port map (
            O => \N__14542\,
            I => \N__14483\
        );

    \I__2606\ : InMux
    port map (
            O => \N__14541\,
            I => \N__14483\
        );

    \I__2605\ : InMux
    port map (
            O => \N__14540\,
            I => \N__14480\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__14535\,
            I => \N__14475\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__14532\,
            I => \N__14475\
        );

    \I__2602\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14472\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__14526\,
            I => \N__14465\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__14519\,
            I => \N__14465\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__14514\,
            I => \N__14462\
        );

    \I__2598\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14459\
        );

    \I__2597\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14454\
        );

    \I__2596\ : InMux
    port map (
            O => \N__14509\,
            I => \N__14454\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__14506\,
            I => \N__14449\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__14499\,
            I => \N__14449\
        );

    \I__2593\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14446\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__14495\,
            I => \N__14443\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__14488\,
            I => \N__14434\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__14483\,
            I => \N__14434\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__14480\,
            I => \N__14434\
        );

    \I__2588\ : Span4Mux_h
    port map (
            O => \N__14475\,
            I => \N__14434\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__14472\,
            I => \N__14431\
        );

    \I__2586\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14428\
        );

    \I__2585\ : InMux
    port map (
            O => \N__14470\,
            I => \N__14425\
        );

    \I__2584\ : Span4Mux_v
    port map (
            O => \N__14465\,
            I => \N__14420\
        );

    \I__2583\ : Span4Mux_h
    port map (
            O => \N__14462\,
            I => \N__14420\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__14459\,
            I => \N__14415\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__14454\,
            I => \N__14415\
        );

    \I__2580\ : Span4Mux_v
    port map (
            O => \N__14449\,
            I => \N__14410\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__14446\,
            I => \N__14410\
        );

    \I__2578\ : Span4Mux_v
    port map (
            O => \N__14443\,
            I => \N__14403\
        );

    \I__2577\ : Span4Mux_v
    port map (
            O => \N__14434\,
            I => \N__14403\
        );

    \I__2576\ : Span4Mux_v
    port map (
            O => \N__14431\,
            I => \N__14403\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__14428\,
            I => \N__14400\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__14425\,
            I => \this_vga_signals_M_vcounter_q_2\
        );

    \I__2573\ : Odrv4
    port map (
            O => \N__14420\,
            I => \this_vga_signals_M_vcounter_q_2\
        );

    \I__2572\ : Odrv12
    port map (
            O => \N__14415\,
            I => \this_vga_signals_M_vcounter_q_2\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__14410\,
            I => \this_vga_signals_M_vcounter_q_2\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__14403\,
            I => \this_vga_signals_M_vcounter_q_2\
        );

    \I__2569\ : Odrv4
    port map (
            O => \N__14400\,
            I => \this_vga_signals_M_vcounter_q_2\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__14387\,
            I => \N__14380\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__14386\,
            I => \N__14362\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__14385\,
            I => \N__14359\
        );

    \I__2565\ : InMux
    port map (
            O => \N__14384\,
            I => \N__14356\
        );

    \I__2564\ : InMux
    port map (
            O => \N__14383\,
            I => \N__14351\
        );

    \I__2563\ : InMux
    port map (
            O => \N__14380\,
            I => \N__14351\
        );

    \I__2562\ : InMux
    port map (
            O => \N__14379\,
            I => \N__14348\
        );

    \I__2561\ : InMux
    port map (
            O => \N__14378\,
            I => \N__14339\
        );

    \I__2560\ : InMux
    port map (
            O => \N__14377\,
            I => \N__14336\
        );

    \I__2559\ : InMux
    port map (
            O => \N__14376\,
            I => \N__14330\
        );

    \I__2558\ : InMux
    port map (
            O => \N__14375\,
            I => \N__14327\
        );

    \I__2557\ : InMux
    port map (
            O => \N__14374\,
            I => \N__14324\
        );

    \I__2556\ : InMux
    port map (
            O => \N__14373\,
            I => \N__14321\
        );

    \I__2555\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14312\
        );

    \I__2554\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14312\
        );

    \I__2553\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14312\
        );

    \I__2552\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14312\
        );

    \I__2551\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14307\
        );

    \I__2550\ : InMux
    port map (
            O => \N__14367\,
            I => \N__14307\
        );

    \I__2549\ : InMux
    port map (
            O => \N__14366\,
            I => \N__14296\
        );

    \I__2548\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14296\
        );

    \I__2547\ : InMux
    port map (
            O => \N__14362\,
            I => \N__14291\
        );

    \I__2546\ : InMux
    port map (
            O => \N__14359\,
            I => \N__14291\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__14356\,
            I => \N__14284\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__14351\,
            I => \N__14284\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__14348\,
            I => \N__14284\
        );

    \I__2542\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14281\
        );

    \I__2541\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14276\
        );

    \I__2540\ : InMux
    port map (
            O => \N__14345\,
            I => \N__14276\
        );

    \I__2539\ : InMux
    port map (
            O => \N__14344\,
            I => \N__14271\
        );

    \I__2538\ : InMux
    port map (
            O => \N__14343\,
            I => \N__14271\
        );

    \I__2537\ : InMux
    port map (
            O => \N__14342\,
            I => \N__14267\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__14339\,
            I => \N__14262\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__14336\,
            I => \N__14262\
        );

    \I__2534\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14259\
        );

    \I__2533\ : InMux
    port map (
            O => \N__14334\,
            I => \N__14256\
        );

    \I__2532\ : InMux
    port map (
            O => \N__14333\,
            I => \N__14251\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__14330\,
            I => \N__14242\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__14327\,
            I => \N__14242\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__14324\,
            I => \N__14242\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__14321\,
            I => \N__14242\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__14312\,
            I => \N__14237\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__14307\,
            I => \N__14237\
        );

    \I__2525\ : InMux
    port map (
            O => \N__14306\,
            I => \N__14234\
        );

    \I__2524\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14227\
        );

    \I__2523\ : InMux
    port map (
            O => \N__14304\,
            I => \N__14227\
        );

    \I__2522\ : InMux
    port map (
            O => \N__14303\,
            I => \N__14227\
        );

    \I__2521\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14224\
        );

    \I__2520\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14221\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__14296\,
            I => \N__14214\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__14291\,
            I => \N__14214\
        );

    \I__2517\ : Span4Mux_h
    port map (
            O => \N__14284\,
            I => \N__14214\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__14281\,
            I => \N__14207\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__14276\,
            I => \N__14207\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__14271\,
            I => \N__14207\
        );

    \I__2513\ : InMux
    port map (
            O => \N__14270\,
            I => \N__14204\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__14267\,
            I => \N__14197\
        );

    \I__2511\ : Span4Mux_v
    port map (
            O => \N__14262\,
            I => \N__14197\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__14259\,
            I => \N__14197\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__14256\,
            I => \N__14194\
        );

    \I__2508\ : InMux
    port map (
            O => \N__14255\,
            I => \N__14191\
        );

    \I__2507\ : InMux
    port map (
            O => \N__14254\,
            I => \N__14188\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__14251\,
            I => \N__14185\
        );

    \I__2505\ : Span4Mux_v
    port map (
            O => \N__14242\,
            I => \N__14180\
        );

    \I__2504\ : Span4Mux_h
    port map (
            O => \N__14237\,
            I => \N__14180\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__14234\,
            I => \N__14173\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__14227\,
            I => \N__14173\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__14224\,
            I => \N__14173\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__14221\,
            I => \N__14164\
        );

    \I__2499\ : Span4Mux_v
    port map (
            O => \N__14214\,
            I => \N__14164\
        );

    \I__2498\ : Span4Mux_v
    port map (
            O => \N__14207\,
            I => \N__14164\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__14204\,
            I => \N__14164\
        );

    \I__2496\ : Span4Mux_v
    port map (
            O => \N__14197\,
            I => \N__14157\
        );

    \I__2495\ : Span4Mux_v
    port map (
            O => \N__14194\,
            I => \N__14157\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__14191\,
            I => \N__14157\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__14188\,
            I => \this_vga_signals_M_vcounter_q_3\
        );

    \I__2492\ : Odrv12
    port map (
            O => \N__14185\,
            I => \this_vga_signals_M_vcounter_q_3\
        );

    \I__2491\ : Odrv4
    port map (
            O => \N__14180\,
            I => \this_vga_signals_M_vcounter_q_3\
        );

    \I__2490\ : Odrv4
    port map (
            O => \N__14173\,
            I => \this_vga_signals_M_vcounter_q_3\
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__14164\,
            I => \this_vga_signals_M_vcounter_q_3\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__14157\,
            I => \this_vga_signals_M_vcounter_q_3\
        );

    \I__2487\ : InMux
    port map (
            O => \N__14144\,
            I => \N__14141\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__14141\,
            I => \N__14138\
        );

    \I__2485\ : Span4Mux_h
    port map (
            O => \N__14138\,
            I => \N__14135\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__14135\,
            I => \N_184_0\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__14132\,
            I => \N__14123\
        );

    \I__2482\ : InMux
    port map (
            O => \N__14131\,
            I => \N__14119\
        );

    \I__2481\ : InMux
    port map (
            O => \N__14130\,
            I => \N__14115\
        );

    \I__2480\ : CascadeMux
    port map (
            O => \N__14129\,
            I => \N__14110\
        );

    \I__2479\ : InMux
    port map (
            O => \N__14128\,
            I => \N__14104\
        );

    \I__2478\ : InMux
    port map (
            O => \N__14127\,
            I => \N__14101\
        );

    \I__2477\ : InMux
    port map (
            O => \N__14126\,
            I => \N__14098\
        );

    \I__2476\ : InMux
    port map (
            O => \N__14123\,
            I => \N__14095\
        );

    \I__2475\ : InMux
    port map (
            O => \N__14122\,
            I => \N__14092\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__14119\,
            I => \N__14088\
        );

    \I__2473\ : InMux
    port map (
            O => \N__14118\,
            I => \N__14085\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__14115\,
            I => \N__14082\
        );

    \I__2471\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14075\
        );

    \I__2470\ : InMux
    port map (
            O => \N__14113\,
            I => \N__14075\
        );

    \I__2469\ : InMux
    port map (
            O => \N__14110\,
            I => \N__14075\
        );

    \I__2468\ : InMux
    port map (
            O => \N__14109\,
            I => \N__14068\
        );

    \I__2467\ : InMux
    port map (
            O => \N__14108\,
            I => \N__14068\
        );

    \I__2466\ : InMux
    port map (
            O => \N__14107\,
            I => \N__14068\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__14104\,
            I => \N__14063\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__14101\,
            I => \N__14060\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__14098\,
            I => \N__14057\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__14095\,
            I => \N__14054\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__14092\,
            I => \N__14051\
        );

    \I__2460\ : InMux
    port map (
            O => \N__14091\,
            I => \N__14048\
        );

    \I__2459\ : Span4Mux_h
    port map (
            O => \N__14088\,
            I => \N__14045\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__14085\,
            I => \N__14042\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__14082\,
            I => \N__14035\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__14075\,
            I => \N__14035\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__14068\,
            I => \N__14035\
        );

    \I__2454\ : InMux
    port map (
            O => \N__14067\,
            I => \N__14032\
        );

    \I__2453\ : InMux
    port map (
            O => \N__14066\,
            I => \N__14029\
        );

    \I__2452\ : Span4Mux_v
    port map (
            O => \N__14063\,
            I => \N__14022\
        );

    \I__2451\ : Span4Mux_v
    port map (
            O => \N__14060\,
            I => \N__14022\
        );

    \I__2450\ : Span4Mux_v
    port map (
            O => \N__14057\,
            I => \N__14022\
        );

    \I__2449\ : Span4Mux_v
    port map (
            O => \N__14054\,
            I => \N__14017\
        );

    \I__2448\ : Span4Mux_v
    port map (
            O => \N__14051\,
            I => \N__14017\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__14048\,
            I => \N__14014\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__14045\,
            I => \N__14007\
        );

    \I__2445\ : Span4Mux_v
    port map (
            O => \N__14042\,
            I => \N__14007\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__14035\,
            I => \N__14007\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__14032\,
            I => \N__14004\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__14029\,
            I => \this_vga_signals_M_vcounter_q_1\
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__14022\,
            I => \this_vga_signals_M_vcounter_q_1\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__14017\,
            I => \this_vga_signals_M_vcounter_q_1\
        );

    \I__2439\ : Odrv12
    port map (
            O => \N__14014\,
            I => \this_vga_signals_M_vcounter_q_1\
        );

    \I__2438\ : Odrv4
    port map (
            O => \N__14007\,
            I => \this_vga_signals_M_vcounter_q_1\
        );

    \I__2437\ : Odrv12
    port map (
            O => \N__14004\,
            I => \this_vga_signals_M_vcounter_q_1\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__13991\,
            I => \N_184_0_cascade_\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__13988\,
            I => \N__13982\
        );

    \I__2434\ : InMux
    port map (
            O => \N__13987\,
            I => \N__13978\
        );

    \I__2433\ : InMux
    port map (
            O => \N__13986\,
            I => \N__13974\
        );

    \I__2432\ : InMux
    port map (
            O => \N__13985\,
            I => \N__13967\
        );

    \I__2431\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13967\
        );

    \I__2430\ : InMux
    port map (
            O => \N__13981\,
            I => \N__13967\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__13978\,
            I => \N__13962\
        );

    \I__2428\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13959\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__13974\,
            I => \N__13954\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__13967\,
            I => \N__13954\
        );

    \I__2425\ : InMux
    port map (
            O => \N__13966\,
            I => \N__13951\
        );

    \I__2424\ : InMux
    port map (
            O => \N__13965\,
            I => \N__13948\
        );

    \I__2423\ : Sp12to4
    port map (
            O => \N__13962\,
            I => \N__13943\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__13959\,
            I => \N__13943\
        );

    \I__2421\ : Span4Mux_v
    port map (
            O => \N__13954\,
            I => \N__13938\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__13951\,
            I => \N__13938\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__13948\,
            I => \this_vga_signals_M_vcounter_q_0\
        );

    \I__2418\ : Odrv12
    port map (
            O => \N__13943\,
            I => \this_vga_signals_M_vcounter_q_0\
        );

    \I__2417\ : Odrv4
    port map (
            O => \N__13938\,
            I => \this_vga_signals_M_vcounter_q_0\
        );

    \I__2416\ : InMux
    port map (
            O => \N__13931\,
            I => \N__13920\
        );

    \I__2415\ : InMux
    port map (
            O => \N__13930\,
            I => \N__13913\
        );

    \I__2414\ : InMux
    port map (
            O => \N__13929\,
            I => \N__13913\
        );

    \I__2413\ : InMux
    port map (
            O => \N__13928\,
            I => \N__13913\
        );

    \I__2412\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13908\
        );

    \I__2411\ : InMux
    port map (
            O => \N__13926\,
            I => \N__13903\
        );

    \I__2410\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13903\
        );

    \I__2409\ : InMux
    port map (
            O => \N__13924\,
            I => \N__13900\
        );

    \I__2408\ : InMux
    port map (
            O => \N__13923\,
            I => \N__13897\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__13920\,
            I => \N__13892\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__13913\,
            I => \N__13892\
        );

    \I__2405\ : InMux
    port map (
            O => \N__13912\,
            I => \N__13887\
        );

    \I__2404\ : InMux
    port map (
            O => \N__13911\,
            I => \N__13887\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__13908\,
            I => \N__13881\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__13903\,
            I => \N__13874\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__13900\,
            I => \N__13874\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__13897\,
            I => \N__13874\
        );

    \I__2399\ : Span4Mux_v
    port map (
            O => \N__13892\,
            I => \N__13869\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__13887\,
            I => \N__13869\
        );

    \I__2397\ : InMux
    port map (
            O => \N__13886\,
            I => \N__13866\
        );

    \I__2396\ : InMux
    port map (
            O => \N__13885\,
            I => \N__13863\
        );

    \I__2395\ : InMux
    port map (
            O => \N__13884\,
            I => \N__13860\
        );

    \I__2394\ : Odrv4
    port map (
            O => \N__13881\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__13874\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__13869\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__13866\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__13863\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__13860\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2388\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13844\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__13844\,
            I => \this_vga_signals.if_N_8_0\
        );

    \I__2386\ : InMux
    port map (
            O => \N__13841\,
            I => \N__13838\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__13838\,
            I => \N__13835\
        );

    \I__2384\ : Span4Mux_v
    port map (
            O => \N__13835\,
            I => \N__13832\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__13832\,
            I => \this_vga_signals.mult1_un54_sum_i_0\
        );

    \I__2382\ : IoInMux
    port map (
            O => \N__13829\,
            I => \N__13826\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__13826\,
            I => \N__13823\
        );

    \I__2380\ : IoSpan4Mux
    port map (
            O => \N__13823\,
            I => \N__13820\
        );

    \I__2379\ : IoSpan4Mux
    port map (
            O => \N__13820\,
            I => \N__13817\
        );

    \I__2378\ : Span4Mux_s2_v
    port map (
            O => \N__13817\,
            I => \N__13814\
        );

    \I__2377\ : Sp12to4
    port map (
            O => \N__13814\,
            I => \N__13811\
        );

    \I__2376\ : Span12Mux_v
    port map (
            O => \N__13811\,
            I => \N__13808\
        );

    \I__2375\ : Odrv12
    port map (
            O => \N__13808\,
            I => \N_31\
        );

    \I__2374\ : InMux
    port map (
            O => \N__13805\,
            I => \N__13794\
        );

    \I__2373\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13785\
        );

    \I__2372\ : InMux
    port map (
            O => \N__13803\,
            I => \N__13782\
        );

    \I__2371\ : InMux
    port map (
            O => \N__13802\,
            I => \N__13777\
        );

    \I__2370\ : InMux
    port map (
            O => \N__13801\,
            I => \N__13777\
        );

    \I__2369\ : InMux
    port map (
            O => \N__13800\,
            I => \N__13774\
        );

    \I__2368\ : InMux
    port map (
            O => \N__13799\,
            I => \N__13770\
        );

    \I__2367\ : InMux
    port map (
            O => \N__13798\,
            I => \N__13767\
        );

    \I__2366\ : InMux
    port map (
            O => \N__13797\,
            I => \N__13764\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__13794\,
            I => \N__13761\
        );

    \I__2364\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13758\
        );

    \I__2363\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13751\
        );

    \I__2362\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13751\
        );

    \I__2361\ : InMux
    port map (
            O => \N__13790\,
            I => \N__13751\
        );

    \I__2360\ : InMux
    port map (
            O => \N__13789\,
            I => \N__13746\
        );

    \I__2359\ : InMux
    port map (
            O => \N__13788\,
            I => \N__13746\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__13785\,
            I => \N__13743\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__13782\,
            I => \N__13736\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__13777\,
            I => \N__13736\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__13774\,
            I => \N__13736\
        );

    \I__2354\ : InMux
    port map (
            O => \N__13773\,
            I => \N__13733\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__13770\,
            I => \N__13728\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__13767\,
            I => \N__13728\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__13764\,
            I => \N__13723\
        );

    \I__2350\ : Span4Mux_v
    port map (
            O => \N__13761\,
            I => \N__13723\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__13758\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__13751\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__13746\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2346\ : Odrv4
    port map (
            O => \N__13743\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__13736\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__13733\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__13728\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__13723\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2341\ : InMux
    port map (
            O => \N__13706\,
            I => \N__13702\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__13705\,
            I => \N__13694\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__13702\,
            I => \N__13691\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__13701\,
            I => \N__13687\
        );

    \I__2337\ : InMux
    port map (
            O => \N__13700\,
            I => \N__13684\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13699\,
            I => \N__13678\
        );

    \I__2335\ : InMux
    port map (
            O => \N__13698\,
            I => \N__13678\
        );

    \I__2334\ : InMux
    port map (
            O => \N__13697\,
            I => \N__13669\
        );

    \I__2333\ : InMux
    port map (
            O => \N__13694\,
            I => \N__13669\
        );

    \I__2332\ : Span4Mux_v
    port map (
            O => \N__13691\,
            I => \N__13666\
        );

    \I__2331\ : InMux
    port map (
            O => \N__13690\,
            I => \N__13663\
        );

    \I__2330\ : InMux
    port map (
            O => \N__13687\,
            I => \N__13660\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__13684\,
            I => \N__13657\
        );

    \I__2328\ : InMux
    port map (
            O => \N__13683\,
            I => \N__13652\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__13678\,
            I => \N__13648\
        );

    \I__2326\ : InMux
    port map (
            O => \N__13677\,
            I => \N__13645\
        );

    \I__2325\ : InMux
    port map (
            O => \N__13676\,
            I => \N__13642\
        );

    \I__2324\ : InMux
    port map (
            O => \N__13675\,
            I => \N__13637\
        );

    \I__2323\ : InMux
    port map (
            O => \N__13674\,
            I => \N__13637\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__13669\,
            I => \N__13634\
        );

    \I__2321\ : Span4Mux_v
    port map (
            O => \N__13666\,
            I => \N__13629\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__13663\,
            I => \N__13629\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__13660\,
            I => \N__13626\
        );

    \I__2318\ : Span4Mux_h
    port map (
            O => \N__13657\,
            I => \N__13623\
        );

    \I__2317\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13618\
        );

    \I__2316\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13618\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__13652\,
            I => \N__13615\
        );

    \I__2314\ : InMux
    port map (
            O => \N__13651\,
            I => \N__13612\
        );

    \I__2313\ : Span4Mux_h
    port map (
            O => \N__13648\,
            I => \N__13601\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__13645\,
            I => \N__13601\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__13642\,
            I => \N__13601\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__13637\,
            I => \N__13601\
        );

    \I__2309\ : Span4Mux_h
    port map (
            O => \N__13634\,
            I => \N__13601\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__13629\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__2307\ : Odrv12
    port map (
            O => \N__13626\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__13623\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__13618\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__2304\ : Odrv4
    port map (
            O => \N__13615\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__13612\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__13601\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__13586\,
            I => \N__13579\
        );

    \I__2300\ : InMux
    port map (
            O => \N__13585\,
            I => \N__13575\
        );

    \I__2299\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13572\
        );

    \I__2298\ : InMux
    port map (
            O => \N__13583\,
            I => \N__13569\
        );

    \I__2297\ : InMux
    port map (
            O => \N__13582\,
            I => \N__13564\
        );

    \I__2296\ : InMux
    port map (
            O => \N__13579\,
            I => \N__13561\
        );

    \I__2295\ : InMux
    port map (
            O => \N__13578\,
            I => \N__13558\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__13575\,
            I => \N__13551\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__13572\,
            I => \N__13546\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__13569\,
            I => \N__13546\
        );

    \I__2291\ : InMux
    port map (
            O => \N__13568\,
            I => \N__13539\
        );

    \I__2290\ : InMux
    port map (
            O => \N__13567\,
            I => \N__13539\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__13564\,
            I => \N__13534\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__13561\,
            I => \N__13534\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__13558\,
            I => \N__13531\
        );

    \I__2286\ : InMux
    port map (
            O => \N__13557\,
            I => \N__13528\
        );

    \I__2285\ : InMux
    port map (
            O => \N__13556\,
            I => \N__13523\
        );

    \I__2284\ : InMux
    port map (
            O => \N__13555\,
            I => \N__13523\
        );

    \I__2283\ : InMux
    port map (
            O => \N__13554\,
            I => \N__13520\
        );

    \I__2282\ : Span4Mux_v
    port map (
            O => \N__13551\,
            I => \N__13515\
        );

    \I__2281\ : Span4Mux_v
    port map (
            O => \N__13546\,
            I => \N__13515\
        );

    \I__2280\ : InMux
    port map (
            O => \N__13545\,
            I => \N__13510\
        );

    \I__2279\ : InMux
    port map (
            O => \N__13544\,
            I => \N__13510\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__13539\,
            I => \N__13507\
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__13534\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__13531\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__13528\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__13523\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__13520\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__13515\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__13510\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2270\ : Odrv4
    port map (
            O => \N__13507\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__13490\,
            I => \this_vga_signals.N_177_0_cascade_\
        );

    \I__2268\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13482\
        );

    \I__2267\ : InMux
    port map (
            O => \N__13486\,
            I => \N__13478\
        );

    \I__2266\ : CascadeMux
    port map (
            O => \N__13485\,
            I => \N__13475\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__13482\,
            I => \N__13472\
        );

    \I__2264\ : InMux
    port map (
            O => \N__13481\,
            I => \N__13469\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__13478\,
            I => \N__13466\
        );

    \I__2262\ : InMux
    port map (
            O => \N__13475\,
            I => \N__13463\
        );

    \I__2261\ : Span4Mux_v
    port map (
            O => \N__13472\,
            I => \N__13458\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__13469\,
            I => \N__13458\
        );

    \I__2259\ : Span4Mux_v
    port map (
            O => \N__13466\,
            I => \N__13453\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__13463\,
            I => \N__13453\
        );

    \I__2257\ : Span4Mux_h
    port map (
            O => \N__13458\,
            I => \N__13450\
        );

    \I__2256\ : Span4Mux_v
    port map (
            O => \N__13453\,
            I => \N__13447\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__13450\,
            I => \N__13444\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__13447\,
            I => \this_vga_signals.CO0_i_0\
        );

    \I__2253\ : Odrv4
    port map (
            O => \N__13444\,
            I => \this_vga_signals.CO0_i_0\
        );

    \I__2252\ : InMux
    port map (
            O => \N__13439\,
            I => \N__13436\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__13436\,
            I => \this_vga_signals.N_269_0\
        );

    \I__2250\ : InMux
    port map (
            O => \N__13433\,
            I => \N__13430\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__13430\,
            I => \this_vga_signals.N_286\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__13427\,
            I => \this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1_cascade_\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__13424\,
            I => \N__13420\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__13423\,
            I => \N__13417\
        );

    \I__2245\ : InMux
    port map (
            O => \N__13420\,
            I => \N__13414\
        );

    \I__2244\ : InMux
    port map (
            O => \N__13417\,
            I => \N__13411\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__13414\,
            I => \N__13408\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__13411\,
            I => \N__13405\
        );

    \I__2241\ : Span4Mux_h
    port map (
            O => \N__13408\,
            I => \N__13402\
        );

    \I__2240\ : Span4Mux_h
    port map (
            O => \N__13405\,
            I => \N__13399\
        );

    \I__2239\ : Odrv4
    port map (
            O => \N__13402\,
            I => \this_vga_signals.N_188_0_0_0\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__13399\,
            I => \this_vga_signals.N_188_0_0_0\
        );

    \I__2237\ : InMux
    port map (
            O => \N__13394\,
            I => \N__13391\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__13391\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_1_0_3\
        );

    \I__2235\ : CascadeMux
    port map (
            O => \N__13388\,
            I => \this_vga_signals.N_188_0_0_0_cascade_\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__13385\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_1_0_2_cascade_\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__13382\,
            I => \N__13379\
        );

    \I__2232\ : InMux
    port map (
            O => \N__13379\,
            I => \N__13376\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__13376\,
            I => \N__13373\
        );

    \I__2230\ : Odrv12
    port map (
            O => \N__13373\,
            I => \this_vga_signals.g1_0_1\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__13370\,
            I => \N__13366\
        );

    \I__2228\ : InMux
    port map (
            O => \N__13369\,
            I => \N__13363\
        );

    \I__2227\ : InMux
    port map (
            O => \N__13366\,
            I => \N__13360\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__13363\,
            I => \N__13355\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__13360\,
            I => \N__13351\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__13359\,
            I => \N__13348\
        );

    \I__2223\ : CascadeMux
    port map (
            O => \N__13358\,
            I => \N__13345\
        );

    \I__2222\ : Span4Mux_v
    port map (
            O => \N__13355\,
            I => \N__13342\
        );

    \I__2221\ : InMux
    port map (
            O => \N__13354\,
            I => \N__13339\
        );

    \I__2220\ : Span4Mux_h
    port map (
            O => \N__13351\,
            I => \N__13336\
        );

    \I__2219\ : InMux
    port map (
            O => \N__13348\,
            I => \N__13331\
        );

    \I__2218\ : InMux
    port map (
            O => \N__13345\,
            I => \N__13331\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__13342\,
            I => \N_183_0\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__13339\,
            I => \N_183_0\
        );

    \I__2215\ : Odrv4
    port map (
            O => \N__13336\,
            I => \N_183_0\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__13331\,
            I => \N_183_0\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__13322\,
            I => \N__13318\
        );

    \I__2212\ : InMux
    port map (
            O => \N__13321\,
            I => \N__13311\
        );

    \I__2211\ : InMux
    port map (
            O => \N__13318\,
            I => \N__13307\
        );

    \I__2210\ : InMux
    port map (
            O => \N__13317\,
            I => \N__13304\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__13316\,
            I => \N__13301\
        );

    \I__2208\ : InMux
    port map (
            O => \N__13315\,
            I => \N__13298\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__13314\,
            I => \N__13294\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__13311\,
            I => \N__13289\
        );

    \I__2205\ : InMux
    port map (
            O => \N__13310\,
            I => \N__13286\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__13307\,
            I => \N__13281\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__13304\,
            I => \N__13281\
        );

    \I__2202\ : InMux
    port map (
            O => \N__13301\,
            I => \N__13278\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__13298\,
            I => \N__13275\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__13297\,
            I => \N__13272\
        );

    \I__2199\ : InMux
    port map (
            O => \N__13294\,
            I => \N__13268\
        );

    \I__2198\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13265\
        );

    \I__2197\ : InMux
    port map (
            O => \N__13292\,
            I => \N__13262\
        );

    \I__2196\ : Span4Mux_h
    port map (
            O => \N__13289\,
            I => \N__13259\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__13286\,
            I => \N__13250\
        );

    \I__2194\ : Span4Mux_h
    port map (
            O => \N__13281\,
            I => \N__13250\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__13278\,
            I => \N__13250\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__13275\,
            I => \N__13250\
        );

    \I__2191\ : InMux
    port map (
            O => \N__13272\,
            I => \N__13245\
        );

    \I__2190\ : InMux
    port map (
            O => \N__13271\,
            I => \N__13245\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__13268\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__13265\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__13262\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2186\ : Odrv4
    port map (
            O => \N__13259\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2185\ : Odrv4
    port map (
            O => \N__13250\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__13245\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__2183\ : InMux
    port map (
            O => \N__13232\,
            I => \N__13229\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__13229\,
            I => \this_vga_signals.mult1_un40_sum_0_axb1_i\
        );

    \I__2181\ : InMux
    port map (
            O => \N__13226\,
            I => \N__13223\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__13223\,
            I => \this_vga_signals.mult1_un40_sum_1_axb1\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__13220\,
            I => \this_vga_signals.mult1_un40_sum_m_x0_1_cascade_\
        );

    \I__2178\ : InMux
    port map (
            O => \N__13217\,
            I => \N__13214\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__13214\,
            I => \this_vga_signals.mult1_un40_sum_m_x1_1\
        );

    \I__2176\ : InMux
    port map (
            O => \N__13211\,
            I => \N__13208\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__13208\,
            I => \N__13203\
        );

    \I__2174\ : InMux
    port map (
            O => \N__13207\,
            I => \N__13200\
        );

    \I__2173\ : InMux
    port map (
            O => \N__13206\,
            I => \N__13197\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__13203\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_1\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__13200\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_1\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__13197\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_1\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__13190\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_1_cascade_\
        );

    \I__2168\ : InMux
    port map (
            O => \N__13187\,
            I => \N__13184\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__13184\,
            I => \N__13181\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__13181\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1\
        );

    \I__2165\ : InMux
    port map (
            O => \N__13178\,
            I => \N__13175\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__13175\,
            I => \N__13170\
        );

    \I__2163\ : InMux
    port map (
            O => \N__13174\,
            I => \N__13165\
        );

    \I__2162\ : InMux
    port map (
            O => \N__13173\,
            I => \N__13165\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__13170\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__13165\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\
        );

    \I__2159\ : InMux
    port map (
            O => \N__13160\,
            I => \N__13156\
        );

    \I__2158\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13150\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__13156\,
            I => \N__13147\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__13155\,
            I => \N__13142\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__13154\,
            I => \N__13139\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__13153\,
            I => \N__13136\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__13150\,
            I => \N__13131\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__13147\,
            I => \N__13131\
        );

    \I__2151\ : InMux
    port map (
            O => \N__13146\,
            I => \N__13128\
        );

    \I__2150\ : InMux
    port map (
            O => \N__13145\,
            I => \N__13119\
        );

    \I__2149\ : InMux
    port map (
            O => \N__13142\,
            I => \N__13119\
        );

    \I__2148\ : InMux
    port map (
            O => \N__13139\,
            I => \N__13119\
        );

    \I__2147\ : InMux
    port map (
            O => \N__13136\,
            I => \N__13119\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__13131\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__13128\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__13119\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__2143\ : InMux
    port map (
            O => \N__13112\,
            I => \N__13108\
        );

    \I__2142\ : InMux
    port map (
            O => \N__13111\,
            I => \N__13104\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__13108\,
            I => \N__13101\
        );

    \I__2140\ : InMux
    port map (
            O => \N__13107\,
            I => \N__13098\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__13104\,
            I => \N__13095\
        );

    \I__2138\ : Span4Mux_h
    port map (
            O => \N__13101\,
            I => \N__13092\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__13098\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__13095\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__13092\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__2134\ : InMux
    port map (
            O => \N__13085\,
            I => \N__13082\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__13082\,
            I => \N__13077\
        );

    \I__2132\ : InMux
    port map (
            O => \N__13081\,
            I => \N__13072\
        );

    \I__2131\ : InMux
    port map (
            O => \N__13080\,
            I => \N__13072\
        );

    \I__2130\ : Odrv12
    port map (
            O => \N__13077\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__13072\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__2128\ : InMux
    port map (
            O => \N__13067\,
            I => \N__13060\
        );

    \I__2127\ : InMux
    port map (
            O => \N__13066\,
            I => \N__13060\
        );

    \I__2126\ : InMux
    port map (
            O => \N__13065\,
            I => \N__13057\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__13060\,
            I => \N__13054\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__13057\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__13054\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__2122\ : InMux
    port map (
            O => \N__13049\,
            I => \N__13046\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__13046\,
            I => \N__13042\
        );

    \I__2120\ : InMux
    port map (
            O => \N__13045\,
            I => \N__13039\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__13042\,
            I => \N__13035\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__13039\,
            I => \N__13032\
        );

    \I__2117\ : InMux
    port map (
            O => \N__13038\,
            I => \N__13029\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__13035\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__2115\ : Odrv12
    port map (
            O => \N__13032\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__13029\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__2113\ : InMux
    port map (
            O => \N__13022\,
            I => \N__13011\
        );

    \I__2112\ : InMux
    port map (
            O => \N__13021\,
            I => \N__13011\
        );

    \I__2111\ : InMux
    port map (
            O => \N__13020\,
            I => \N__13000\
        );

    \I__2110\ : InMux
    port map (
            O => \N__13019\,
            I => \N__13000\
        );

    \I__2109\ : InMux
    port map (
            O => \N__13018\,
            I => \N__13000\
        );

    \I__2108\ : InMux
    port map (
            O => \N__13017\,
            I => \N__13000\
        );

    \I__2107\ : InMux
    port map (
            O => \N__13016\,
            I => \N__13000\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__13011\,
            I => \N__12994\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__13000\,
            I => \N__12994\
        );

    \I__2104\ : InMux
    port map (
            O => \N__12999\,
            I => \N__12988\
        );

    \I__2103\ : Span4Mux_h
    port map (
            O => \N__12994\,
            I => \N__12985\
        );

    \I__2102\ : InMux
    port map (
            O => \N__12993\,
            I => \N__12982\
        );

    \I__2101\ : InMux
    port map (
            O => \N__12992\,
            I => \N__12977\
        );

    \I__2100\ : InMux
    port map (
            O => \N__12991\,
            I => \N__12977\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__12988\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__2098\ : Odrv4
    port map (
            O => \N__12985\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__12982\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__12977\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__2095\ : InMux
    port map (
            O => \N__12968\,
            I => \N__12962\
        );

    \I__2094\ : InMux
    port map (
            O => \N__12967\,
            I => \N__12962\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__12962\,
            I => \N__12958\
        );

    \I__2092\ : InMux
    port map (
            O => \N__12961\,
            I => \N__12955\
        );

    \I__2091\ : Span4Mux_h
    port map (
            O => \N__12958\,
            I => \N__12952\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__12955\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__12952\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__2088\ : InMux
    port map (
            O => \N__12947\,
            I => \N__12944\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__12944\,
            I => \N__12939\
        );

    \I__2086\ : InMux
    port map (
            O => \N__12943\,
            I => \N__12936\
        );

    \I__2085\ : InMux
    port map (
            O => \N__12942\,
            I => \N__12933\
        );

    \I__2084\ : Span4Mux_h
    port map (
            O => \N__12939\,
            I => \N__12930\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__12936\,
            I => \N__12925\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__12933\,
            I => \N__12925\
        );

    \I__2081\ : Span4Mux_v
    port map (
            O => \N__12930\,
            I => \N__12922\
        );

    \I__2080\ : Span4Mux_v
    port map (
            O => \N__12925\,
            I => \N__12919\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__12922\,
            I => \this_vga_signals.N_188_0\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__12919\,
            I => \this_vga_signals.N_188_0\
        );

    \I__2077\ : InMux
    port map (
            O => \N__12914\,
            I => \N__12911\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__12911\,
            I => \N__12908\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__12908\,
            I => \this_vga_signals.M_this_vga_ramdac_en_i_o2_0_0\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__12905\,
            I => \this_vga_signals.M_this_vga_ramdac_en_i_o2_0_0_cascade_\
        );

    \I__2073\ : InMux
    port map (
            O => \N__12902\,
            I => \N__12898\
        );

    \I__2072\ : InMux
    port map (
            O => \N__12901\,
            I => \N__12895\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__12898\,
            I => \this_vga_signals.g1_4\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__12895\,
            I => \this_vga_signals.g1_4\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__12890\,
            I => \N__12887\
        );

    \I__2068\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12881\
        );

    \I__2067\ : InMux
    port map (
            O => \N__12886\,
            I => \N__12881\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__12881\,
            I => \N__12878\
        );

    \I__2065\ : Span4Mux_v
    port map (
            O => \N__12878\,
            I => \N__12874\
        );

    \I__2064\ : InMux
    port map (
            O => \N__12877\,
            I => \N__12871\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__12874\,
            I => \this_vga_signals.mult1_un61_sum_s_3\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__12871\,
            I => \this_vga_signals.mult1_un61_sum_s_3\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__12866\,
            I => \N__12863\
        );

    \I__2060\ : InMux
    port map (
            O => \N__12863\,
            I => \N__12860\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__12860\,
            I => \this_vga_signals.mult1_un61_sum_i_3\
        );

    \I__2058\ : InMux
    port map (
            O => \N__12857\,
            I => \N__12853\
        );

    \I__2057\ : InMux
    port map (
            O => \N__12856\,
            I => \N__12848\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__12853\,
            I => \N__12845\
        );

    \I__2055\ : InMux
    port map (
            O => \N__12852\,
            I => \N__12840\
        );

    \I__2054\ : InMux
    port map (
            O => \N__12851\,
            I => \N__12840\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__12848\,
            I => \this_vga_signals.if_N_3_mux\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__12845\,
            I => \this_vga_signals.if_N_3_mux\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__12840\,
            I => \this_vga_signals.if_N_3_mux\
        );

    \I__2050\ : InMux
    port map (
            O => \N__12833\,
            I => \N__12830\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__12830\,
            I => \N__12826\
        );

    \I__2048\ : InMux
    port map (
            O => \N__12829\,
            I => \N__12823\
        );

    \I__2047\ : Odrv4
    port map (
            O => \N__12826\,
            I => \this_vga_signals.g6_0\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__12823\,
            I => \this_vga_signals.g6_0\
        );

    \I__2045\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12812\
        );

    \I__2044\ : InMux
    port map (
            O => \N__12817\,
            I => \N__12809\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__12816\,
            I => \N__12801\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__12815\,
            I => \N__12798\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__12812\,
            I => \N__12795\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__12809\,
            I => \N__12792\
        );

    \I__2039\ : InMux
    port map (
            O => \N__12808\,
            I => \N__12789\
        );

    \I__2038\ : InMux
    port map (
            O => \N__12807\,
            I => \N__12786\
        );

    \I__2037\ : InMux
    port map (
            O => \N__12806\,
            I => \N__12783\
        );

    \I__2036\ : InMux
    port map (
            O => \N__12805\,
            I => \N__12774\
        );

    \I__2035\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12774\
        );

    \I__2034\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12774\
        );

    \I__2033\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12774\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__12795\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__12792\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__12789\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__12786\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__12783\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__12774\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__12761\,
            I => \N__12758\
        );

    \I__2025\ : InMux
    port map (
            O => \N__12758\,
            I => \N__12755\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__12755\,
            I => \N__12752\
        );

    \I__2023\ : Span4Mux_h
    port map (
            O => \N__12752\,
            I => \N__12749\
        );

    \I__2022\ : Span4Mux_v
    port map (
            O => \N__12749\,
            I => \N__12746\
        );

    \I__2021\ : Odrv4
    port map (
            O => \N__12746\,
            I => \M_this_vga_signals_address_13\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__12743\,
            I => \N__12740\
        );

    \I__2019\ : InMux
    port map (
            O => \N__12740\,
            I => \N__12737\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__12737\,
            I => \N__12734\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__12734\,
            I => \this_vga_signals.g0_0\
        );

    \I__2016\ : InMux
    port map (
            O => \N__12731\,
            I => \N__12728\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__12728\,
            I => \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0ASZ0\
        );

    \I__2014\ : InMux
    port map (
            O => \N__12725\,
            I => \N__12720\
        );

    \I__2013\ : InMux
    port map (
            O => \N__12724\,
            I => \N__12717\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__12723\,
            I => \N__12714\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__12720\,
            I => \N__12710\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__12717\,
            I => \N__12707\
        );

    \I__2009\ : InMux
    port map (
            O => \N__12714\,
            I => \N__12699\
        );

    \I__2008\ : InMux
    port map (
            O => \N__12713\,
            I => \N__12699\
        );

    \I__2007\ : Span4Mux_h
    port map (
            O => \N__12710\,
            I => \N__12694\
        );

    \I__2006\ : Span4Mux_h
    port map (
            O => \N__12707\,
            I => \N__12694\
        );

    \I__2005\ : InMux
    port map (
            O => \N__12706\,
            I => \N__12687\
        );

    \I__2004\ : InMux
    port map (
            O => \N__12705\,
            I => \N__12687\
        );

    \I__2003\ : InMux
    port map (
            O => \N__12704\,
            I => \N__12687\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__12699\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__2001\ : Odrv4
    port map (
            O => \N__12694\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__12687\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1999\ : InMux
    port map (
            O => \N__12680\,
            I => \N__12674\
        );

    \I__1998\ : InMux
    port map (
            O => \N__12679\,
            I => \N__12674\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__12674\,
            I => \N__12670\
        );

    \I__1996\ : InMux
    port map (
            O => \N__12673\,
            I => \N__12667\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__12670\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__12667\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1993\ : InMux
    port map (
            O => \N__12662\,
            I => \N__12657\
        );

    \I__1992\ : InMux
    port map (
            O => \N__12661\,
            I => \N__12652\
        );

    \I__1991\ : InMux
    port map (
            O => \N__12660\,
            I => \N__12652\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__12657\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__12652\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__12647\,
            I => \this_vga_signals.g0_10_1_cascade_\
        );

    \I__1987\ : InMux
    port map (
            O => \N__12644\,
            I => \N__12641\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__12641\,
            I => \N__12636\
        );

    \I__1985\ : InMux
    port map (
            O => \N__12640\,
            I => \N__12633\
        );

    \I__1984\ : InMux
    port map (
            O => \N__12639\,
            I => \N__12625\
        );

    \I__1983\ : Span4Mux_h
    port map (
            O => \N__12636\,
            I => \N__12621\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__12633\,
            I => \N__12618\
        );

    \I__1981\ : InMux
    port map (
            O => \N__12632\,
            I => \N__12615\
        );

    \I__1980\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12606\
        );

    \I__1979\ : InMux
    port map (
            O => \N__12630\,
            I => \N__12606\
        );

    \I__1978\ : InMux
    port map (
            O => \N__12629\,
            I => \N__12606\
        );

    \I__1977\ : InMux
    port map (
            O => \N__12628\,
            I => \N__12606\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__12625\,
            I => \N__12603\
        );

    \I__1975\ : InMux
    port map (
            O => \N__12624\,
            I => \N__12600\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__12621\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__12618\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__12615\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__12606\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1\
        );

    \I__1970\ : Odrv4
    port map (
            O => \N__12603\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__12600\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1\
        );

    \I__1968\ : InMux
    port map (
            O => \N__12587\,
            I => \N__12584\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__12584\,
            I => \N__12581\
        );

    \I__1966\ : Span4Mux_h
    port map (
            O => \N__12581\,
            I => \N__12578\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__12578\,
            I => \this_vga_signals.if_N_18_1\
        );

    \I__1964\ : InMux
    port map (
            O => \N__12575\,
            I => \N__12572\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__12572\,
            I => \this_vga_signals.m48_i_x4_0\
        );

    \I__1962\ : InMux
    port map (
            O => \N__12569\,
            I => \N__12562\
        );

    \I__1961\ : InMux
    port map (
            O => \N__12568\,
            I => \N__12562\
        );

    \I__1960\ : InMux
    port map (
            O => \N__12567\,
            I => \N__12557\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__12562\,
            I => \N__12554\
        );

    \I__1958\ : InMux
    port map (
            O => \N__12561\,
            I => \N__12545\
        );

    \I__1957\ : InMux
    port map (
            O => \N__12560\,
            I => \N__12542\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__12557\,
            I => \N__12539\
        );

    \I__1955\ : Span4Mux_v
    port map (
            O => \N__12554\,
            I => \N__12529\
        );

    \I__1954\ : InMux
    port map (
            O => \N__12553\,
            I => \N__12522\
        );

    \I__1953\ : InMux
    port map (
            O => \N__12552\,
            I => \N__12522\
        );

    \I__1952\ : InMux
    port map (
            O => \N__12551\,
            I => \N__12522\
        );

    \I__1951\ : InMux
    port map (
            O => \N__12550\,
            I => \N__12515\
        );

    \I__1950\ : InMux
    port map (
            O => \N__12549\,
            I => \N__12515\
        );

    \I__1949\ : InMux
    port map (
            O => \N__12548\,
            I => \N__12515\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__12545\,
            I => \N__12510\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__12542\,
            I => \N__12510\
        );

    \I__1946\ : Span4Mux_h
    port map (
            O => \N__12539\,
            I => \N__12507\
        );

    \I__1945\ : InMux
    port map (
            O => \N__12538\,
            I => \N__12498\
        );

    \I__1944\ : InMux
    port map (
            O => \N__12537\,
            I => \N__12498\
        );

    \I__1943\ : InMux
    port map (
            O => \N__12536\,
            I => \N__12498\
        );

    \I__1942\ : InMux
    port map (
            O => \N__12535\,
            I => \N__12498\
        );

    \I__1941\ : InMux
    port map (
            O => \N__12534\,
            I => \N__12491\
        );

    \I__1940\ : InMux
    port map (
            O => \N__12533\,
            I => \N__12491\
        );

    \I__1939\ : InMux
    port map (
            O => \N__12532\,
            I => \N__12491\
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__12529\,
            I => \this_vga_signals.mult1_un47_sum_c3_0\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__12522\,
            I => \this_vga_signals.mult1_un47_sum_c3_0\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__12515\,
            I => \this_vga_signals.mult1_un47_sum_c3_0\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__12510\,
            I => \this_vga_signals.mult1_un47_sum_c3_0\
        );

    \I__1934\ : Odrv4
    port map (
            O => \N__12507\,
            I => \this_vga_signals.mult1_un47_sum_c3_0\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__12498\,
            I => \this_vga_signals.mult1_un47_sum_c3_0\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__12491\,
            I => \this_vga_signals.mult1_un47_sum_c3_0\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__12476\,
            I => \N__12473\
        );

    \I__1930\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12470\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__12470\,
            I => \this_vga_signals.g4_1_0\
        );

    \I__1928\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12461\
        );

    \I__1927\ : InMux
    port map (
            O => \N__12466\,
            I => \N__12461\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__12461\,
            I => \N__12458\
        );

    \I__1925\ : Span4Mux_h
    port map (
            O => \N__12458\,
            I => \N__12453\
        );

    \I__1924\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12448\
        );

    \I__1923\ : InMux
    port map (
            O => \N__12456\,
            I => \N__12448\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__12453\,
            I => \this_vga_signals.g0_1\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__12448\,
            I => \this_vga_signals.g0_1\
        );

    \I__1920\ : InMux
    port map (
            O => \N__12443\,
            I => \this_vga_signals.mult1_un68_sum_cry_0\
        );

    \I__1919\ : InMux
    port map (
            O => \N__12440\,
            I => \N__12437\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__12437\,
            I => \N__12434\
        );

    \I__1917\ : Span12Mux_h
    port map (
            O => \N__12434\,
            I => \N__12431\
        );

    \I__1916\ : Odrv12
    port map (
            O => \N__12431\,
            I => \this_vga_signals.mult1_un61_sum_cry_1_s\
        );

    \I__1915\ : InMux
    port map (
            O => \N__12428\,
            I => \this_vga_signals.mult1_un68_sum_cry_1\
        );

    \I__1914\ : InMux
    port map (
            O => \N__12425\,
            I => \N__12422\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__12422\,
            I => \N__12419\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__12419\,
            I => \N__12416\
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__12416\,
            I => \this_vga_signals.mult1_un68_sum_axb_3\
        );

    \I__1910\ : InMux
    port map (
            O => \N__12413\,
            I => \this_vga_signals.mult1_un68_sum_cry_2\
        );

    \I__1909\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12407\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__12407\,
            I => \N__12401\
        );

    \I__1907\ : InMux
    port map (
            O => \N__12406\,
            I => \N__12398\
        );

    \I__1906\ : InMux
    port map (
            O => \N__12405\,
            I => \N__12395\
        );

    \I__1905\ : InMux
    port map (
            O => \N__12404\,
            I => \N__12392\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__12401\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__12398\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__12395\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__12392\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__1900\ : InMux
    port map (
            O => \N__12383\,
            I => \N__12380\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__12380\,
            I => \this_vga_signals.N_3_2\
        );

    \I__1898\ : InMux
    port map (
            O => \N__12377\,
            I => \N__12369\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__12376\,
            I => \N__12358\
        );

    \I__1896\ : InMux
    port map (
            O => \N__12375\,
            I => \N__12348\
        );

    \I__1895\ : InMux
    port map (
            O => \N__12374\,
            I => \N__12348\
        );

    \I__1894\ : InMux
    port map (
            O => \N__12373\,
            I => \N__12348\
        );

    \I__1893\ : InMux
    port map (
            O => \N__12372\,
            I => \N__12348\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__12369\,
            I => \N__12345\
        );

    \I__1891\ : InMux
    port map (
            O => \N__12368\,
            I => \N__12340\
        );

    \I__1890\ : InMux
    port map (
            O => \N__12367\,
            I => \N__12340\
        );

    \I__1889\ : InMux
    port map (
            O => \N__12366\,
            I => \N__12337\
        );

    \I__1888\ : InMux
    port map (
            O => \N__12365\,
            I => \N__12330\
        );

    \I__1887\ : InMux
    port map (
            O => \N__12364\,
            I => \N__12330\
        );

    \I__1886\ : InMux
    port map (
            O => \N__12363\,
            I => \N__12330\
        );

    \I__1885\ : InMux
    port map (
            O => \N__12362\,
            I => \N__12323\
        );

    \I__1884\ : InMux
    port map (
            O => \N__12361\,
            I => \N__12323\
        );

    \I__1883\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12323\
        );

    \I__1882\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12320\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__12348\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__12345\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__12340\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__12337\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__12330\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__12323\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__12320\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__1874\ : InMux
    port map (
            O => \N__12305\,
            I => \N__12302\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__12302\,
            I => \this_vga_signals.g0_16_x1\
        );

    \I__1872\ : InMux
    port map (
            O => \N__12299\,
            I => \N__12295\
        );

    \I__1871\ : InMux
    port map (
            O => \N__12298\,
            I => \N__12292\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__12295\,
            I => \this_vga_signals.N_81_1\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__12292\,
            I => \this_vga_signals.N_81_1\
        );

    \I__1868\ : InMux
    port map (
            O => \N__12287\,
            I => \N__12284\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__12284\,
            I => \this_vga_signals.g1_2\
        );

    \I__1866\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12277\
        );

    \I__1865\ : InMux
    port map (
            O => \N__12280\,
            I => \N__12274\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__12277\,
            I => \this_vga_signals.if_N_7_i\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__12274\,
            I => \this_vga_signals.if_N_7_i\
        );

    \I__1862\ : InMux
    port map (
            O => \N__12269\,
            I => \N__12265\
        );

    \I__1861\ : InMux
    port map (
            O => \N__12268\,
            I => \N__12262\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__12265\,
            I => \this_vga_signals.if_N_11\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__12262\,
            I => \this_vga_signals.if_N_11\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__12257\,
            I => \this_vga_signals.if_i3_mux_0_1_cascade_\
        );

    \I__1857\ : InMux
    port map (
            O => \N__12254\,
            I => \N__12251\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__12251\,
            I => \this_vga_signals.m48_i_x4_3\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__12248\,
            I => \N__12245\
        );

    \I__1854\ : InMux
    port map (
            O => \N__12245\,
            I => \N__12242\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__12242\,
            I => \N__12239\
        );

    \I__1852\ : Odrv4
    port map (
            O => \N__12239\,
            I => \this_vga_signals.if_i3_mux_0_1\
        );

    \I__1851\ : InMux
    port map (
            O => \N__12236\,
            I => \N__12230\
        );

    \I__1850\ : InMux
    port map (
            O => \N__12235\,
            I => \N__12230\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__12230\,
            I => \this_vga_signals.mult1_un68_sum_axb1_0_0\
        );

    \I__1848\ : InMux
    port map (
            O => \N__12227\,
            I => \N__12224\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__12224\,
            I => \this_vga_signals.N_57_0\
        );

    \I__1846\ : InMux
    port map (
            O => \N__12221\,
            I => \N__12218\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__12218\,
            I => \this_vga_signals.N_57_i_i_0\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__12215\,
            I => \this_vga_signals.g1_0_cascade_\
        );

    \I__1843\ : InMux
    port map (
            O => \N__12212\,
            I => \N__12209\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__12209\,
            I => \this_vga_signals.if_N_6_mux_0_0_0\
        );

    \I__1841\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12203\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__12203\,
            I => \this_vga_signals.g2_1_0_0\
        );

    \I__1839\ : InMux
    port map (
            O => \N__12200\,
            I => \N__12195\
        );

    \I__1838\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12184\
        );

    \I__1837\ : InMux
    port map (
            O => \N__12198\,
            I => \N__12184\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__12195\,
            I => \N__12181\
        );

    \I__1835\ : InMux
    port map (
            O => \N__12194\,
            I => \N__12176\
        );

    \I__1834\ : InMux
    port map (
            O => \N__12193\,
            I => \N__12176\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__12192\,
            I => \N__12161\
        );

    \I__1832\ : InMux
    port map (
            O => \N__12191\,
            I => \N__12156\
        );

    \I__1831\ : InMux
    port map (
            O => \N__12190\,
            I => \N__12156\
        );

    \I__1830\ : InMux
    port map (
            O => \N__12189\,
            I => \N__12153\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__12184\,
            I => \N__12150\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__12181\,
            I => \N__12145\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__12176\,
            I => \N__12145\
        );

    \I__1826\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12140\
        );

    \I__1825\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12140\
        );

    \I__1824\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12137\
        );

    \I__1823\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12126\
        );

    \I__1822\ : InMux
    port map (
            O => \N__12171\,
            I => \N__12126\
        );

    \I__1821\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12126\
        );

    \I__1820\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12126\
        );

    \I__1819\ : InMux
    port map (
            O => \N__12168\,
            I => \N__12126\
        );

    \I__1818\ : InMux
    port map (
            O => \N__12167\,
            I => \N__12117\
        );

    \I__1817\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12117\
        );

    \I__1816\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12117\
        );

    \I__1815\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12117\
        );

    \I__1814\ : InMux
    port map (
            O => \N__12161\,
            I => \N__12114\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__12156\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__12153\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__12150\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__12145\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__12140\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__12137\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__12126\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__12117\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__12114\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1804\ : InMux
    port map (
            O => \N__12095\,
            I => \N__12092\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__12092\,
            I => \N__12085\
        );

    \I__1802\ : InMux
    port map (
            O => \N__12091\,
            I => \N__12079\
        );

    \I__1801\ : InMux
    port map (
            O => \N__12090\,
            I => \N__12074\
        );

    \I__1800\ : InMux
    port map (
            O => \N__12089\,
            I => \N__12074\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__12088\,
            I => \N__12062\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__12085\,
            I => \N__12058\
        );

    \I__1797\ : InMux
    port map (
            O => \N__12084\,
            I => \N__12053\
        );

    \I__1796\ : InMux
    port map (
            O => \N__12083\,
            I => \N__12053\
        );

    \I__1795\ : InMux
    port map (
            O => \N__12082\,
            I => \N__12050\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__12079\,
            I => \N__12047\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__12074\,
            I => \N__12044\
        );

    \I__1792\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12041\
        );

    \I__1791\ : InMux
    port map (
            O => \N__12072\,
            I => \N__12036\
        );

    \I__1790\ : InMux
    port map (
            O => \N__12071\,
            I => \N__12036\
        );

    \I__1789\ : InMux
    port map (
            O => \N__12070\,
            I => \N__12029\
        );

    \I__1788\ : InMux
    port map (
            O => \N__12069\,
            I => \N__12029\
        );

    \I__1787\ : InMux
    port map (
            O => \N__12068\,
            I => \N__12029\
        );

    \I__1786\ : InMux
    port map (
            O => \N__12067\,
            I => \N__12020\
        );

    \I__1785\ : InMux
    port map (
            O => \N__12066\,
            I => \N__12020\
        );

    \I__1784\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12020\
        );

    \I__1783\ : InMux
    port map (
            O => \N__12062\,
            I => \N__12020\
        );

    \I__1782\ : InMux
    port map (
            O => \N__12061\,
            I => \N__12017\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__12058\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__12053\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__12050\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__12047\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1777\ : Odrv4
    port map (
            O => \N__12044\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__12041\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__12036\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__12029\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__12020\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__12017\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11996\,
            I => \N__11992\
        );

    \I__1770\ : CascadeMux
    port map (
            O => \N__11995\,
            I => \N__11989\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__11992\,
            I => \N__11986\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11989\,
            I => \N__11983\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__11986\,
            I => \this_vga_signals.N_5_i_1_0\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__11983\,
            I => \this_vga_signals.N_5_i_1_0\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__11978\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_1_0_x1_cascade_\
        );

    \I__1764\ : InMux
    port map (
            O => \N__11975\,
            I => \N__11972\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__11972\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_1_0\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11969\,
            I => \N__11966\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__11966\,
            I => \this_vga_signals.mult1_un61_sum_ac0_2_2_1\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__11963\,
            I => \this_vga_signals.mult1_un61_sum_ac0_2_2_1_cascade_\
        );

    \I__1759\ : InMux
    port map (
            O => \N__11960\,
            I => \N__11957\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__11957\,
            I => \N__11950\
        );

    \I__1757\ : InMux
    port map (
            O => \N__11956\,
            I => \N__11943\
        );

    \I__1756\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11943\
        );

    \I__1755\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11943\
        );

    \I__1754\ : InMux
    port map (
            O => \N__11953\,
            I => \N__11940\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__11950\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__11943\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__11940\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0
        );

    \I__1750\ : InMux
    port map (
            O => \N__11933\,
            I => \N__11930\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__11930\,
            I => \N__11926\
        );

    \I__1748\ : InMux
    port map (
            O => \N__11929\,
            I => \N__11923\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__11926\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__11923\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__1745\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11909\
        );

    \I__1744\ : InMux
    port map (
            O => \N__11917\,
            I => \N__11909\
        );

    \I__1743\ : InMux
    port map (
            O => \N__11916\,
            I => \N__11909\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__11909\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_2\
        );

    \I__1741\ : InMux
    port map (
            O => \N__11906\,
            I => \N__11903\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__11903\,
            I => \this_vga_signals.mult1_un61_sum_ac0_sx\
        );

    \I__1739\ : InMux
    port map (
            O => \N__11900\,
            I => \N__11896\
        );

    \I__1738\ : InMux
    port map (
            O => \N__11899\,
            I => \N__11893\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__11896\,
            I => \this_vga_signals.mult1_un61_sum_ac0_2_4_tz\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__11893\,
            I => \this_vga_signals.mult1_un61_sum_ac0_2_4_tz\
        );

    \I__1735\ : InMux
    port map (
            O => \N__11888\,
            I => \N__11884\
        );

    \I__1734\ : InMux
    port map (
            O => \N__11887\,
            I => \N__11881\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__11884\,
            I => \N__11874\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__11881\,
            I => \N__11874\
        );

    \I__1731\ : InMux
    port map (
            O => \N__11880\,
            I => \N__11871\
        );

    \I__1730\ : InMux
    port map (
            O => \N__11879\,
            I => \N__11868\
        );

    \I__1729\ : Odrv4
    port map (
            O => \N__11874\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__11871\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__11868\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__11861\,
            I => \this_vga_signals.mult1_un61_sum_ac0_2_cascade_\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11858\,
            I => \N__11854\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__11857\,
            I => \N__11850\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__11854\,
            I => \N__11845\
        );

    \I__1722\ : InMux
    port map (
            O => \N__11853\,
            I => \N__11841\
        );

    \I__1721\ : InMux
    port map (
            O => \N__11850\,
            I => \N__11836\
        );

    \I__1720\ : InMux
    port map (
            O => \N__11849\,
            I => \N__11836\
        );

    \I__1719\ : InMux
    port map (
            O => \N__11848\,
            I => \N__11832\
        );

    \I__1718\ : Span4Mux_v
    port map (
            O => \N__11845\,
            I => \N__11826\
        );

    \I__1717\ : InMux
    port map (
            O => \N__11844\,
            I => \N__11823\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__11841\,
            I => \N__11820\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__11836\,
            I => \N__11817\
        );

    \I__1714\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11814\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__11832\,
            I => \N__11811\
        );

    \I__1712\ : InMux
    port map (
            O => \N__11831\,
            I => \N__11806\
        );

    \I__1711\ : InMux
    port map (
            O => \N__11830\,
            I => \N__11806\
        );

    \I__1710\ : InMux
    port map (
            O => \N__11829\,
            I => \N__11803\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__11826\,
            I => this_vga_signals_un4_lcounter_if_i3_mux
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__11823\,
            I => this_vga_signals_un4_lcounter_if_i3_mux
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__11820\,
            I => this_vga_signals_un4_lcounter_if_i3_mux
        );

    \I__1706\ : Odrv4
    port map (
            O => \N__11817\,
            I => this_vga_signals_un4_lcounter_if_i3_mux
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__11814\,
            I => this_vga_signals_un4_lcounter_if_i3_mux
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__11811\,
            I => this_vga_signals_un4_lcounter_if_i3_mux
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__11806\,
            I => this_vga_signals_un4_lcounter_if_i3_mux
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__11803\,
            I => this_vga_signals_un4_lcounter_if_i3_mux
        );

    \I__1701\ : InMux
    port map (
            O => \N__11786\,
            I => \N__11783\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__11783\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__1699\ : InMux
    port map (
            O => \N__11780\,
            I => \N__11777\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__11777\,
            I => \this_delay_clk.M_pipe_qZ0Z_2\
        );

    \I__1697\ : InMux
    port map (
            O => \N__11774\,
            I => \N__11771\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__11771\,
            I => \this_delay_clk.M_pipe_qZ0Z_3\
        );

    \I__1695\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11764\
        );

    \I__1694\ : InMux
    port map (
            O => \N__11767\,
            I => \N__11761\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__11764\,
            I => \this_vga_signals.N_81_0\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__11761\,
            I => \this_vga_signals.N_81_0\
        );

    \I__1691\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11749\
        );

    \I__1690\ : InMux
    port map (
            O => \N__11755\,
            I => \N__11749\
        );

    \I__1689\ : InMux
    port map (
            O => \N__11754\,
            I => \N__11746\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__11749\,
            I => \N__11743\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__11746\,
            I => \this_vga_signals.N_370_0\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__11743\,
            I => \this_vga_signals.N_370_0\
        );

    \I__1685\ : InMux
    port map (
            O => \N__11738\,
            I => \N__11735\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__11735\,
            I => \this_vga_signals.mult1_un40_sum1_2\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__11732\,
            I => \N__11729\
        );

    \I__1682\ : InMux
    port map (
            O => \N__11729\,
            I => \N__11716\
        );

    \I__1681\ : InMux
    port map (
            O => \N__11728\,
            I => \N__11716\
        );

    \I__1680\ : InMux
    port map (
            O => \N__11727\,
            I => \N__11716\
        );

    \I__1679\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11716\
        );

    \I__1678\ : InMux
    port map (
            O => \N__11725\,
            I => \N__11712\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__11716\,
            I => \N__11709\
        );

    \I__1676\ : InMux
    port map (
            O => \N__11715\,
            I => \N__11706\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__11712\,
            I => \this_vga_signals_M_vcounter_q_7_rep1\
        );

    \I__1674\ : Odrv4
    port map (
            O => \N__11709\,
            I => \this_vga_signals_M_vcounter_q_7_rep1\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__11706\,
            I => \this_vga_signals_M_vcounter_q_7_rep1\
        );

    \I__1672\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11685\
        );

    \I__1671\ : InMux
    port map (
            O => \N__11698\,
            I => \N__11685\
        );

    \I__1670\ : InMux
    port map (
            O => \N__11697\,
            I => \N__11685\
        );

    \I__1669\ : InMux
    port map (
            O => \N__11696\,
            I => \N__11685\
        );

    \I__1668\ : InMux
    port map (
            O => \N__11695\,
            I => \N__11680\
        );

    \I__1667\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11680\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__11685\,
            I => \this_vga_signals_M_vcounter_q_8_rep1\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__11680\,
            I => \this_vga_signals_M_vcounter_q_8_rep1\
        );

    \I__1664\ : InMux
    port map (
            O => \N__11675\,
            I => \N__11671\
        );

    \I__1663\ : InMux
    port map (
            O => \N__11674\,
            I => \N__11668\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__11671\,
            I => \this_vga_signals.N_330_0\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__11668\,
            I => \this_vga_signals.N_330_0\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__11663\,
            I => \N__11660\
        );

    \I__1659\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11657\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__11657\,
            I => \N__11654\
        );

    \I__1657\ : Span4Mux_v
    port map (
            O => \N__11654\,
            I => \N__11651\
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__11651\,
            I => \this_vga_signals.vsync_1_0_a2_6_a2_0\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__11648\,
            I => \this_vga_signals.if_m11_1_cascade_\
        );

    \I__1654\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11642\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__11642\,
            I => \N__11639\
        );

    \I__1652\ : Span4Mux_h
    port map (
            O => \N__11639\,
            I => \N__11636\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__11636\,
            I => \this_vga_signals.mult1_un47_sum_i_0\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__11633\,
            I => \this_vga_signals.mult1_un61_sum_ac0_2_2_cascade_\
        );

    \I__1649\ : InMux
    port map (
            O => \N__11630\,
            I => \N__11627\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__11627\,
            I => \N__11624\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__11624\,
            I => \this_vga_signals.mult1_un61_sum_axb2_i\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__11621\,
            I => \N__11617\
        );

    \I__1645\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11613\
        );

    \I__1644\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11610\
        );

    \I__1643\ : InMux
    port map (
            O => \N__11616\,
            I => \N__11606\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__11613\,
            I => \N__11603\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__11610\,
            I => \N__11600\
        );

    \I__1640\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11597\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__11606\,
            I => \N__11592\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__11603\,
            I => \N__11585\
        );

    \I__1637\ : Span4Mux_h
    port map (
            O => \N__11600\,
            I => \N__11585\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__11597\,
            I => \N__11585\
        );

    \I__1635\ : InMux
    port map (
            O => \N__11596\,
            I => \N__11580\
        );

    \I__1634\ : InMux
    port map (
            O => \N__11595\,
            I => \N__11580\
        );

    \I__1633\ : Odrv4
    port map (
            O => \N__11592\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__11585\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__11580\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__11573\,
            I => \N__11570\
        );

    \I__1629\ : InMux
    port map (
            O => \N__11570\,
            I => \N__11564\
        );

    \I__1628\ : InMux
    port map (
            O => \N__11569\,
            I => \N__11564\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__11564\,
            I => \this_vga_signals.if_m5_0_1\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__11561\,
            I => \N__11558\
        );

    \I__1625\ : InMux
    port map (
            O => \N__11558\,
            I => \N__11554\
        );

    \I__1624\ : InMux
    port map (
            O => \N__11557\,
            I => \N__11551\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__11554\,
            I => \N__11548\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__11551\,
            I => \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41Z0Z_1\
        );

    \I__1621\ : Odrv4
    port map (
            O => \N__11548\,
            I => \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41Z0Z_1\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__11543\,
            I => \this_vga_signals.mult1_un40_sum_0_axb1_i_cascade_\
        );

    \I__1619\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11535\
        );

    \I__1618\ : InMux
    port map (
            O => \N__11539\,
            I => \N__11530\
        );

    \I__1617\ : InMux
    port map (
            O => \N__11538\,
            I => \N__11530\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__11535\,
            I => \this_vga_signals.mult1_un47_sum_ac0_1\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__11530\,
            I => \this_vga_signals.mult1_un47_sum_ac0_1\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__11525\,
            I => \N__11521\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__11524\,
            I => \N__11517\
        );

    \I__1612\ : InMux
    port map (
            O => \N__11521\,
            I => \N__11512\
        );

    \I__1611\ : InMux
    port map (
            O => \N__11520\,
            I => \N__11512\
        );

    \I__1610\ : InMux
    port map (
            O => \N__11517\,
            I => \N__11509\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__11512\,
            I => \N__11506\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__11509\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_c\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__11506\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_c\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__11501\,
            I => \N_475_cascade_\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__11498\,
            I => \this_vga_signals.if_N_3_mux_cascade_\
        );

    \I__1604\ : InMux
    port map (
            O => \N__11495\,
            I => \N__11491\
        );

    \I__1603\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11488\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__11491\,
            I => \N__11483\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__11488\,
            I => \N__11483\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__11483\,
            I => \this_vga_signals.mult1_un47_sum_axb2_0\
        );

    \I__1599\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11477\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__11477\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_x1\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__11474\,
            I => \this_vga_signals.mult1_un47_sum_axb2_0_cascade_\
        );

    \I__1596\ : InMux
    port map (
            O => \N__11471\,
            I => \N__11468\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__11468\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_x0\
        );

    \I__1594\ : InMux
    port map (
            O => \N__11465\,
            I => \N__11459\
        );

    \I__1593\ : InMux
    port map (
            O => \N__11464\,
            I => \N__11459\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__11459\,
            I => \N__11456\
        );

    \I__1591\ : Odrv4
    port map (
            O => \N__11456\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__1590\ : InMux
    port map (
            O => \N__11453\,
            I => \N__11450\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__11450\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_1_0_x1\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__11447\,
            I => \N__11444\
        );

    \I__1587\ : InMux
    port map (
            O => \N__11444\,
            I => \N__11440\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__11443\,
            I => \N__11436\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__11440\,
            I => \N__11432\
        );

    \I__1584\ : InMux
    port map (
            O => \N__11439\,
            I => \N__11425\
        );

    \I__1583\ : InMux
    port map (
            O => \N__11436\,
            I => \N__11425\
        );

    \I__1582\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11425\
        );

    \I__1581\ : Odrv4
    port map (
            O => \N__11432\,
            I => \this_vga_signals_M_vcounter_q_fast_6\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__11425\,
            I => \this_vga_signals_M_vcounter_q_fast_6\
        );

    \I__1579\ : InMux
    port map (
            O => \N__11420\,
            I => \N__11417\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__11417\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_1_0_x0\
        );

    \I__1577\ : InMux
    port map (
            O => \N__11414\,
            I => \N__11411\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__11411\,
            I => \this_vga_signals.if_m10_0_a4_1_0_x1\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__11408\,
            I => \this_vga_signals.if_m10_0_a4_1_0_x0_cascade_\
        );

    \I__1574\ : InMux
    port map (
            O => \N__11405\,
            I => \N__11402\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__11402\,
            I => \this_vga_signals.if_m10_0_a4_1\
        );

    \I__1572\ : InMux
    port map (
            O => \N__11399\,
            I => \N__11394\
        );

    \I__1571\ : InMux
    port map (
            O => \N__11398\,
            I => \N__11391\
        );

    \I__1570\ : InMux
    port map (
            O => \N__11397\,
            I => \N__11388\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__11394\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__11391\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__11388\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__1566\ : InMux
    port map (
            O => \N__11381\,
            I => \N__11375\
        );

    \I__1565\ : InMux
    port map (
            O => \N__11380\,
            I => \N__11375\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__11375\,
            I => \this_vga_signals.g0_0_a3_0\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__11372\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNISGOSZ0Z_4_cascade_\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__11369\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1_x0_cascade_\
        );

    \I__1561\ : InMux
    port map (
            O => \N__11366\,
            I => \N__11363\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__11363\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1_x1\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__11360\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1_cascade_\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__11357\,
            I => \this_vga_signals.if_m10_0_x2_0_0_cascade_\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__11354\,
            I => \N__11351\
        );

    \I__1556\ : InMux
    port map (
            O => \N__11351\,
            I => \N__11348\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__11348\,
            I => \this_vga_signals.mult1_un47_sum_c2_0\
        );

    \I__1554\ : CascadeMux
    port map (
            O => \N__11345\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_\
        );

    \I__1553\ : CascadeMux
    port map (
            O => \N__11342\,
            I => \this_vga_signals.mult1_un47_sum_c3_0_cascade_\
        );

    \I__1552\ : InMux
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__11336\,
            I => \N__11333\
        );

    \I__1550\ : Odrv4
    port map (
            O => \N__11333\,
            I => \this_vga_signals.if_m2_1\
        );

    \I__1549\ : InMux
    port map (
            O => \N__11330\,
            I => \N__11326\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__11329\,
            I => \N__11321\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__11326\,
            I => \N__11318\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__11325\,
            I => \N__11315\
        );

    \I__1545\ : InMux
    port map (
            O => \N__11324\,
            I => \N__11311\
        );

    \I__1544\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11308\
        );

    \I__1543\ : Span4Mux_v
    port map (
            O => \N__11318\,
            I => \N__11305\
        );

    \I__1542\ : InMux
    port map (
            O => \N__11315\,
            I => \N__11300\
        );

    \I__1541\ : InMux
    port map (
            O => \N__11314\,
            I => \N__11300\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__11311\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__11308\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__1538\ : Odrv4
    port map (
            O => \N__11305\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__11300\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__11291\,
            I => \this_vga_signals.g1_2_cascade_\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__11288\,
            I => \N__11280\
        );

    \I__1534\ : InMux
    port map (
            O => \N__11287\,
            I => \N__11266\
        );

    \I__1533\ : InMux
    port map (
            O => \N__11286\,
            I => \N__11266\
        );

    \I__1532\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11263\
        );

    \I__1531\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11258\
        );

    \I__1530\ : InMux
    port map (
            O => \N__11283\,
            I => \N__11258\
        );

    \I__1529\ : InMux
    port map (
            O => \N__11280\,
            I => \N__11249\
        );

    \I__1528\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11249\
        );

    \I__1527\ : InMux
    port map (
            O => \N__11278\,
            I => \N__11249\
        );

    \I__1526\ : InMux
    port map (
            O => \N__11277\,
            I => \N__11249\
        );

    \I__1525\ : InMux
    port map (
            O => \N__11276\,
            I => \N__11244\
        );

    \I__1524\ : InMux
    port map (
            O => \N__11275\,
            I => \N__11244\
        );

    \I__1523\ : InMux
    port map (
            O => \N__11274\,
            I => \N__11235\
        );

    \I__1522\ : InMux
    port map (
            O => \N__11273\,
            I => \N__11235\
        );

    \I__1521\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11235\
        );

    \I__1520\ : InMux
    port map (
            O => \N__11271\,
            I => \N__11235\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__11266\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__11263\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__11258\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__11249\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__11244\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__11235\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__11222\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_0_cascade_\
        );

    \I__1512\ : InMux
    port map (
            O => \N__11219\,
            I => \N__11216\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__11216\,
            I => \this_vga_signals.g1_1\
        );

    \I__1510\ : InMux
    port map (
            O => \N__11213\,
            I => \N__11210\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__11210\,
            I => \N__11207\
        );

    \I__1508\ : Odrv4
    port map (
            O => \N__11207\,
            I => \this_vga_signals.N_4_i_0_x\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__11204\,
            I => \N__11201\
        );

    \I__1506\ : InMux
    port map (
            O => \N__11201\,
            I => \N__11195\
        );

    \I__1505\ : InMux
    port map (
            O => \N__11200\,
            I => \N__11195\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__11195\,
            I => \N__11190\
        );

    \I__1503\ : InMux
    port map (
            O => \N__11194\,
            I => \N__11185\
        );

    \I__1502\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11185\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__11190\,
            I => \this_vga_signals.N_4_i_0_1\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__11185\,
            I => \this_vga_signals.N_4_i_0_1\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__11180\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_0_1_cascade_\
        );

    \I__1498\ : CascadeMux
    port map (
            O => \N__11177\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\
        );

    \I__1497\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11171\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__11171\,
            I => \this_vga_signals.N_57_i_i_0_0\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__11168\,
            I => \this_vga_signals.g0_1_0_cascade_\
        );

    \I__1494\ : InMux
    port map (
            O => \N__11165\,
            I => \N__11162\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__11162\,
            I => \this_vga_signals.N_5_0_0_1\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__11159\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_3_0_0_0_cascade_\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__11156\,
            I => \N__11153\
        );

    \I__1490\ : InMux
    port map (
            O => \N__11153\,
            I => \N__11150\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__11150\,
            I => \N__11147\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__11147\,
            I => this_vga_signals_address_0_i_7
        );

    \I__1487\ : InMux
    port map (
            O => \N__11144\,
            I => \N__11141\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__11141\,
            I => \this_vga_signals.N_6_0_0\
        );

    \I__1485\ : InMux
    port map (
            O => \N__11138\,
            I => \N__11135\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__11135\,
            I => \this_vga_signals.mult1_un75_sum_c2_0_0_0_1\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__11132\,
            I => \N__11129\
        );

    \I__1482\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11126\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__11126\,
            I => \this_vga_signals.g3_3_0\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__11123\,
            I => \N__11120\
        );

    \I__1479\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11117\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__11117\,
            I => \this_vga_signals.g3_1_0\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__11114\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i_cascade_\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__11111\,
            I => \N__11108\
        );

    \I__1475\ : CascadeBuf
    port map (
            O => \N__11108\,
            I => \N__11105\
        );

    \I__1474\ : CascadeMux
    port map (
            O => \N__11105\,
            I => \N__11102\
        );

    \I__1473\ : CascadeBuf
    port map (
            O => \N__11102\,
            I => \N__11099\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__11099\,
            I => \N__11096\
        );

    \I__1471\ : CascadeBuf
    port map (
            O => \N__11096\,
            I => \N__11093\
        );

    \I__1470\ : CascadeMux
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__1469\ : CascadeBuf
    port map (
            O => \N__11090\,
            I => \N__11087\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__11087\,
            I => \N__11084\
        );

    \I__1467\ : CascadeBuf
    port map (
            O => \N__11084\,
            I => \N__11081\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__11081\,
            I => \N__11078\
        );

    \I__1465\ : CascadeBuf
    port map (
            O => \N__11078\,
            I => \N__11075\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__11075\,
            I => \N__11072\
        );

    \I__1463\ : CascadeBuf
    port map (
            O => \N__11072\,
            I => \N__11069\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__11069\,
            I => \N__11066\
        );

    \I__1461\ : CascadeBuf
    port map (
            O => \N__11066\,
            I => \N__11063\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__11063\,
            I => \N__11060\
        );

    \I__1459\ : CascadeBuf
    port map (
            O => \N__11060\,
            I => \N__11057\
        );

    \I__1458\ : CascadeMux
    port map (
            O => \N__11057\,
            I => \N__11054\
        );

    \I__1457\ : CascadeBuf
    port map (
            O => \N__11054\,
            I => \N__11051\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__11051\,
            I => \N__11048\
        );

    \I__1455\ : CascadeBuf
    port map (
            O => \N__11048\,
            I => \N__11045\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__11045\,
            I => \N__11042\
        );

    \I__1453\ : CascadeBuf
    port map (
            O => \N__11042\,
            I => \N__11039\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__11039\,
            I => \N__11036\
        );

    \I__1451\ : CascadeBuf
    port map (
            O => \N__11036\,
            I => \N__11033\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__11033\,
            I => \N__11030\
        );

    \I__1449\ : CascadeBuf
    port map (
            O => \N__11030\,
            I => \N__11027\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__11027\,
            I => \N__11024\
        );

    \I__1447\ : CascadeBuf
    port map (
            O => \N__11024\,
            I => \N__11021\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__11021\,
            I => \N__11018\
        );

    \I__1445\ : InMux
    port map (
            O => \N__11018\,
            I => \N__11014\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__11017\,
            I => \N__11011\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__11014\,
            I => \N__11008\
        );

    \I__1442\ : InMux
    port map (
            O => \N__11011\,
            I => \N__11005\
        );

    \I__1441\ : Span4Mux_v
    port map (
            O => \N__11008\,
            I => \N__11002\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__11005\,
            I => \N__10999\
        );

    \I__1439\ : Span4Mux_h
    port map (
            O => \N__11002\,
            I => \N__10996\
        );

    \I__1438\ : Sp12to4
    port map (
            O => \N__10999\,
            I => \N__10991\
        );

    \I__1437\ : Sp12to4
    port map (
            O => \N__10996\,
            I => \N__10988\
        );

    \I__1436\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10985\
        );

    \I__1435\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10982\
        );

    \I__1434\ : Span12Mux_v
    port map (
            O => \N__10991\,
            I => \N__10977\
        );

    \I__1433\ : Span12Mux_h
    port map (
            O => \N__10988\,
            I => \N__10977\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__10985\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__10982\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__1430\ : Odrv12
    port map (
            O => \N__10977\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__10970\,
            I => \N__10967\
        );

    \I__1428\ : CascadeBuf
    port map (
            O => \N__10967\,
            I => \N__10964\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__10964\,
            I => \N__10961\
        );

    \I__1426\ : CascadeBuf
    port map (
            O => \N__10961\,
            I => \N__10958\
        );

    \I__1425\ : CascadeMux
    port map (
            O => \N__10958\,
            I => \N__10955\
        );

    \I__1424\ : CascadeBuf
    port map (
            O => \N__10955\,
            I => \N__10952\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__10952\,
            I => \N__10949\
        );

    \I__1422\ : CascadeBuf
    port map (
            O => \N__10949\,
            I => \N__10946\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__10946\,
            I => \N__10943\
        );

    \I__1420\ : CascadeBuf
    port map (
            O => \N__10943\,
            I => \N__10940\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__10940\,
            I => \N__10937\
        );

    \I__1418\ : CascadeBuf
    port map (
            O => \N__10937\,
            I => \N__10934\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__10934\,
            I => \N__10931\
        );

    \I__1416\ : CascadeBuf
    port map (
            O => \N__10931\,
            I => \N__10928\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__10928\,
            I => \N__10925\
        );

    \I__1414\ : CascadeBuf
    port map (
            O => \N__10925\,
            I => \N__10922\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__10922\,
            I => \N__10919\
        );

    \I__1412\ : CascadeBuf
    port map (
            O => \N__10919\,
            I => \N__10916\
        );

    \I__1411\ : CascadeMux
    port map (
            O => \N__10916\,
            I => \N__10913\
        );

    \I__1410\ : CascadeBuf
    port map (
            O => \N__10913\,
            I => \N__10910\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__10910\,
            I => \N__10907\
        );

    \I__1408\ : CascadeBuf
    port map (
            O => \N__10907\,
            I => \N__10904\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__10904\,
            I => \N__10901\
        );

    \I__1406\ : CascadeBuf
    port map (
            O => \N__10901\,
            I => \N__10898\
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__10898\,
            I => \N__10895\
        );

    \I__1404\ : CascadeBuf
    port map (
            O => \N__10895\,
            I => \N__10892\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__10892\,
            I => \N__10889\
        );

    \I__1402\ : CascadeBuf
    port map (
            O => \N__10889\,
            I => \N__10886\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__10886\,
            I => \N__10883\
        );

    \I__1400\ : CascadeBuf
    port map (
            O => \N__10883\,
            I => \N__10879\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__10882\,
            I => \N__10876\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__10879\,
            I => \N__10873\
        );

    \I__1397\ : InMux
    port map (
            O => \N__10876\,
            I => \N__10870\
        );

    \I__1396\ : InMux
    port map (
            O => \N__10873\,
            I => \N__10867\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__10870\,
            I => \N__10864\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__10867\,
            I => \N__10861\
        );

    \I__1393\ : Sp12to4
    port map (
            O => \N__10864\,
            I => \N__10856\
        );

    \I__1392\ : Span12Mux_s11_h
    port map (
            O => \N__10861\,
            I => \N__10853\
        );

    \I__1391\ : InMux
    port map (
            O => \N__10860\,
            I => \N__10850\
        );

    \I__1390\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10847\
        );

    \I__1389\ : Span12Mux_v
    port map (
            O => \N__10856\,
            I => \N__10842\
        );

    \I__1388\ : Span12Mux_h
    port map (
            O => \N__10853\,
            I => \N__10842\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__10850\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__10847\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__1385\ : Odrv12
    port map (
            O => \N__10842\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__10835\,
            I => \N__10832\
        );

    \I__1383\ : CascadeBuf
    port map (
            O => \N__10832\,
            I => \N__10829\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__10829\,
            I => \N__10826\
        );

    \I__1381\ : CascadeBuf
    port map (
            O => \N__10826\,
            I => \N__10823\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__10823\,
            I => \N__10820\
        );

    \I__1379\ : CascadeBuf
    port map (
            O => \N__10820\,
            I => \N__10817\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__10817\,
            I => \N__10814\
        );

    \I__1377\ : CascadeBuf
    port map (
            O => \N__10814\,
            I => \N__10811\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__10811\,
            I => \N__10808\
        );

    \I__1375\ : CascadeBuf
    port map (
            O => \N__10808\,
            I => \N__10805\
        );

    \I__1374\ : CascadeMux
    port map (
            O => \N__10805\,
            I => \N__10802\
        );

    \I__1373\ : CascadeBuf
    port map (
            O => \N__10802\,
            I => \N__10799\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__10799\,
            I => \N__10796\
        );

    \I__1371\ : CascadeBuf
    port map (
            O => \N__10796\,
            I => \N__10793\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__10793\,
            I => \N__10790\
        );

    \I__1369\ : CascadeBuf
    port map (
            O => \N__10790\,
            I => \N__10787\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__10787\,
            I => \N__10784\
        );

    \I__1367\ : CascadeBuf
    port map (
            O => \N__10784\,
            I => \N__10781\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__10781\,
            I => \N__10778\
        );

    \I__1365\ : CascadeBuf
    port map (
            O => \N__10778\,
            I => \N__10775\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__10775\,
            I => \N__10772\
        );

    \I__1363\ : CascadeBuf
    port map (
            O => \N__10772\,
            I => \N__10769\
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__10769\,
            I => \N__10766\
        );

    \I__1361\ : CascadeBuf
    port map (
            O => \N__10766\,
            I => \N__10763\
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__10763\,
            I => \N__10760\
        );

    \I__1359\ : CascadeBuf
    port map (
            O => \N__10760\,
            I => \N__10757\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__10757\,
            I => \N__10754\
        );

    \I__1357\ : CascadeBuf
    port map (
            O => \N__10754\,
            I => \N__10751\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__10751\,
            I => \N__10748\
        );

    \I__1355\ : CascadeBuf
    port map (
            O => \N__10748\,
            I => \N__10745\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__10745\,
            I => \N__10742\
        );

    \I__1353\ : InMux
    port map (
            O => \N__10742\,
            I => \N__10739\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__10739\,
            I => \N__10735\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__10738\,
            I => \N__10732\
        );

    \I__1350\ : Span4Mux_s3_v
    port map (
            O => \N__10735\,
            I => \N__10729\
        );

    \I__1349\ : InMux
    port map (
            O => \N__10732\,
            I => \N__10725\
        );

    \I__1348\ : Span4Mux_h
    port map (
            O => \N__10729\,
            I => \N__10722\
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__10728\,
            I => \N__10718\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__10725\,
            I => \N__10715\
        );

    \I__1345\ : Sp12to4
    port map (
            O => \N__10722\,
            I => \N__10712\
        );

    \I__1344\ : InMux
    port map (
            O => \N__10721\,
            I => \N__10709\
        );

    \I__1343\ : InMux
    port map (
            O => \N__10718\,
            I => \N__10706\
        );

    \I__1342\ : Sp12to4
    port map (
            O => \N__10715\,
            I => \N__10703\
        );

    \I__1341\ : Span12Mux_h
    port map (
            O => \N__10712\,
            I => \N__10700\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__10709\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__10706\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__1338\ : Odrv12
    port map (
            O => \N__10703\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__1337\ : Odrv12
    port map (
            O => \N__10700\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__1336\ : InMux
    port map (
            O => \N__10691\,
            I => \N__10688\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__10688\,
            I => \this_ppu.un1_M_state_d8_5_0\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__10685\,
            I => \M_this_sprites_ram_read_data_0_cascade_\
        );

    \I__1333\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10679\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__10679\,
            I => \N__10676\
        );

    \I__1331\ : Span12Mux_v
    port map (
            O => \N__10676\,
            I => \N__10673\
        );

    \I__1330\ : Odrv12
    port map (
            O => \N__10673\,
            I => \M_this_vram_write_data_0\
        );

    \I__1329\ : InMux
    port map (
            O => \N__10670\,
            I => \N__10667\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__10667\,
            I => \N__10664\
        );

    \I__1327\ : Span12Mux_h
    port map (
            O => \N__10664\,
            I => \N__10661\
        );

    \I__1326\ : Odrv12
    port map (
            O => \N__10661\,
            I => port_clk_c
        );

    \I__1325\ : InMux
    port map (
            O => \N__10658\,
            I => \N__10655\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__10655\,
            I => \N__10652\
        );

    \I__1323\ : Span4Mux_v
    port map (
            O => \N__10652\,
            I => \N__10649\
        );

    \I__1322\ : Odrv4
    port map (
            O => \N__10649\,
            I => \this_vga_signals.vsync_1_0_a2_6_a2_1_0\
        );

    \I__1321\ : IoInMux
    port map (
            O => \N__10646\,
            I => \N__10643\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__10643\,
            I => \N__10640\
        );

    \I__1319\ : Span4Mux_s0_v
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__1318\ : Sp12to4
    port map (
            O => \N__10637\,
            I => \N__10634\
        );

    \I__1317\ : Span12Mux_s7_h
    port map (
            O => \N__10634\,
            I => \N__10631\
        );

    \I__1316\ : Span12Mux_v
    port map (
            O => \N__10631\,
            I => \N__10628\
        );

    \I__1315\ : Odrv12
    port map (
            O => \N__10628\,
            I => this_vga_signals_vsync_1_i
        );

    \I__1314\ : InMux
    port map (
            O => \N__10625\,
            I => \N__10622\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__10622\,
            I => \this_delay_clk.M_pipe_qZ0Z_0\
        );

    \I__1312\ : InMux
    port map (
            O => \N__10619\,
            I => \N__10616\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__10616\,
            I => \this_delay_clk.M_pipe_qZ0Z_1\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__10613\,
            I => \this_vga_signals.g0_16_x0_cascade_\
        );

    \I__1309\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10607\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__10607\,
            I => \this_vga_signals.g3_0\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__10604\,
            I => \this_vga_signals_un4_lcounter_if_i1_mux_cascade_\
        );

    \I__1306\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10595\
        );

    \I__1305\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10592\
        );

    \I__1304\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10587\
        );

    \I__1303\ : InMux
    port map (
            O => \N__10598\,
            I => \N__10587\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__10595\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__10592\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__10587\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0
        );

    \I__1299\ : CascadeMux
    port map (
            O => \N__10580\,
            I => \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_cascade_\
        );

    \I__1298\ : InMux
    port map (
            O => \N__10577\,
            I => \N__10573\
        );

    \I__1297\ : InMux
    port map (
            O => \N__10576\,
            I => \N__10570\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__10573\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_1
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__10570\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_1
        );

    \I__1294\ : InMux
    port map (
            O => \N__10565\,
            I => \N__10562\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__10562\,
            I => \this_ppu.M_m7Z0Z_1\
        );

    \I__1292\ : InMux
    port map (
            O => \N__10559\,
            I => \N__10556\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__10556\,
            I => \N__10553\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__10553\,
            I => \this_ppu.M_m12_0_o2_381_10Z0Z_1\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__10550\,
            I => \this_ppu.M_N_11_mux_cascade_\
        );

    \I__1288\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10543\
        );

    \I__1287\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10540\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__10543\,
            I => \this_ppu.M_m12_0_o2_381_10\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__10540\,
            I => \this_ppu.M_m12_0_o2_381_10\
        );

    \I__1284\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10531\
        );

    \I__1283\ : InMux
    port map (
            O => \N__10534\,
            I => \N__10528\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__10531\,
            I => this_vga_signals_un4_lcounter_if_i1_mux
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__10528\,
            I => this_vga_signals_un4_lcounter_if_i1_mux
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__10523\,
            I => \N__10520\
        );

    \I__1279\ : InMux
    port map (
            O => \N__10520\,
            I => \N__10515\
        );

    \I__1278\ : InMux
    port map (
            O => \N__10519\,
            I => \N__10512\
        );

    \I__1277\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10509\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__10515\,
            I => \N__10504\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__10512\,
            I => \N__10504\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__10509\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1
        );

    \I__1273\ : Odrv4
    port map (
            O => \N__10504\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1
        );

    \I__1272\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10496\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__10496\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_1
        );

    \I__1270\ : InMux
    port map (
            O => \N__10493\,
            I => \N__10486\
        );

    \I__1269\ : InMux
    port map (
            O => \N__10492\,
            I => \N__10486\
        );

    \I__1268\ : InMux
    port map (
            O => \N__10491\,
            I => \N__10483\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__10486\,
            I => \this_vga_signals_un4_lcounter_if_N_7_i_i\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__10483\,
            I => \this_vga_signals_un4_lcounter_if_N_7_i_i\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__10478\,
            I => \N__10475\
        );

    \I__1264\ : CascadeBuf
    port map (
            O => \N__10475\,
            I => \N__10472\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__10472\,
            I => \N__10469\
        );

    \I__1262\ : CascadeBuf
    port map (
            O => \N__10469\,
            I => \N__10466\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__10466\,
            I => \N__10463\
        );

    \I__1260\ : CascadeBuf
    port map (
            O => \N__10463\,
            I => \N__10460\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__10460\,
            I => \N__10457\
        );

    \I__1258\ : CascadeBuf
    port map (
            O => \N__10457\,
            I => \N__10454\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__10454\,
            I => \N__10451\
        );

    \I__1256\ : CascadeBuf
    port map (
            O => \N__10451\,
            I => \N__10448\
        );

    \I__1255\ : CascadeMux
    port map (
            O => \N__10448\,
            I => \N__10445\
        );

    \I__1254\ : CascadeBuf
    port map (
            O => \N__10445\,
            I => \N__10442\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__10442\,
            I => \N__10439\
        );

    \I__1252\ : CascadeBuf
    port map (
            O => \N__10439\,
            I => \N__10436\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__10436\,
            I => \N__10433\
        );

    \I__1250\ : CascadeBuf
    port map (
            O => \N__10433\,
            I => \N__10430\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__10430\,
            I => \N__10427\
        );

    \I__1248\ : CascadeBuf
    port map (
            O => \N__10427\,
            I => \N__10424\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__10424\,
            I => \N__10421\
        );

    \I__1246\ : CascadeBuf
    port map (
            O => \N__10421\,
            I => \N__10418\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__10418\,
            I => \N__10415\
        );

    \I__1244\ : CascadeBuf
    port map (
            O => \N__10415\,
            I => \N__10412\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__10412\,
            I => \N__10409\
        );

    \I__1242\ : CascadeBuf
    port map (
            O => \N__10409\,
            I => \N__10406\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__10406\,
            I => \N__10403\
        );

    \I__1240\ : CascadeBuf
    port map (
            O => \N__10403\,
            I => \N__10400\
        );

    \I__1239\ : CascadeMux
    port map (
            O => \N__10400\,
            I => \N__10397\
        );

    \I__1238\ : CascadeBuf
    port map (
            O => \N__10397\,
            I => \N__10394\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__10394\,
            I => \N__10391\
        );

    \I__1236\ : CascadeBuf
    port map (
            O => \N__10391\,
            I => \N__10388\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__1234\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__10382\,
            I => \N__10378\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__10381\,
            I => \N__10375\
        );

    \I__1231\ : Span4Mux_h
    port map (
            O => \N__10378\,
            I => \N__10372\
        );

    \I__1230\ : InMux
    port map (
            O => \N__10375\,
            I => \N__10369\
        );

    \I__1229\ : Span4Mux_h
    port map (
            O => \N__10372\,
            I => \N__10366\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__10369\,
            I => \N__10361\
        );

    \I__1227\ : Sp12to4
    port map (
            O => \N__10366\,
            I => \N__10358\
        );

    \I__1226\ : InMux
    port map (
            O => \N__10365\,
            I => \N__10355\
        );

    \I__1225\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10352\
        );

    \I__1224\ : Span12Mux_v
    port map (
            O => \N__10361\,
            I => \N__10347\
        );

    \I__1223\ : Span12Mux_v
    port map (
            O => \N__10358\,
            I => \N__10347\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__10355\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__10352\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__1220\ : Odrv12
    port map (
            O => \N__10347\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__1218\ : CascadeBuf
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__10334\,
            I => \N__10331\
        );

    \I__1216\ : CascadeBuf
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__10328\,
            I => \N__10325\
        );

    \I__1214\ : CascadeBuf
    port map (
            O => \N__10325\,
            I => \N__10322\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__10322\,
            I => \N__10319\
        );

    \I__1212\ : CascadeBuf
    port map (
            O => \N__10319\,
            I => \N__10316\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__10316\,
            I => \N__10313\
        );

    \I__1210\ : CascadeBuf
    port map (
            O => \N__10313\,
            I => \N__10310\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__10310\,
            I => \N__10307\
        );

    \I__1208\ : CascadeBuf
    port map (
            O => \N__10307\,
            I => \N__10304\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__10304\,
            I => \N__10301\
        );

    \I__1206\ : CascadeBuf
    port map (
            O => \N__10301\,
            I => \N__10298\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__10298\,
            I => \N__10295\
        );

    \I__1204\ : CascadeBuf
    port map (
            O => \N__10295\,
            I => \N__10292\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__10292\,
            I => \N__10289\
        );

    \I__1202\ : CascadeBuf
    port map (
            O => \N__10289\,
            I => \N__10286\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__10286\,
            I => \N__10283\
        );

    \I__1200\ : CascadeBuf
    port map (
            O => \N__10283\,
            I => \N__10280\
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__10280\,
            I => \N__10277\
        );

    \I__1198\ : CascadeBuf
    port map (
            O => \N__10277\,
            I => \N__10274\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__10274\,
            I => \N__10271\
        );

    \I__1196\ : CascadeBuf
    port map (
            O => \N__10271\,
            I => \N__10268\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__10268\,
            I => \N__10265\
        );

    \I__1194\ : CascadeBuf
    port map (
            O => \N__10265\,
            I => \N__10262\
        );

    \I__1193\ : CascadeMux
    port map (
            O => \N__10262\,
            I => \N__10259\
        );

    \I__1192\ : CascadeBuf
    port map (
            O => \N__10259\,
            I => \N__10256\
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__10256\,
            I => \N__10253\
        );

    \I__1190\ : CascadeBuf
    port map (
            O => \N__10253\,
            I => \N__10250\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__10250\,
            I => \N__10247\
        );

    \I__1188\ : InMux
    port map (
            O => \N__10247\,
            I => \N__10243\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__10246\,
            I => \N__10240\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__10243\,
            I => \N__10237\
        );

    \I__1185\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10234\
        );

    \I__1184\ : Span4Mux_s2_v
    port map (
            O => \N__10237\,
            I => \N__10231\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__10234\,
            I => \N__10228\
        );

    \I__1182\ : Span4Mux_h
    port map (
            O => \N__10231\,
            I => \N__10225\
        );

    \I__1181\ : Span4Mux_v
    port map (
            O => \N__10228\,
            I => \N__10220\
        );

    \I__1180\ : Sp12to4
    port map (
            O => \N__10225\,
            I => \N__10217\
        );

    \I__1179\ : InMux
    port map (
            O => \N__10224\,
            I => \N__10214\
        );

    \I__1178\ : InMux
    port map (
            O => \N__10223\,
            I => \N__10211\
        );

    \I__1177\ : Span4Mux_v
    port map (
            O => \N__10220\,
            I => \N__10208\
        );

    \I__1176\ : Span12Mux_v
    port map (
            O => \N__10217\,
            I => \N__10205\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__10214\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__10211\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__1173\ : Odrv4
    port map (
            O => \N__10208\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__1172\ : Odrv12
    port map (
            O => \N__10205\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__10196\,
            I => \N__10193\
        );

    \I__1170\ : CascadeBuf
    port map (
            O => \N__10193\,
            I => \N__10190\
        );

    \I__1169\ : CascadeMux
    port map (
            O => \N__10190\,
            I => \N__10187\
        );

    \I__1168\ : CascadeBuf
    port map (
            O => \N__10187\,
            I => \N__10184\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__10184\,
            I => \N__10181\
        );

    \I__1166\ : CascadeBuf
    port map (
            O => \N__10181\,
            I => \N__10178\
        );

    \I__1165\ : CascadeMux
    port map (
            O => \N__10178\,
            I => \N__10175\
        );

    \I__1164\ : CascadeBuf
    port map (
            O => \N__10175\,
            I => \N__10172\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__10172\,
            I => \N__10169\
        );

    \I__1162\ : CascadeBuf
    port map (
            O => \N__10169\,
            I => \N__10166\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__10166\,
            I => \N__10163\
        );

    \I__1160\ : CascadeBuf
    port map (
            O => \N__10163\,
            I => \N__10160\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__10160\,
            I => \N__10157\
        );

    \I__1158\ : CascadeBuf
    port map (
            O => \N__10157\,
            I => \N__10154\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__10154\,
            I => \N__10151\
        );

    \I__1156\ : CascadeBuf
    port map (
            O => \N__10151\,
            I => \N__10148\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__10148\,
            I => \N__10145\
        );

    \I__1154\ : CascadeBuf
    port map (
            O => \N__10145\,
            I => \N__10142\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__10142\,
            I => \N__10139\
        );

    \I__1152\ : CascadeBuf
    port map (
            O => \N__10139\,
            I => \N__10136\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__10136\,
            I => \N__10133\
        );

    \I__1150\ : CascadeBuf
    port map (
            O => \N__10133\,
            I => \N__10130\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__10130\,
            I => \N__10127\
        );

    \I__1148\ : CascadeBuf
    port map (
            O => \N__10127\,
            I => \N__10124\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__10124\,
            I => \N__10121\
        );

    \I__1146\ : CascadeBuf
    port map (
            O => \N__10121\,
            I => \N__10118\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__10118\,
            I => \N__10115\
        );

    \I__1144\ : CascadeBuf
    port map (
            O => \N__10115\,
            I => \N__10112\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__10112\,
            I => \N__10109\
        );

    \I__1142\ : CascadeBuf
    port map (
            O => \N__10109\,
            I => \N__10106\
        );

    \I__1141\ : CascadeMux
    port map (
            O => \N__10106\,
            I => \N__10103\
        );

    \I__1140\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10100\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__10100\,
            I => \N__10096\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__10099\,
            I => \N__10093\
        );

    \I__1137\ : Span4Mux_s2_v
    port map (
            O => \N__10096\,
            I => \N__10090\
        );

    \I__1136\ : InMux
    port map (
            O => \N__10093\,
            I => \N__10087\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__10090\,
            I => \N__10084\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__10087\,
            I => \N__10080\
        );

    \I__1133\ : Span4Mux_v
    port map (
            O => \N__10084\,
            I => \N__10077\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__10083\,
            I => \N__10074\
        );

    \I__1131\ : Span4Mux_v
    port map (
            O => \N__10080\,
            I => \N__10070\
        );

    \I__1130\ : Sp12to4
    port map (
            O => \N__10077\,
            I => \N__10067\
        );

    \I__1129\ : InMux
    port map (
            O => \N__10074\,
            I => \N__10064\
        );

    \I__1128\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10061\
        );

    \I__1127\ : Sp12to4
    port map (
            O => \N__10070\,
            I => \N__10056\
        );

    \I__1126\ : Span12Mux_h
    port map (
            O => \N__10067\,
            I => \N__10056\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__10064\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__10061\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__1123\ : Odrv12
    port map (
            O => \N__10056\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__10049\,
            I => \N__10046\
        );

    \I__1121\ : CascadeBuf
    port map (
            O => \N__10046\,
            I => \N__10043\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__10043\,
            I => \N__10040\
        );

    \I__1119\ : CascadeBuf
    port map (
            O => \N__10040\,
            I => \N__10037\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__10037\,
            I => \N__10034\
        );

    \I__1117\ : CascadeBuf
    port map (
            O => \N__10034\,
            I => \N__10031\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__10031\,
            I => \N__10028\
        );

    \I__1115\ : CascadeBuf
    port map (
            O => \N__10028\,
            I => \N__10025\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__10025\,
            I => \N__10022\
        );

    \I__1113\ : CascadeBuf
    port map (
            O => \N__10022\,
            I => \N__10019\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__10019\,
            I => \N__10016\
        );

    \I__1111\ : CascadeBuf
    port map (
            O => \N__10016\,
            I => \N__10013\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__10013\,
            I => \N__10010\
        );

    \I__1109\ : CascadeBuf
    port map (
            O => \N__10010\,
            I => \N__10007\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__10007\,
            I => \N__10004\
        );

    \I__1107\ : CascadeBuf
    port map (
            O => \N__10004\,
            I => \N__10001\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__10001\,
            I => \N__9998\
        );

    \I__1105\ : CascadeBuf
    port map (
            O => \N__9998\,
            I => \N__9995\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__9995\,
            I => \N__9992\
        );

    \I__1103\ : CascadeBuf
    port map (
            O => \N__9992\,
            I => \N__9989\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__1101\ : CascadeBuf
    port map (
            O => \N__9986\,
            I => \N__9983\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__9983\,
            I => \N__9980\
        );

    \I__1099\ : CascadeBuf
    port map (
            O => \N__9980\,
            I => \N__9977\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__9977\,
            I => \N__9974\
        );

    \I__1097\ : CascadeBuf
    port map (
            O => \N__9974\,
            I => \N__9971\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__9971\,
            I => \N__9968\
        );

    \I__1095\ : CascadeBuf
    port map (
            O => \N__9968\,
            I => \N__9965\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__9965\,
            I => \N__9962\
        );

    \I__1093\ : CascadeBuf
    port map (
            O => \N__9962\,
            I => \N__9959\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__9959\,
            I => \N__9956\
        );

    \I__1091\ : InMux
    port map (
            O => \N__9956\,
            I => \N__9953\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__9953\,
            I => \N__9949\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__9952\,
            I => \N__9946\
        );

    \I__1088\ : Span4Mux_s2_v
    port map (
            O => \N__9949\,
            I => \N__9943\
        );

    \I__1087\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9940\
        );

    \I__1086\ : Span4Mux_h
    port map (
            O => \N__9943\,
            I => \N__9937\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__9940\,
            I => \N__9932\
        );

    \I__1084\ : Sp12to4
    port map (
            O => \N__9937\,
            I => \N__9929\
        );

    \I__1083\ : InMux
    port map (
            O => \N__9936\,
            I => \N__9926\
        );

    \I__1082\ : InMux
    port map (
            O => \N__9935\,
            I => \N__9923\
        );

    \I__1081\ : Span12Mux_s8_h
    port map (
            O => \N__9932\,
            I => \N__9920\
        );

    \I__1080\ : Span12Mux_h
    port map (
            O => \N__9929\,
            I => \N__9917\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__9926\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__9923\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__1077\ : Odrv12
    port map (
            O => \N__9920\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__1076\ : Odrv12
    port map (
            O => \N__9917\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__9908\,
            I => \this_ppu.un1_M_state_d8_4_0_cascade_\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__9902\,
            I => \this_ppu.M_N_3_mux_0_0\
        );

    \I__1072\ : InMux
    port map (
            O => \N__9899\,
            I => \N__9896\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__9896\,
            I => \N__9891\
        );

    \I__1070\ : InMux
    port map (
            O => \N__9895\,
            I => \N__9888\
        );

    \I__1069\ : InMux
    port map (
            O => \N__9894\,
            I => \N__9885\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__9891\,
            I => \this_vga_signals.CO1_5_0\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__9888\,
            I => \this_vga_signals.CO1_5_0\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__9885\,
            I => \this_vga_signals.CO1_5_0\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__9878\,
            I => \this_vga_signals.mult1_un40_sum0_2_cascade_\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__9875\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_2_cascade_\
        );

    \I__1063\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9869\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__9869\,
            I => \N__9865\
        );

    \I__1061\ : InMux
    port map (
            O => \N__9868\,
            I => \N__9862\
        );

    \I__1060\ : Span4Mux_h
    port map (
            O => \N__9865\,
            I => \N__9859\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__9862\,
            I => \N__9856\
        );

    \I__1058\ : Odrv4
    port map (
            O => \N__9859\,
            I => \this_vga_signals.N_196_0\
        );

    \I__1057\ : Odrv4
    port map (
            O => \N__9856\,
            I => \this_vga_signals.N_196_0\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__9851\,
            I => \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0_cascade_\
        );

    \I__1055\ : InMux
    port map (
            O => \N__9848\,
            I => \N__9842\
        );

    \I__1054\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9842\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__9842\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un54_sum_axb1
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__9839\,
            I => \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un54_sum_axb1_cascade_\
        );

    \I__1051\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9832\
        );

    \I__1050\ : InMux
    port map (
            O => \N__9835\,
            I => \N__9829\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__9832\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_c3_0
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__9829\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_c3_0
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__9824\,
            I => \this_vga_signals.mult1_un40_sum_0_c3_0_cascade_\
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__9821\,
            I => \N__9818\
        );

    \I__1045\ : InMux
    port map (
            O => \N__9818\,
            I => \N__9814\
        );

    \I__1044\ : InMux
    port map (
            O => \N__9817\,
            I => \N__9811\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__9814\,
            I => \N__9808\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__9811\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__9808\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__1040\ : InMux
    port map (
            O => \N__9803\,
            I => \N__9799\
        );

    \I__1039\ : InMux
    port map (
            O => \N__9802\,
            I => \N__9796\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__9799\,
            I => \N__9793\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__9796\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__1036\ : Odrv4
    port map (
            O => \N__9793\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__1035\ : InMux
    port map (
            O => \N__9788\,
            I => \N__9785\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__9785\,
            I => \N__9781\
        );

    \I__1033\ : InMux
    port map (
            O => \N__9784\,
            I => \N__9778\
        );

    \I__1032\ : Odrv4
    port map (
            O => \N__9781\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__9778\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__1030\ : InMux
    port map (
            O => \N__9773\,
            I => \N__9770\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__9770\,
            I => \this_vga_signals.mult1_un40_sum_0_c3_0\
        );

    \I__1028\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9764\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__9764\,
            I => \this_vga_signals.mult1_un40_sum_1_c2_0\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__9761\,
            I => \this_vga_signals.mult1_un40_sum_m_x1_3_cascade_\
        );

    \I__1025\ : InMux
    port map (
            O => \N__9758\,
            I => \N__9755\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__9755\,
            I => \this_vga_signals.mult1_un40_sum_m_x0_3\
        );

    \I__1023\ : InMux
    port map (
            O => \N__9752\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_1\
        );

    \I__1022\ : InMux
    port map (
            O => \N__9749\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_2\
        );

    \I__1021\ : InMux
    port map (
            O => \N__9746\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3\
        );

    \I__1020\ : InMux
    port map (
            O => \N__9743\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4\
        );

    \I__1019\ : InMux
    port map (
            O => \N__9740\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5\
        );

    \I__1018\ : InMux
    port map (
            O => \N__9737\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6\
        );

    \I__1017\ : InMux
    port map (
            O => \N__9734\,
            I => \bfn_10_15_0_\
        );

    \I__1016\ : InMux
    port map (
            O => \N__9731\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__9728\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_1_0_cascade_\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__9725\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\
        );

    \I__1013\ : InMux
    port map (
            O => \N__9722\,
            I => \N__9719\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__9719\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_1_0_0\
        );

    \I__1011\ : InMux
    port map (
            O => \N__9716\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_0\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__9713\,
            I => \this_vga_signals.g0_3_0_a3_2_cascade_\
        );

    \I__1009\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9707\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__9707\,
            I => \this_vga_signals.g2_1\
        );

    \I__1007\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9701\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__9701\,
            I => \N__9698\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__9698\,
            I => \this_vga_signals.g1_0_0_0\
        );

    \I__1004\ : CascadeMux
    port map (
            O => \N__9695\,
            I => \this_vga_signals.N_188_0_cascade_\
        );

    \I__1003\ : CascadeMux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__1002\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9686\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__9686\,
            I => \this_vga_signals.if_m10_0_a4_0_0\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__9683\,
            I => \this_vga_signals.g1_3_0_cascade_\
        );

    \I__999\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9677\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__9677\,
            I => \this_vga_signals.if_m10_0_a4_1_1\
        );

    \I__997\ : InMux
    port map (
            O => \N__9674\,
            I => \N__9671\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__9671\,
            I => \this_vga_signals.if_N_18_0\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__9668\,
            I => \N__9664\
        );

    \I__994\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9661\
        );

    \I__993\ : InMux
    port map (
            O => \N__9664\,
            I => \N__9658\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__9661\,
            I => \this_vga_signals.N_3_1\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__9658\,
            I => \this_vga_signals.N_3_1\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__9653\,
            I => \N__9650\
        );

    \I__989\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9644\
        );

    \I__988\ : InMux
    port map (
            O => \N__9649\,
            I => \N__9644\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__9644\,
            I => \this_vga_signals.m6_2\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__9641\,
            I => \N__9638\
        );

    \I__985\ : InMux
    port map (
            O => \N__9638\,
            I => \N__9635\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__9635\,
            I => \N__9632\
        );

    \I__983\ : Odrv4
    port map (
            O => \N__9632\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_0_0\
        );

    \I__982\ : InMux
    port map (
            O => \N__9629\,
            I => \N__9626\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__9626\,
            I => \N__9621\
        );

    \I__980\ : InMux
    port map (
            O => \N__9625\,
            I => \N__9618\
        );

    \I__979\ : InMux
    port map (
            O => \N__9624\,
            I => \N__9615\
        );

    \I__978\ : Odrv4
    port map (
            O => \N__9621\,
            I => \this_vga_signals.if_i3_mux_0_0\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__9618\,
            I => \this_vga_signals.if_i3_mux_0_0\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__9615\,
            I => \this_vga_signals.if_i3_mux_0_0\
        );

    \I__975\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9605\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__9605\,
            I => \this_vga_signals.M_vcounter_q_RNI820378Z0Z_2\
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__9602\,
            I => \this_vga_signals.N_3_0_cascade_\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__9599\,
            I => \this_vga_signals.g1_cascade_\
        );

    \I__971\ : InMux
    port map (
            O => \N__9596\,
            I => \N__9593\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__9593\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__969\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9587\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__9587\,
            I => \this_vga_signals.M_vcounter_q_RNI820378_0Z0Z_2\
        );

    \I__967\ : InMux
    port map (
            O => \N__9584\,
            I => \N__9580\
        );

    \I__966\ : InMux
    port map (
            O => \N__9583\,
            I => \N__9577\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__9580\,
            I => \this_vga_signals.N_9_0_0\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__9577\,
            I => \this_vga_signals.N_9_0_0\
        );

    \I__963\ : CascadeMux
    port map (
            O => \N__9572\,
            I => \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3Z0Z_5_cascade_\
        );

    \I__962\ : InMux
    port map (
            O => \N__9569\,
            I => \N__9566\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__9566\,
            I => \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_0Z0Z_5\
        );

    \I__960\ : InMux
    port map (
            O => \N__9563\,
            I => \N__9560\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__9560\,
            I => \N__9557\
        );

    \I__958\ : Odrv4
    port map (
            O => \N__9557\,
            I => \this_vga_signals.N_5\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__9554\,
            I => \this_vga_signals.g0_0_x2_0_0_a3_3_cascade_\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__9551\,
            I => \this_vga_signals.N_9_i_0_0_cascade_\
        );

    \I__955\ : InMux
    port map (
            O => \N__9548\,
            I => \N__9545\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9545\,
            I => \this_vga_signals.N_9_i_0_0\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__9542\,
            I => \this_vga_signals.g0_2_x0_cascade_\
        );

    \I__952\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9536\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__9536\,
            I => \this_vga_signals.g0_2_x1\
        );

    \I__950\ : InMux
    port map (
            O => \N__9533\,
            I => \this_ppu.un1_M_current_q_cry_0\
        );

    \I__949\ : InMux
    port map (
            O => \N__9530\,
            I => \this_ppu.un1_M_current_q_cry_1\
        );

    \I__948\ : InMux
    port map (
            O => \N__9527\,
            I => \this_ppu.un1_M_current_q_cry_2\
        );

    \I__947\ : InMux
    port map (
            O => \N__9524\,
            I => \this_ppu.un1_M_current_q_cry_3\
        );

    \I__946\ : InMux
    port map (
            O => \N__9521\,
            I => \this_ppu.un1_M_current_q_cry_4\
        );

    \I__945\ : InMux
    port map (
            O => \N__9518\,
            I => \this_ppu.un1_M_current_q_cry_5\
        );

    \I__944\ : SRMux
    port map (
            O => \N__9515\,
            I => \N__9512\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__9512\,
            I => \N__9509\
        );

    \I__942\ : Odrv12
    port map (
            O => \N__9509\,
            I => \this_ppu.N_256_1_i\
        );

    \I__941\ : InMux
    port map (
            O => \N__9506\,
            I => \N__9501\
        );

    \I__940\ : InMux
    port map (
            O => \N__9505\,
            I => \N__9496\
        );

    \I__939\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9496\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__9501\,
            I => \this_vga_signals.mult1_un68_sum_axb1_0\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__9496\,
            I => \this_vga_signals.mult1_un68_sum_axb1_0\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__9491\,
            I => \N__9488\
        );

    \I__935\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9485\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__9485\,
            I => \N__9482\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__9482\,
            I => \M_this_vga_signals_address_10\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__9479\,
            I => \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_c3_0_cascade_\
        );

    \I__931\ : InMux
    port map (
            O => \N__9476\,
            I => \N__9470\
        );

    \I__930\ : InMux
    port map (
            O => \N__9475\,
            I => \N__9470\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__9470\,
            I => \this_ppu.N_277\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__9467\,
            I => \this_ppu.M_mZ0Z1_cascade_\
        );

    \I__927\ : IoInMux
    port map (
            O => \N__9464\,
            I => \N__9461\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__9461\,
            I => \N__9458\
        );

    \I__925\ : IoSpan4Mux
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__924\ : IoSpan4Mux
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__923\ : Span4Mux_s3_v
    port map (
            O => \N__9452\,
            I => \N__9449\
        );

    \I__922\ : Sp12to4
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__921\ : Odrv12
    port map (
            O => \N__9446\,
            I => \N_92\
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__9443\,
            I => \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axb1_cascade_\
        );

    \I__919\ : InMux
    port map (
            O => \N__9440\,
            I => \N__9437\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__9437\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_c3_0
        );

    \I__917\ : InMux
    port map (
            O => \N__9434\,
            I => \N__9431\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__9431\,
            I => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axb1
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__9428\,
            I => \this_ppu.M_N_16_1_cascade_\
        );

    \I__914\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9422\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__9422\,
            I => \N__9418\
        );

    \I__912\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9415\
        );

    \I__911\ : Odrv4
    port map (
            O => \N__9418\,
            I => \this_ppu.M_m9_i_x3Z0Z_0\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__9415\,
            I => \this_ppu.M_m9_i_x3Z0Z_0\
        );

    \I__909\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9407\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__9407\,
            I => \this_ppu.M_mZ0Z1\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__9404\,
            I => \this_ppu.M_m1_e_0_1_0_cascade_\
        );

    \I__906\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9398\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__9398\,
            I => \this_ppu.M_m1_e_0_1_1\
        );

    \I__904\ : InMux
    port map (
            O => \N__9395\,
            I => \N__9389\
        );

    \I__903\ : InMux
    port map (
            O => \N__9394\,
            I => \N__9389\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__9389\,
            I => \this_ppu.M_m12_0_x3_out_0\
        );

    \I__901\ : InMux
    port map (
            O => \N__9386\,
            I => \N__9383\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__9383\,
            I => \this_ppu.M_N_16_1\
        );

    \I__899\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9377\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__9377\,
            I => \this_ppu.M_m1_e_0_0\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__9374\,
            I => \this_ppu.M_N_6_0_cascade_\
        );

    \I__896\ : InMux
    port map (
            O => \N__9371\,
            I => \N__9368\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__9368\,
            I => \this_ppu.M_N_13_mux\
        );

    \I__894\ : InMux
    port map (
            O => \N__9365\,
            I => \N__9362\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__9362\,
            I => \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_c_0\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__9359\,
            I => \this_ppu.M_N_15_mux_cascade_\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__9356\,
            I => \this_ppu.M_m12_0_x3_s_0_1Z0Z_0_cascade_\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__9353\,
            I => \this_ppu.M_m12_0_x3_out_0_cascade_\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__9350\,
            I => \this_vga_signals.if_m12_cascade_\
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__9347\,
            I => \N__9344\
        );

    \I__887\ : InMux
    port map (
            O => \N__9344\,
            I => \N__9341\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__9341\,
            I => \this_vga_signals.mult1_un54_sum_cry_1_s\
        );

    \I__885\ : InMux
    port map (
            O => \N__9338\,
            I => \this_vga_signals.mult1_un54_sum_cry_0\
        );

    \I__884\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9332\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__9332\,
            I => \N__9329\
        );

    \I__882\ : Odrv12
    port map (
            O => \N__9329\,
            I => \this_vga_signals.mult1_un47_sum_cry_1_s\
        );

    \I__881\ : InMux
    port map (
            O => \N__9326\,
            I => \N__9323\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__9323\,
            I => \this_vga_signals.mult1_un61_sum_axb_3\
        );

    \I__879\ : InMux
    port map (
            O => \N__9320\,
            I => \this_vga_signals.mult1_un54_sum_cry_1\
        );

    \I__878\ : InMux
    port map (
            O => \N__9317\,
            I => \N__9314\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__9314\,
            I => \N__9311\
        );

    \I__876\ : Odrv4
    port map (
            O => \N__9311\,
            I => \this_vga_signals.mult1_un54_sum_axb_3\
        );

    \I__875\ : InMux
    port map (
            O => \N__9308\,
            I => \this_vga_signals.mult1_un54_sum_cry_2\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__9305\,
            I => \N__9302\
        );

    \I__873\ : InMux
    port map (
            O => \N__9302\,
            I => \N__9295\
        );

    \I__872\ : InMux
    port map (
            O => \N__9301\,
            I => \N__9295\
        );

    \I__871\ : InMux
    port map (
            O => \N__9300\,
            I => \N__9292\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__9295\,
            I => \this_vga_signals.mult1_un54_sum_s_3\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__9292\,
            I => \this_vga_signals.mult1_un54_sum_s_3\
        );

    \I__868\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9284\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__9284\,
            I => \N__9281\
        );

    \I__866\ : Span4Mux_v
    port map (
            O => \N__9281\,
            I => \N__9278\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__9278\,
            I => \this_vga_signals.M_hcounter_q_i_0_5\
        );

    \I__864\ : CascadeMux
    port map (
            O => \N__9275\,
            I => \N__9272\
        );

    \I__863\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9266\
        );

    \I__862\ : InMux
    port map (
            O => \N__9271\,
            I => \N__9266\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__9266\,
            I => \N__9262\
        );

    \I__860\ : InMux
    port map (
            O => \N__9265\,
            I => \N__9259\
        );

    \I__859\ : Odrv12
    port map (
            O => \N__9262\,
            I => \this_vga_signals.mult1_un47_sum_s_3\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__9259\,
            I => \this_vga_signals.mult1_un47_sum_s_3\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__9254\,
            I => \N__9251\
        );

    \I__856\ : InMux
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__9248\,
            I => \this_vga_signals.mult1_un47_sum_i_3\
        );

    \I__854\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9242\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__9242\,
            I => \this_vga_signals.mult1_un40_sum_axb_2\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__851\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9233\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__9233\,
            I => \N__9230\
        );

    \I__849\ : Odrv4
    port map (
            O => \N__9230\,
            I => \this_vga_signals.mult1_un40_sum_axb_1_l_fx\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__9227\,
            I => \N__9224\
        );

    \I__847\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9217\
        );

    \I__846\ : InMux
    port map (
            O => \N__9223\,
            I => \N__9217\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__9222\,
            I => \N__9214\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__9217\,
            I => \N__9211\
        );

    \I__843\ : InMux
    port map (
            O => \N__9214\,
            I => \N__9208\
        );

    \I__842\ : Odrv4
    port map (
            O => \N__9211\,
            I => \this_vga_signals.mult1_un40_sum_cry_2_THRU_CO\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__9208\,
            I => \this_vga_signals.mult1_un40_sum_cry_2_THRU_CO\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__839\ : InMux
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__9197\,
            I => \this_vga_signals.mult1_un40_sum_s_3\
        );

    \I__837\ : InMux
    port map (
            O => \N__9194\,
            I => \this_vga_signals.mult1_un61_sum_cry_0\
        );

    \I__836\ : InMux
    port map (
            O => \N__9191\,
            I => \this_vga_signals.mult1_un61_sum_cry_1\
        );

    \I__835\ : InMux
    port map (
            O => \N__9188\,
            I => \this_vga_signals.mult1_un61_sum_cry_2\
        );

    \I__834\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9181\
        );

    \I__833\ : InMux
    port map (
            O => \N__9184\,
            I => \N__9178\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__9181\,
            I => \N__9172\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__9178\,
            I => \N__9172\
        );

    \I__830\ : InMux
    port map (
            O => \N__9177\,
            I => \N__9169\
        );

    \I__829\ : Odrv4
    port map (
            O => \N__9172\,
            I => \this_vga_signals.N_70_0\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__9169\,
            I => \this_vga_signals.N_70_0\
        );

    \I__827\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9161\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__9161\,
            I => \this_vga_signals.mult1_un54_sum_i_3\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__9158\,
            I => \N_70_cascade_\
        );

    \I__824\ : InMux
    port map (
            O => \N__9155\,
            I => \N__9152\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__9152\,
            I => \this_vga_signals.mult1_un40_sum_cry_1_THRU_CO\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__9149\,
            I => \N__9146\
        );

    \I__821\ : InMux
    port map (
            O => \N__9146\,
            I => \N__9141\
        );

    \I__820\ : InMux
    port map (
            O => \N__9145\,
            I => \N__9136\
        );

    \I__819\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9136\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__9141\,
            I => \G_501\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__9136\,
            I => \G_501\
        );

    \I__816\ : InMux
    port map (
            O => \N__9131\,
            I => \N__9126\
        );

    \I__815\ : InMux
    port map (
            O => \N__9130\,
            I => \N__9121\
        );

    \I__814\ : InMux
    port map (
            O => \N__9129\,
            I => \N__9121\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__9126\,
            I => \N_70\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__9121\,
            I => \N_70\
        );

    \I__811\ : CEMux
    port map (
            O => \N__9116\,
            I => \N__9113\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__9113\,
            I => \N__9110\
        );

    \I__809\ : Span4Mux_v
    port map (
            O => \N__9110\,
            I => \N__9107\
        );

    \I__808\ : Odrv4
    port map (
            O => \N__9107\,
            I => \N_26\
        );

    \I__807\ : InMux
    port map (
            O => \N__9104\,
            I => \this_vga_signals.mult1_un47_sum_cry_0\
        );

    \I__806\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__9098\,
            I => \N__9095\
        );

    \I__804\ : Odrv4
    port map (
            O => \N__9095\,
            I => \this_vga_signals.mult1_un40_sum_cry_1_s\
        );

    \I__803\ : InMux
    port map (
            O => \N__9092\,
            I => \this_vga_signals.mult1_un47_sum_cry_1\
        );

    \I__802\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9086\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__9086\,
            I => \this_vga_signals.mult1_un47_sum_axb_3\
        );

    \I__800\ : InMux
    port map (
            O => \N__9083\,
            I => \this_vga_signals.mult1_un47_sum_cry_2\
        );

    \I__799\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9074\
        );

    \I__798\ : InMux
    port map (
            O => \N__9079\,
            I => \N__9074\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__9074\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1\
        );

    \I__796\ : InMux
    port map (
            O => \N__9071\,
            I => \N__9068\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__9068\,
            I => \this_vga_signals.g2_0_x1\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__9065\,
            I => \this_vga_signals.g2_0_x0_cascade_\
        );

    \I__793\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__9059\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0_0\
        );

    \I__791\ : InMux
    port map (
            O => \N__9056\,
            I => \N__9053\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__9053\,
            I => \this_vga_signals.g2_0\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__788\ : InMux
    port map (
            O => \N__9047\,
            I => \N__9044\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__786\ : Odrv4
    port map (
            O => \N__9041\,
            I => \M_this_vga_signals_address_12\
        );

    \I__785\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__9035\,
            I => \this_vga_signals.g0_2\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__9032\,
            I => \N__9029\
        );

    \I__782\ : InMux
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__9026\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_1\
        );

    \I__780\ : InMux
    port map (
            O => \N__9023\,
            I => \this_vga_signals.mult1_un40_sum_cry_0\
        );

    \I__779\ : InMux
    port map (
            O => \N__9020\,
            I => \this_vga_signals.mult1_un40_sum_cry_1\
        );

    \I__778\ : InMux
    port map (
            O => \N__9017\,
            I => \this_vga_signals.mult1_un40_sum_cry_2\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__9014\,
            I => \this_vga_signals.if_N_6_mux_0_0_cascade_\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__9011\,
            I => \N__9008\
        );

    \I__775\ : InMux
    port map (
            O => \N__9008\,
            I => \N__9005\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__9005\,
            I => \M_this_vga_signals_address_8\
        );

    \I__773\ : CascadeMux
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__772\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8996\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__8996\,
            I => \M_this_vga_signals_address_11\
        );

    \I__770\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8990\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__8990\,
            I => \this_vga_signals.g0_0_a2_1\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__8987\,
            I => \N__8984\
        );

    \I__767\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__8981\,
            I => \M_this_vga_signals_address_9\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__8978\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_cascade_\
        );

    \I__764\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8972\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__8972\,
            I => \this_vga_ramdac.m16\
        );

    \I__762\ : IoInMux
    port map (
            O => \N__8969\,
            I => \N__8966\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__8966\,
            I => \N__8963\
        );

    \I__760\ : IoSpan4Mux
    port map (
            O => \N__8963\,
            I => \N__8960\
        );

    \I__759\ : IoSpan4Mux
    port map (
            O => \N__8960\,
            I => \N__8957\
        );

    \I__758\ : Span4Mux_s2_h
    port map (
            O => \N__8957\,
            I => \N__8954\
        );

    \I__757\ : Odrv4
    port map (
            O => \N__8954\,
            I => \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_2\
        );

    \I__756\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8948\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__8948\,
            I => \this_vga_ramdac.m19\
        );

    \I__754\ : IoInMux
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__752\ : Span4Mux_s2_h
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__751\ : Sp12to4
    port map (
            O => \N__8936\,
            I => \N__8933\
        );

    \I__750\ : Span12Mux_v
    port map (
            O => \N__8933\,
            I => \N__8930\
        );

    \I__749\ : Odrv12
    port map (
            O => \N__8930\,
            I => \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_3\
        );

    \I__748\ : IoInMux
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__746\ : Span4Mux_s2_h
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__8918\,
            I => \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_1\
        );

    \I__744\ : InMux
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__8912\,
            I => \this_vga_ramdac.i2_mux\
        );

    \I__742\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__8906\,
            I => \N__8900\
        );

    \I__740\ : InMux
    port map (
            O => \N__8905\,
            I => \N__8897\
        );

    \I__739\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8892\
        );

    \I__738\ : InMux
    port map (
            O => \N__8903\,
            I => \N__8892\
        );

    \I__737\ : Span4Mux_s3_h
    port map (
            O => \N__8900\,
            I => \N__8885\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__8897\,
            I => \N__8885\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__8892\,
            I => \N__8882\
        );

    \I__734\ : InMux
    port map (
            O => \N__8891\,
            I => \N__8877\
        );

    \I__733\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8877\
        );

    \I__732\ : Span4Mux_v
    port map (
            O => \N__8885\,
            I => \N__8870\
        );

    \I__731\ : Span4Mux_s3_h
    port map (
            O => \N__8882\,
            I => \N__8870\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__8877\,
            I => \N__8870\
        );

    \I__729\ : Span4Mux_h
    port map (
            O => \N__8870\,
            I => \N__8867\
        );

    \I__728\ : Odrv4
    port map (
            O => \N__8867\,
            I => \M_this_vram_read_data_0\
        );

    \I__727\ : InMux
    port map (
            O => \N__8864\,
            I => \N__8856\
        );

    \I__726\ : InMux
    port map (
            O => \N__8863\,
            I => \N__8856\
        );

    \I__725\ : InMux
    port map (
            O => \N__8862\,
            I => \N__8851\
        );

    \I__724\ : InMux
    port map (
            O => \N__8861\,
            I => \N__8851\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__8856\,
            I => \N__8846\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__8851\,
            I => \N__8843\
        );

    \I__721\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8838\
        );

    \I__720\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8838\
        );

    \I__719\ : Span4Mux_v
    port map (
            O => \N__8846\,
            I => \N__8835\
        );

    \I__718\ : Span4Mux_s3_h
    port map (
            O => \N__8843\,
            I => \N__8830\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__8838\,
            I => \N__8830\
        );

    \I__716\ : Span4Mux_h
    port map (
            O => \N__8835\,
            I => \N__8825\
        );

    \I__715\ : Span4Mux_h
    port map (
            O => \N__8830\,
            I => \N__8825\
        );

    \I__714\ : Odrv4
    port map (
            O => \N__8825\,
            I => \M_this_vram_read_data_2\
        );

    \I__713\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__8819\,
            I => \N__8812\
        );

    \I__711\ : InMux
    port map (
            O => \N__8818\,
            I => \N__8809\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__8817\,
            I => \N__8805\
        );

    \I__709\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8800\
        );

    \I__708\ : InMux
    port map (
            O => \N__8815\,
            I => \N__8800\
        );

    \I__707\ : Span4Mux_s3_h
    port map (
            O => \N__8812\,
            I => \N__8795\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__8809\,
            I => \N__8795\
        );

    \I__705\ : InMux
    port map (
            O => \N__8808\,
            I => \N__8790\
        );

    \I__704\ : InMux
    port map (
            O => \N__8805\,
            I => \N__8790\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__8800\,
            I => \N__8787\
        );

    \I__702\ : Span4Mux_v
    port map (
            O => \N__8795\,
            I => \N__8784\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__8790\,
            I => \N__8779\
        );

    \I__700\ : Span4Mux_s3_h
    port map (
            O => \N__8787\,
            I => \N__8779\
        );

    \I__699\ : Span4Mux_h
    port map (
            O => \N__8784\,
            I => \N__8774\
        );

    \I__698\ : Span4Mux_h
    port map (
            O => \N__8779\,
            I => \N__8774\
        );

    \I__697\ : Odrv4
    port map (
            O => \N__8774\,
            I => \M_this_vram_read_data_1\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__8771\,
            I => \N__8768\
        );

    \I__695\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8763\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__8767\,
            I => \N__8759\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__8766\,
            I => \N__8756\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__8763\,
            I => \N__8752\
        );

    \I__691\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8749\
        );

    \I__690\ : InMux
    port map (
            O => \N__8759\,
            I => \N__8744\
        );

    \I__689\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8744\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__8755\,
            I => \N__8740\
        );

    \I__687\ : Span4Mux_s3_h
    port map (
            O => \N__8752\,
            I => \N__8735\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__8749\,
            I => \N__8735\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__8744\,
            I => \N__8732\
        );

    \I__684\ : InMux
    port map (
            O => \N__8743\,
            I => \N__8727\
        );

    \I__683\ : InMux
    port map (
            O => \N__8740\,
            I => \N__8727\
        );

    \I__682\ : Span4Mux_v
    port map (
            O => \N__8735\,
            I => \N__8720\
        );

    \I__681\ : Span4Mux_s3_h
    port map (
            O => \N__8732\,
            I => \N__8720\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__8727\,
            I => \N__8720\
        );

    \I__679\ : Span4Mux_h
    port map (
            O => \N__8720\,
            I => \N__8717\
        );

    \I__678\ : Odrv4
    port map (
            O => \N__8717\,
            I => \M_this_vram_read_data_3\
        );

    \I__677\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8711\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__8711\,
            I => \N__8708\
        );

    \I__675\ : Span4Mux_s3_h
    port map (
            O => \N__8708\,
            I => \N__8700\
        );

    \I__674\ : InMux
    port map (
            O => \N__8707\,
            I => \N__8697\
        );

    \I__673\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8690\
        );

    \I__672\ : InMux
    port map (
            O => \N__8705\,
            I => \N__8690\
        );

    \I__671\ : InMux
    port map (
            O => \N__8704\,
            I => \N__8690\
        );

    \I__670\ : InMux
    port map (
            O => \N__8703\,
            I => \N__8687\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__8700\,
            I => \this_vga_ramdac.N_706_0\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__8697\,
            I => \this_vga_ramdac.N_706_0\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__8690\,
            I => \this_vga_ramdac.N_706_0\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__8687\,
            I => \this_vga_ramdac.N_706_0\
        );

    \I__665\ : InMux
    port map (
            O => \N__8678\,
            I => \N__8675\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__8675\,
            I => \this_vga_ramdac.i2_mux_0\
        );

    \I__663\ : IoInMux
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__661\ : IoSpan4Mux
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__660\ : IoSpan4Mux
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__659\ : IoSpan4Mux
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__658\ : Span4Mux_s3_h
    port map (
            O => \N__8657\,
            I => \N__8654\
        );

    \I__657\ : Odrv4
    port map (
            O => \N__8654\,
            I => \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_4\
        );

    \I__656\ : IoInMux
    port map (
            O => \N__8651\,
            I => \N__8648\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__654\ : Span4Mux_s2_h
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__653\ : Span4Mux_h
    port map (
            O => \N__8642\,
            I => \N__8639\
        );

    \I__652\ : Odrv4
    port map (
            O => \N__8639\,
            I => \N_94\
        );

    \I__651\ : IoInMux
    port map (
            O => \N__8636\,
            I => \N__8633\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__8633\,
            I => \N__8630\
        );

    \I__649\ : Span4Mux_s3_v
    port map (
            O => \N__8630\,
            I => \N__8627\
        );

    \I__648\ : Span4Mux_v
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__647\ : Span4Mux_v
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__646\ : Span4Mux_v
    port map (
            O => \N__8621\,
            I => \N__8618\
        );

    \I__645\ : Odrv4
    port map (
            O => \N__8618\,
            I => \N_274_i\
        );

    \I__644\ : IoInMux
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__8612\,
            I => \this_vga_signals.N_517_1\
        );

    \I__642\ : IoInMux
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__8606\,
            I => \N_205_i\
        );

    \I__640\ : IoInMux
    port map (
            O => \N__8603\,
            I => \N__8600\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__8600\,
            I => \N__8597\
        );

    \I__638\ : IoSpan4Mux
    port map (
            O => \N__8597\,
            I => \N__8594\
        );

    \I__637\ : Span4Mux_s0_h
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__8591\,
            I => \this_vga_ramdac.M_this_rgb_d_3_0_dreg\
        );

    \I__635\ : CascadeMux
    port map (
            O => \N__8588\,
            I => \this_vga_ramdac.m5_cascade_\
        );

    \I__634\ : IoInMux
    port map (
            O => \N__8585\,
            I => \N__8582\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__8582\,
            I => \N__8579\
        );

    \I__632\ : IoSpan4Mux
    port map (
            O => \N__8579\,
            I => \N__8576\
        );

    \I__631\ : Span4Mux_s2_h
    port map (
            O => \N__8576\,
            I => \N__8573\
        );

    \I__630\ : Odrv4
    port map (
            O => \N__8573\,
            I => \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_0\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_1_cry_8\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_16_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_21_0_\
        );

    \IN_MUX_bfv_16_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_internal_address_q_cry_7\,
            carryinitout => \bfn_16_22_0_\
        );

    \IN_MUX_bfv_31_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_31_23_0_\
        );

    \IN_MUX_bfv_31_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_external_address_q_cry_7\,
            carryinitout => \bfn_31_24_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_data_count_q_cry_7\,
            carryinitout => \bfn_15_24_0_\
        );

    \IN_MUX_bfv_15_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO\,
            carryinitout => \bfn_15_25_0_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIRV75_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__16529\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_684_g\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI6RKH5_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8615\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_517_1_g\
        );

    \this_reset_cond.M_stage_q_RNI6VB7_3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19594\,
            GLOBALBUFFEROUTPUT => \M_this_state_q_nss_g_0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI6RKH5_9_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17143\,
            in2 => \_gnd_net_\,
            in3 => \N__15497\,
            lcout => \this_vga_signals.N_517_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_205_i_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__20214\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20641\,
            lcout => \N_205_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_0_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000000000"
        )
    port map (
            in0 => \N__8822\,
            in1 => \N__8909\,
            in2 => \N__8771\,
            in3 => \N__8714\,
            lcout => \this_vga_ramdac.M_this_rgb_d_3_0_dreg\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m5_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__8863\,
            in1 => \N__8818\,
            in2 => \_gnd_net_\,
            in3 => \N__8905\,
            lcout => OPEN,
            ltout => \this_vga_ramdac.m5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_1_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__8762\,
            in1 => \N__8864\,
            in2 => \N__8588\,
            in3 => \N__8707\,
            lcout => \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001110010111"
        )
    port map (
            in0 => \N__8861\,
            in1 => \N__8816\,
            in2 => \N__8766\,
            in3 => \N__8903\,
            lcout => \this_vga_ramdac.m16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010100101011"
        )
    port map (
            in0 => \N__8862\,
            in1 => \N__8815\,
            in2 => \N__8767\,
            in3 => \N__8904\,
            lcout => \this_vga_ramdac.m19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_3_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__8975\,
            in1 => \N__8705\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_4_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8706\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8951\,
            lcout => \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_2_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8704\,
            in2 => \_gnd_net_\,
            in3 => \N__8915\,
            lcout => \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111101"
        )
    port map (
            in0 => \N__8849\,
            in1 => \N__8808\,
            in2 => \N__8755\,
            in3 => \N__8890\,
            lcout => \this_vga_ramdac.i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_q_250_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23823\,
            in2 => \_gnd_net_\,
            in3 => \N__24787\,
            lcout => \this_vga_ramdac.N_706_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010000111011"
        )
    port map (
            in0 => \N__8891\,
            in1 => \N__8850\,
            in2 => \N__8817\,
            in3 => \N__8743\,
            lcout => \this_vga_ramdac.i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_5_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8703\,
            in2 => \_gnd_net_\,
            in3 => \N__8678\,
            lcout => \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNID8NA3_9_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010111"
        )
    port map (
            in0 => \N__20218\,
            in1 => \N__9872\,
            in2 => \N__13485\,
            in3 => \N__16642\,
            lcout => \N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIJVML2_9_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__16643\,
            in1 => \N__9868\,
            in2 => \_gnd_net_\,
            in3 => \N__13486\,
            lcout => \N_274_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000110111"
        )
    port map (
            in0 => \N__9506\,
            in1 => \N__9629\,
            in2 => \N__14132\,
            in3 => \N__14572\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_6_mux_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNINGUT4R3_7_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000100010"
        )
    port map (
            in0 => \N__23853\,
            in1 => \N__8993\,
            in2 => \N__9014\,
            in3 => \N__9056\,
            lcout => \M_this_vga_signals_address_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI6UL1Q3_7_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__23852\,
            in1 => \N__12095\,
            in2 => \_gnd_net_\,
            in3 => \N__12200\,
            lcout => \M_this_vga_signals_address_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_a2_1_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011111101000"
        )
    port map (
            in0 => \N__9584\,
            in1 => \N__14376\,
            in2 => \N__14582\,
            in3 => \N__9667\,
            lcout => \this_vga_signals.g0_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_x2_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13987\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14122\,
            lcout => \this_vga_signals.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIR4HAL91_7_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__23851\,
            in1 => \N__9596\,
            in2 => \_gnd_net_\,
            in3 => \N__9080\,
            lcout => \M_this_vga_signals_address_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_7_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101001111010"
        )
    port map (
            in0 => \N__14375\,
            in1 => \N__9583\,
            in2 => \N__9668\,
            in3 => \N__14565\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_N_3_i_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9038\,
            in1 => \N__11285\,
            in2 => \N__9032\,
            in3 => \N__12377\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_0_x1_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110101111000"
        )
    port map (
            in0 => \N__14564\,
            in1 => \N__9504\,
            in2 => \N__8978\,
            in3 => \N__9624\,
            lcout => \this_vga_signals.g2_0_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI9OGF9_5_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15135\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12567\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_0_x0_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000110101"
        )
    port map (
            in0 => \N__9625\,
            in1 => \N__9505\,
            in2 => \N__14581\,
            in3 => \N__9079\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_0_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_0_ns_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9071\,
            in2 => \N__9065\,
            in3 => \N__9062\,
            lcout => \this_vga_signals.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNINSNSM_7_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__12569\,
            in1 => \N__23860\,
            in2 => \_gnd_net_\,
            in3 => \N__12644\,
            lcout => \M_this_vga_signals_address_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12089\,
            in1 => \N__12568\,
            in2 => \N__15155\,
            in3 => \N__12194\,
            lcout => \this_vga_signals.g0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100101011"
        )
    port map (
            in0 => \N__12193\,
            in1 => \N__14377\,
            in2 => \N__15449\,
            in3 => \N__12090\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_0_c_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16343\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \this_vga_signals.mult1_un40_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_1_s_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9185\,
            in2 => \N__9239\,
            in3 => \N__9023\,
            lcout => \this_vga_signals.mult1_un40_sum_cry_1_s\,
            ltout => OPEN,
            carryin => \this_vga_signals.mult1_un40_sum_cry_0\,
            carryout => \this_vga_signals.mult1_un40_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.mult1_un40_sum_cry_1_THRU_LUT4_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9131\,
            in2 => \N__9149\,
            in3 => \N__9020\,
            lcout => \this_vga_signals.mult1_un40_sum_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_vga_signals.mult1_un40_sum_cry_1\,
            carryout => \this_vga_signals.mult1_un40_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.mult1_un40_sum_cry_2_THRU_LUT4_0_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9017\,
            lcout => \this_vga_signals.mult1_un40_sum_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_2_c_inv_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9184\,
            in1 => \N__9144\,
            in2 => \_gnd_net_\,
            in3 => \N__9129\,
            lcout => \N_70\,
            ltout => \N_70_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_2_l_fx_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9158\,
            in3 => \N__9245\,
            lcout => \G_501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_axb_3_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9155\,
            in1 => \N__9145\,
            in2 => \N__9222\,
            in3 => \N__9130\,
            lcout => \this_vga_signals.mult1_un47_sum_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_vram_write_en_i_0_i_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__22385\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23552\,
            lcout => \N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_cry_0_c_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16220\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \this_vga_signals.mult1_un47_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_cry_1_s_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9287\,
            in2 => \N__9203\,
            in3 => \N__9104\,
            lcout => \this_vga_signals.mult1_un47_sum_cry_1_s\,
            ltout => OPEN,
            carryin => \this_vga_signals.mult1_un47_sum_cry_0\,
            carryout => \this_vga_signals.mult1_un47_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_axb_3_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9265\,
            in1 => \N__9101\,
            in2 => \N__9227\,
            in3 => \N__9092\,
            lcout => \this_vga_signals.mult1_un54_sum_axb_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.mult1_un47_sum_cry_1\,
            carryout => \this_vga_signals.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_s_3_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__9089\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9083\,
            lcout => \this_vga_signals.mult1_un47_sum_s_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_2_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011110011110"
        )
    port map (
            in0 => \N__15794\,
            in1 => \N__15890\,
            in2 => \N__16004\,
            in3 => \N__16101\,
            lcout => \this_vga_signals.mult1_un40_sum_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_1_l_fx_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15793\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9177\,
            lcout => \this_vga_signals.mult1_un40_sum_axb_1_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_s_3_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9223\,
            lcout => \this_vga_signals.mult1_un40_sum_s_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_cry_0_c_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18106\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \this_vga_signals.mult1_un61_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_cry_1_s_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13841\,
            in2 => \N__9305\,
            in3 => \N__9194\,
            lcout => \this_vga_signals.mult1_un61_sum_cry_1_s\,
            ltout => OPEN,
            carryin => \this_vga_signals.mult1_un61_sum_cry_0\,
            carryout => \this_vga_signals.mult1_un61_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_axb_3_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12877\,
            in1 => \N__9164\,
            in2 => \N__9347\,
            in3 => \N__9191\,
            lcout => \this_vga_signals.mult1_un68_sum_axb_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.mult1_un61_sum_cry_1\,
            carryout => \this_vga_signals.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_s_3_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9326\,
            in2 => \_gnd_net_\,
            in3 => \N__9188\,
            lcout => \this_vga_signals.mult1_un61_sum_s_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNITQQM_9_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16581\,
            in2 => \_gnd_net_\,
            in3 => \N__13804\,
            lcout => \this_vga_signals.CO1_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNICJJV_9_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000110100111"
        )
    port map (
            in0 => \N__15889\,
            in1 => \N__15792\,
            in2 => \N__16003\,
            in3 => \N__16100\,
            lcout => \this_vga_signals.N_70_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_sbtinv_3_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9301\,
            lcout => \this_vga_signals.mult1_un54_sum_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_cry_0_c_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17006\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \this_vga_signals.mult1_un54_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_cry_1_s_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11645\,
            in2 => \N__9275\,
            in3 => \N__9338\,
            lcout => \this_vga_signals.mult1_un54_sum_cry_1_s\,
            ltout => OPEN,
            carryin => \this_vga_signals.mult1_un54_sum_cry_0\,
            carryout => \this_vga_signals.mult1_un54_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_axb_3_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9300\,
            in1 => \N__9335\,
            in2 => \N__9254\,
            in3 => \N__9320\,
            lcout => \this_vga_signals.mult1_un61_sum_axb_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.mult1_un54_sum_cry_1\,
            carryout => \this_vga_signals.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_s_3_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__9317\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9308\,
            lcout => \this_vga_signals.mult1_un54_sum_s_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI54V41_5_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__14342\,
            in1 => \N__15423\,
            in2 => \_gnd_net_\,
            in3 => \N__15150\,
            lcout => \this_vga_signals.vsync_1_0_a2_6_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_sbtinv_5_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16338\,
            lcout => \this_vga_signals.M_hcounter_q_i_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_sbtinv_3_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9271\,
            lcout => \this_vga_signals.mult1_un47_sum_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m8_0_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001101010101"
        )
    port map (
            in0 => \N__9848\,
            in1 => \N__11849\,
            in2 => \N__13988\,
            in3 => \N__10598\,
            lcout => \this_ppu.M_N_13_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m9_i_x3_0_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14109\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13985\,
            lcout => \this_ppu.M_m9_i_x3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_c_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14498\,
            in1 => \N__14107\,
            in2 => \_gnd_net_\,
            in3 => \N__14335\,
            lcout => \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m5_0_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101010100"
        )
    port map (
            in0 => \N__10599\,
            in1 => \N__13981\,
            in2 => \N__11857\,
            in3 => \N__9847\,
            lcout => OPEN,
            ltout => \this_ppu.M_N_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m11_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__14144\,
            in1 => \N__14108\,
            in2 => \N__9374\,
            in3 => \N__9371\,
            lcout => OPEN,
            ltout => \this_ppu.M_N_15_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_0_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9365\,
            in1 => \N__15202\,
            in2 => \N__9359\,
            in3 => \N__15422\,
            lcout => \this_ppu.N_277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m12_0_x3_s_0_1_0_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001011101101"
        )
    port map (
            in0 => \N__14556\,
            in1 => \N__10499\,
            in2 => \N__14129\,
            in3 => \N__10492\,
            lcout => OPEN,
            ltout => \this_ppu.M_m12_0_x3_s_0_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m12_0_x3_s_0_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011111100001"
        )
    port map (
            in0 => \N__14118\,
            in1 => \N__14557\,
            in2 => \N__9356\,
            in3 => \N__9836\,
            lcout => \this_ppu.M_m12_0_x3_out_0\,
            ltout => \this_ppu.M_m12_0_x3_out_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_4_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111011"
        )
    port map (
            in0 => \N__14114\,
            in1 => \N__13986\,
            in2 => \N__9353\,
            in3 => \N__9475\,
            lcout => \this_ppu.M_m1_e_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_m12_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__15398\,
            in1 => \N__10518\,
            in2 => \_gnd_net_\,
            in3 => \N__10535\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_m14_0_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101001010001"
        )
    port map (
            in0 => \N__10493\,
            in1 => \N__14113\,
            in2 => \N__9350\,
            in3 => \N__14555\,
            lcout => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_c3_0,
            ltout => \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m1_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9479\,
            in3 => \N__10577\,
            lcout => \this_ppu.M_mZ0Z1\,
            ltout => \this_ppu.M_mZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIMJNMSC_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100000000"
        )
    port map (
            in0 => \N__9476\,
            in1 => \N__9421\,
            in2 => \N__9467\,
            in3 => \N__10547\,
            lcout => \this_ppu.M_m1_e_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__16103\,
            in1 => \N__15888\,
            in2 => \_gnd_net_\,
            in3 => \N__16002\,
            lcout => \N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un68_sum_axb1_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11858\,
            in1 => \N__10601\,
            in2 => \N__14580\,
            in3 => \N__9835\,
            lcout => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axb1,
            ltout => \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m12_0_o3_0_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001101"
        )
    port map (
            in0 => \N__10576\,
            in1 => \N__14130\,
            in2 => \N__9443\,
            in3 => \N__9440\,
            lcout => \this_ppu.M_N_16_1\,
            ltout => \this_ppu.M_N_16_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_3_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100000000"
        )
    port map (
            in0 => \N__9434\,
            in1 => \N__9394\,
            in2 => \N__9428\,
            in3 => \N__10546\,
            lcout => OPEN,
            ltout => \this_ppu.M_m1_e_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_2_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000000000"
        )
    port map (
            in0 => \N__9425\,
            in1 => \N__9410\,
            in2 => \N__9404\,
            in3 => \N__9401\,
            lcout => \this_ppu.M_N_3_mux_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI8H768U_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011110000"
        )
    port map (
            in0 => \N__9395\,
            in1 => \N__9386\,
            in2 => \N__24800\,
            in3 => \N__9380\,
            lcout => \this_ppu.N_256_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_current_q_0_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10995\,
            in2 => \N__22378\,
            in3 => \N__22386\,
            lcout => \M_this_ppu_vram_addr_0\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \this_ppu.un1_M_current_q_cry_0\,
            clk => \N__25021\,
            ce => 'H',
            sr => \N__9515\
        );

    \this_ppu.M_current_q_1_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10721\,
            in2 => \_gnd_net_\,
            in3 => \N__9533\,
            lcout => \M_this_ppu_vram_addr_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_current_q_cry_0\,
            carryout => \this_ppu.un1_M_current_q_cry_1\,
            clk => \N__25021\,
            ce => 'H',
            sr => \N__9515\
        );

    \this_ppu.M_current_q_2_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9936\,
            in2 => \_gnd_net_\,
            in3 => \N__9530\,
            lcout => \M_this_ppu_vram_addr_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_current_q_cry_1\,
            carryout => \this_ppu.un1_M_current_q_cry_2\,
            clk => \N__25021\,
            ce => 'H',
            sr => \N__9515\
        );

    \this_ppu.M_current_q_3_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10860\,
            in2 => \_gnd_net_\,
            in3 => \N__9527\,
            lcout => \M_this_ppu_vram_addr_3\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_current_q_cry_2\,
            carryout => \this_ppu.un1_M_current_q_cry_3\,
            clk => \N__25021\,
            ce => 'H',
            sr => \N__9515\
        );

    \this_ppu.M_current_q_4_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10223\,
            in2 => \_gnd_net_\,
            in3 => \N__9524\,
            lcout => \M_this_ppu_vram_addr_4\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_current_q_cry_3\,
            carryout => \this_ppu.un1_M_current_q_cry_4\,
            clk => \N__25021\,
            ce => 'H',
            sr => \N__9515\
        );

    \this_ppu.M_current_q_5_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10364\,
            in2 => \_gnd_net_\,
            in3 => \N__9521\,
            lcout => \M_this_ppu_vram_addr_5\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_current_q_cry_4\,
            carryout => \this_ppu.un1_M_current_q_cry_5\,
            clk => \N__25021\,
            ce => 'H',
            sr => \N__9515\
        );

    \this_ppu.M_current_q_6_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10073\,
            in2 => \_gnd_net_\,
            in3 => \N__9518\,
            lcout => \M_this_ppu_vram_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25021\,
            ce => 'H',
            sr => \N__9515\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_0_5_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12198\,
            in1 => \N__12466\,
            in2 => \N__11204\,
            in3 => \N__9649\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12364\,
            in1 => \N__11277\,
            in2 => \_gnd_net_\,
            in3 => \N__14373\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIN3CPT8_7_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__23850\,
            in1 => \_gnd_net_\,
            in2 => \N__11288\,
            in3 => \N__12365\,
            lcout => \M_this_vga_signals_address_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_9_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11278\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12363\,
            lcout => \this_vga_signals.N_9_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12467\,
            in1 => \N__11200\,
            in2 => \N__9653\,
            in3 => \N__12199\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIGU2FNB_5_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__11279\,
            in1 => \_gnd_net_\,
            in2 => \N__9572\,
            in3 => \N__9569\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_x2_0_0_a3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_14_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110111010111"
        )
    port map (
            in0 => \N__9563\,
            in1 => \N__9704\,
            in2 => \N__9554\,
            in3 => \N__10610\,
            lcout => \this_vga_signals.N_5_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_19_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12069\,
            in1 => \N__15442\,
            in2 => \_gnd_net_\,
            in3 => \N__12166\,
            lcout => \this_vga_signals.N_9_i_0_0\,
            ltout => \this_vga_signals.N_9_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_x1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001111100011"
        )
    port map (
            in0 => \N__14541\,
            in1 => \N__14333\,
            in2 => \N__9551\,
            in3 => \N__12367\,
            lcout => \this_vga_signals.g0_2_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI6CQQNK_2_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9608\,
            in1 => \N__9590\,
            in2 => \_gnd_net_\,
            in3 => \N__11284\,
            lcout => \this_vga_signals.N_57_i_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_x0_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100110010001"
        )
    port map (
            in0 => \N__14374\,
            in1 => \N__9548\,
            in2 => \N__14576\,
            in3 => \N__12368\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_2_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_ns_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11283\,
            in2 => \N__9542\,
            in3 => \N__9539\,
            lcout => \this_vga_signals.N_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__12167\,
            in1 => \_gnd_net_\,
            in2 => \N__15452\,
            in3 => \N__12070\,
            lcout => \this_vga_signals.N_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI5RUBJ1_5_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15136\,
            in1 => \N__12560\,
            in2 => \N__14579\,
            in3 => \N__12165\,
            lcout => \this_vga_signals.m6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010010111000"
        )
    port map (
            in0 => \N__12164\,
            in1 => \N__11339\,
            in2 => \N__9641\,
            in3 => \N__12068\,
            lcout => \this_vga_signals.mult1_un61_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_11_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__9674\,
            in1 => \N__12280\,
            in2 => \N__9692\,
            in3 => \N__12268\,
            lcout => \this_vga_signals.if_i3_mux_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI820378_2_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110000110110"
        )
    port map (
            in0 => \N__14369\,
            in1 => \N__11381\,
            in2 => \N__14577\,
            in3 => \N__12373\,
            lcout => \this_vga_signals.M_vcounter_q_RNI820378Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_8_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15362\,
            in1 => \N__12084\,
            in2 => \_gnd_net_\,
            in3 => \N__12191\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101001111010"
        )
    port map (
            in0 => \N__14372\,
            in1 => \N__11287\,
            in2 => \N__9602\,
            in3 => \N__12375\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14551\,
            in2 => \N__9599\,
            in3 => \N__9710\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI820378_0_2_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011001101100"
        )
    port map (
            in0 => \N__14370\,
            in1 => \N__11380\,
            in2 => \N__14578\,
            in3 => \N__12372\,
            lcout => \this_vga_signals.M_vcounter_q_RNI820378_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_0_a3_2_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14378\,
            in1 => \N__12083\,
            in2 => \N__15425\,
            in3 => \N__12190\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_3_0_a3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_1_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011110111101"
        )
    port map (
            in0 => \N__14371\,
            in1 => \N__11286\,
            in2 => \N__9713\,
            in3 => \N__12374\,
            lcout => \this_vga_signals.g2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m10_0_a4_1_1_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__12548\,
            in1 => \N__14303\,
            in2 => \N__15125\,
            in3 => \N__15414\,
            lcout => \this_vga_signals.if_m10_0_a4_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_1_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__14305\,
            in1 => \N__12082\,
            in2 => \N__15448\,
            in3 => \N__12189\,
            lcout => \this_vga_signals.g1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_4_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12724\,
            lcout => \this_vga_signals.N_188_0\,
            ltout => \this_vga_signals.N_188_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIEC471_9_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15191\,
            in2 => \N__9695\,
            in3 => \N__16613\,
            lcout => \this_vga_signals.CO0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m10_0_a4_0_0_0_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__12550\,
            in1 => \N__14304\,
            in2 => \N__15126\,
            in3 => \N__15415\,
            lcout => \this_vga_signals.if_m10_0_a4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_3_0_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11324\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12632\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_12_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \N__12549\,
            in1 => \N__11398\,
            in2 => \N__9683\,
            in3 => \N__9680\,
            lcout => \this_vga_signals.if_N_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000110110111"
        )
    port map (
            in0 => \N__15044\,
            in1 => \N__13700\,
            in2 => \N__15447\,
            in3 => \N__12808\,
            lcout => \this_vga_signals.mult1_un47_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_ns_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11453\,
            in1 => \N__9722\,
            in2 => \_gnd_net_\,
            in3 => \N__11420\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_c3_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011010000"
        )
    port map (
            in0 => \N__13805\,
            in1 => \N__13160\,
            in2 => \N__9728\,
            in3 => \N__11725\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__13697\,
            in1 => \N__13912\,
            in2 => \N__9725\,
            in3 => \N__15029\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_5_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13038\,
            lcout => \this_vga_signals_M_vcounter_q_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24981\,
            ce => \N__15520\,
            sr => \N__15493\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_0_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9803\,
            in2 => \N__9821\,
            in3 => \N__9784\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_1_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001100000"
        )
    port map (
            in0 => \N__13315\,
            in1 => \N__13911\,
            in2 => \N__13705\,
            in3 => \N__12806\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13107\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24981\,
            ce => \N__15520\,
            sr => \N__15493\
        );

    \this_vga_signals.M_vcounter_q_0_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17144\,
            in1 => \N__13965\,
            in2 => \N__16682\,
            in3 => \N__16678\,
            lcout => \this_vga_signals_M_vcounter_q_0\,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            clk => \N__24986\,
            ce => 'H',
            sr => \N__15492\
        );

    \this_vga_signals.M_vcounter_q_1_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17146\,
            in1 => \N__14066\,
            in2 => \_gnd_net_\,
            in3 => \N__9716\,
            lcout => \this_vga_signals_M_vcounter_q_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            clk => \N__24986\,
            ce => 'H',
            sr => \N__15492\
        );

    \this_vga_signals.M_vcounter_q_2_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17145\,
            in1 => \N__14470\,
            in2 => \_gnd_net_\,
            in3 => \N__9752\,
            lcout => \this_vga_signals_M_vcounter_q_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            clk => \N__24986\,
            ce => 'H',
            sr => \N__15492\
        );

    \this_vga_signals.M_vcounter_q_3_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17147\,
            in1 => \N__14254\,
            in2 => \_gnd_net_\,
            in3 => \N__9749\,
            lcout => \this_vga_signals_M_vcounter_q_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            clk => \N__24986\,
            ce => 'H',
            sr => \N__15492\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15358\,
            in2 => \_gnd_net_\,
            in3 => \N__9746\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15083\,
            in2 => \_gnd_net_\,
            in3 => \N__9743\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13690\,
            in2 => \_gnd_net_\,
            in3 => \N__9740\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13584\,
            in2 => \_gnd_net_\,
            in3 => \N__9737\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13797\,
            in2 => \_gnd_net_\,
            in3 => \N__9734\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16630\,
            in2 => \_gnd_net_\,
            in3 => \N__9731\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_9_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13173\,
            lcout => \this_vga_signals_M_vcounter_q_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24994\,
            ce => \N__15518\,
            sr => \N__15490\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_9_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13174\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24994\,
            ce => \N__15518\,
            sr => \N__15490\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13081\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24994\,
            ce => \N__15518\,
            sr => \N__15490\
        );

    \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13080\,
            lcout => \this_vga_signals_M_vcounter_q_8_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24994\,
            ce => \N__15518\,
            sr => \N__15490\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_c2_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010111011"
        )
    port map (
            in0 => \N__13022\,
            in1 => \N__11767\,
            in2 => \_gnd_net_\,
            in3 => \N__12725\,
            lcout => \this_vga_signals.mult1_un40_sum_1_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_ac0_3_0_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100010011"
        )
    port map (
            in0 => \N__13321\,
            in1 => \N__11674\,
            in2 => \N__11561\,
            in3 => \N__13021\,
            lcout => \this_vga_signals.mult1_un40_sum_0_c3_0\,
            ltout => \this_vga_signals.mult1_un40_sum_0_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x0_3_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001011000000"
        )
    port map (
            in0 => \N__11569\,
            in1 => \N__9894\,
            in2 => \N__9824\,
            in3 => \N__11755\,
            lcout => \this_vga_signals.mult1_un40_sum_m_x0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_7_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110110011001"
        )
    port map (
            in0 => \N__9817\,
            in1 => \N__9802\,
            in2 => \N__11447\,
            in3 => \N__9788\,
            lcout => \this_vga_signals.N_81_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x1_3_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000010100"
        )
    port map (
            in0 => \N__9895\,
            in1 => \N__11756\,
            in2 => \N__11573\,
            in3 => \N__9773\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_m_x1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_3_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9767\,
            in2 => \N__9761\,
            in3 => \N__9758\,
            lcout => \this_vga_signals.mult1_un40_sum_m_ns_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m12_0_o2_381_10_1_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101010101"
        )
    port map (
            in0 => \N__15201\,
            in1 => \N__14301\,
            in2 => \N__13370\,
            in3 => \N__15127\,
            lcout => \this_ppu.M_m12_0_o2_381_10Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_axbxc2_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111011101"
        )
    port map (
            in0 => \N__13698\,
            in1 => \N__11557\,
            in2 => \_gnd_net_\,
            in3 => \N__13317\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_2_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__11738\,
            in1 => \N__9899\,
            in2 => \N__9878\,
            in3 => \N__11675\,
            lcout => \this_vga_signals.mult1_un40_sum_m_ns_2\,
            ltout => \this_vga_signals.mult1_un40_sum_m_ns_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__13929\,
            in1 => \_gnd_net_\,
            in2 => \N__9875\,
            in3 => \N__15093\,
            lcout => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI65531_6_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__12943\,
            in1 => \N__13369\,
            in2 => \_gnd_net_\,
            in3 => \N__13699\,
            lcout => \this_vga_signals.N_196_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100110001"
        )
    port map (
            in0 => \N__13928\,
            in1 => \N__13211\,
            in2 => \N__13322\,
            in3 => \N__11879\,
            lcout => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0,
            ltout => \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axb1_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9851\,
            in3 => \N__13930\,
            lcout => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un54_sum_axb1,
            ltout => \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un54_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m7_1_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110000001"
        )
    port map (
            in0 => \N__13977\,
            in1 => \N__11835\,
            in2 => \N__9839\,
            in3 => \N__10600\,
            lcout => \this_ppu.M_m7Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100000000"
        )
    port map (
            in0 => \N__11630\,
            in1 => \N__10491\,
            in2 => \N__14561\,
            in3 => \N__11975\,
            lcout => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_c3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_m3_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011011101"
        )
    port map (
            in0 => \N__14345\,
            in1 => \N__13931\,
            in2 => \_gnd_net_\,
            in3 => \N__11954\,
            lcout => this_vga_signals_un4_lcounter_if_i1_mux,
            ltout => \this_vga_signals_un4_lcounter_if_i1_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__11955\,
            in1 => \_gnd_net_\,
            in2 => \N__10604\,
            in3 => \N__10519\,
            lcout => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0,
            ltout => \this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011111100001"
        )
    port map (
            in0 => \N__11933\,
            in1 => \N__11831\,
            in2 => \N__10580\,
            in3 => \N__11786\,
            lcout => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m7_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__14512\,
            in1 => \N__14091\,
            in2 => \_gnd_net_\,
            in3 => \N__10565\,
            lcout => OPEN,
            ltout => \this_ppu.M_N_11_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIFN38L2_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__10559\,
            in1 => \N__14699\,
            in2 => \N__10550\,
            in3 => \N__15094\,
            lcout => \this_ppu.M_m12_0_o2_381_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d_m1_0_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11956\,
            in1 => \N__10534\,
            in2 => \N__10523\,
            in3 => \N__11844\,
            lcout => this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_m14_0_x3_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__14346\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11830\,
            lcout => \this_vga_signals_un4_lcounter_if_N_7_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10365\,
            in1 => \N__10224\,
            in2 => \N__10083\,
            in3 => \N__9935\,
            lcout => OPEN,
            ltout => \this_ppu.un1_M_state_d8_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100101010"
        )
    port map (
            in0 => \N__22365\,
            in1 => \N__10691\,
            in2 => \N__9908\,
            in3 => \N__9905\,
            lcout => \M_this_ppu_vram_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25012\,
            ce => 'H',
            sr => \N__24743\
        );

    \this_ppu.M_state_q_RNO_1_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10994\,
            in1 => \N__10859\,
            in2 => \N__10728\,
            in3 => \N__22363\,
            lcout => \this_ppu.un1_M_state_d8_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__22811\,
            in1 => \N__22085\,
            in2 => \N__22301\,
            in3 => \N__21818\,
            lcout => OPEN,
            ltout => \M_this_sprites_ram_read_data_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_vram_write_data_0_i_0_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__20882\,
            in1 => \N__23501\,
            in2 => \N__10685\,
            in3 => \N__22364\,
            lcout => \M_this_vram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_0_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10670\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_2_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10619\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__10658\,
            in1 => \N__14513\,
            in2 => \N__11663\,
            in3 => \N__13706\,
            lcout => this_vga_signals_vsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_1_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10625\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_16_x0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001101110"
        )
    port map (
            in0 => \N__11996\,
            in1 => \N__14384\,
            in2 => \N__12376\,
            in3 => \N__14574\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_16_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_16_ns_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__11273\,
            in1 => \_gnd_net_\,
            in2 => \N__10613\,
            in3 => \N__12305\,
            lcout => \this_vga_signals.g3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_a2_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12091\,
            in1 => \N__11271\,
            in2 => \N__14387\,
            in3 => \N__11213\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__11274\,
            in1 => \N__14126\,
            in2 => \_gnd_net_\,
            in3 => \N__12362\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__14383\,
            in1 => \N__11174\,
            in2 => \N__11168\,
            in3 => \N__11165\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_axbxc3_3_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI5DK9PN1_7_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__23854\,
            in1 => \N__12206\,
            in2 => \N__11159\,
            in3 => \N__11138\,
            lcout => this_vga_signals_address_0_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011100100001"
        )
    port map (
            in0 => \N__11144\,
            in1 => \N__14127\,
            in2 => \N__11132\,
            in3 => \N__14575\,
            lcout => \this_vga_signals.mult1_un75_sum_c2_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11272\,
            in1 => \N__11219\,
            in2 => \N__11123\,
            in3 => \N__12361\,
            lcout => \this_vga_signals.g3_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_1_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12171\,
            in1 => \N__12065\,
            in2 => \N__15153\,
            in3 => \N__12561\,
            lcout => \this_vga_signals.g3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_N_4_i_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12456\,
            in1 => \N__11193\,
            in2 => \N__12088\,
            in3 => \N__12169\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_2_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011101000"
        )
    port map (
            in0 => \N__14540\,
            in1 => \N__14365\,
            in2 => \N__11114\,
            in3 => \N__11275\,
            lcout => \this_vga_signals.g1_2\,
            ltout => \this_vga_signals.g1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_m2_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011100010010"
        )
    port map (
            in0 => \N__14366\,
            in1 => \N__15446\,
            in2 => \N__11291\,
            in3 => \N__12298\,
            lcout => \this_vga_signals.N_57_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100101011"
        )
    port map (
            in0 => \N__12172\,
            in1 => \N__15429\,
            in2 => \N__14386\,
            in3 => \N__12067\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIOH6PPC_5_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11276\,
            in1 => \N__12575\,
            in2 => \N__11222\,
            in3 => \N__12366\,
            lcout => \this_vga_signals.m48_i_x4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011010100"
        )
    port map (
            in0 => \N__12170\,
            in1 => \N__15430\,
            in2 => \N__14385\,
            in3 => \N__12066\,
            lcout => \this_vga_signals.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_N_4_i_0_x_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__12457\,
            in1 => \N__11194\,
            in2 => \_gnd_net_\,
            in3 => \N__12168\,
            lcout => \this_vga_signals.N_4_i_0_x\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_N_4_i_0_1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110011011110"
        )
    port map (
            in0 => \N__12533\,
            in1 => \N__15105\,
            in2 => \N__15450\,
            in3 => \N__12383\,
            lcout => \this_vga_signals.N_4_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100011010"
        )
    port map (
            in0 => \N__15104\,
            in1 => \N__12532\,
            in2 => \N__15424\,
            in3 => \N__12639\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110001000101"
        )
    port map (
            in0 => \N__11330\,
            in1 => \N__12660\,
            in2 => \N__11180\,
            in3 => \N__11465\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.g0_0_i_o3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11177\,
            in3 => \N__12175\,
            lcout => \this_vga_signals.N_81_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m10_0_x2_0_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12534\,
            in1 => \N__14306\,
            in2 => \N__15451\,
            in3 => \N__15106\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m10_0_x2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m10_0_a4_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__11405\,
            in1 => \N__12071\,
            in2 => \N__11357\,
            in3 => \N__12174\,
            lcout => \this_vga_signals.if_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12817\,
            in1 => \N__11495\,
            in2 => \N__11354\,
            in3 => \N__11464\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1\,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m10_0_x2_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12661\,
            in1 => \N__11399\,
            in2 => \N__11345\,
            in3 => \N__12072\,
            lcout => \this_vga_signals.if_N_7_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000001"
        )
    port map (
            in0 => \N__11494\,
            in1 => \N__11540\,
            in2 => \N__11524\,
            in3 => \N__12807\,
            lcout => \this_vga_signals.mult1_un47_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un47_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11314\,
            in2 => \N__11342\,
            in3 => \N__12628\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m2_1_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000100100100"
        )
    port map (
            in0 => \N__14302\,
            in1 => \N__15064\,
            in2 => \N__15427\,
            in3 => \N__12538\,
            lcout => \this_vga_signals.if_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_x1_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__12536\,
            in1 => \N__15369\,
            in2 => \N__11329\,
            in3 => \N__12630\,
            lcout => \this_vga_signals.if_m10_0_a4_1_0_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_x0_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100010000100"
        )
    port map (
            in0 => \N__12631\,
            in1 => \N__15432\,
            in2 => \N__11325\,
            in3 => \N__12537\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m10_0_a4_1_0_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_ns_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11414\,
            in2 => \N__11408\,
            in3 => \N__11397\,
            lcout => \this_vga_signals.if_m10_0_a4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000110111100"
        )
    port map (
            in0 => \N__12629\,
            in1 => \N__15063\,
            in2 => \N__15426\,
            in3 => \N__12535\,
            lcout => \this_vga_signals.mult1_un54_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIK5K7M3_4_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15433\,
            in1 => \N__12073\,
            in2 => \_gnd_net_\,
            in3 => \N__12173\,
            lcout => \this_vga_signals.g0_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_x1_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100111100001"
        )
    port map (
            in0 => \N__13066\,
            in1 => \N__12851\,
            in2 => \N__12816\,
            in3 => \N__12967\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_1_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__11616\,
            in1 => \N__13187\,
            in2 => \N__12723\,
            in3 => \N__13651\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNISGOS_4_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000001"
        )
    port map (
            in0 => \N__13583\,
            in1 => \N__12999\,
            in2 => \N__11621\,
            in3 => \N__13799\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_fast_esr_RNISGOSZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIP2HP1_5_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__12713\,
            in1 => \_gnd_net_\,
            in2 => \N__11372\,
            in3 => \N__12731\,
            lcout => \this_vga_signals.vaddress_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_x0_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111001111000"
        )
    port map (
            in0 => \N__13067\,
            in1 => \N__12852\,
            in2 => \N__12815\,
            in3 => \N__12968\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un47_sum_axbxc3_1_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_ns_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12404\,
            in2 => \N__11369\,
            in3 => \N__11366\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_1\,
            ltout => \this_vga_signals.mult1_un47_sum_axbxc3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110100111100"
        )
    port map (
            in0 => \N__12804\,
            in1 => \N__11520\,
            in2 => \N__11360\,
            in3 => \N__11538\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011111011"
        )
    port map (
            in0 => \N__11539\,
            in1 => \N__12805\,
            in2 => \N__11525\,
            in3 => \N__12624\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_d_0_sqmuxa_i_0_0_a2_1_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11439\,
            in1 => \N__11715\,
            in2 => \_gnd_net_\,
            in3 => \N__11695\,
            lcout => \N_475\,
            ltout => \N_475_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m1_e_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000001010"
        )
    port map (
            in0 => \N__13146\,
            in1 => \N__12706\,
            in2 => \N__11501\,
            in3 => \N__11609\,
            lcout => \this_vga_signals.if_N_3_mux\,
            ltout => \this_vga_signals.if_N_3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axbxc1_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010110"
        )
    port map (
            in0 => \N__13065\,
            in1 => \N__12961\,
            in2 => \N__11498\,
            in3 => \N__12405\,
            lcout => \this_vga_signals.mult1_un47_sum_axb2_0\,
            ltout => \this_vga_signals.mult1_un47_sum_axb2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11480\,
            in2 => \N__11474\,
            in3 => \N__11471\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13111\,
            lcout => \this_vga_signals_M_vcounter_q_7_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24982\,
            ce => \N__15521\,
            sr => \N__15491\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12673\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals_M_vcounter_q_fast_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24982\,
            ce => \N__15521\,
            sr => \N__15491\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_x1_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__12705\,
            in1 => \N__11596\,
            in2 => \N__11443\,
            in3 => \N__11694\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0_1_0_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_x0_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__11595\,
            in1 => \N__12704\,
            in2 => \_gnd_net_\,
            in3 => \N__11435\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0_1_0_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axb2_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__14623\,
            in1 => \N__11848\,
            in2 => \_gnd_net_\,
            in3 => \N__11960\,
            lcout => \this_vga_signals.mult1_un61_sum_axb2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15537\,
            lcout => \this_vga_signals.M_vcounter_q_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24987\,
            ce => \N__15519\,
            sr => \N__15488\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_4_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15538\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24987\,
            ce => \N__15519\,
            sr => \N__15488\
        );

    \this_vga_signals.un4_lcounter_if_m5_0_1_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110111111001"
        )
    port map (
            in0 => \N__11699\,
            in1 => \N__13145\,
            in2 => \N__11732\,
            in3 => \N__13019\,
            lcout => \this_vga_signals.if_m5_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_1_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011100001"
        )
    port map (
            in0 => \N__13018\,
            in1 => \N__11727\,
            in2 => \N__13154\,
            in3 => \N__11697\,
            lcout => \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_axb1_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100010010110"
        )
    port map (
            in0 => \N__13791\,
            in1 => \N__13674\,
            in2 => \N__16615\,
            in3 => \N__13556\,
            lcout => \this_vga_signals.mult1_un40_sum_1_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101001"
        )
    port map (
            in0 => \N__13017\,
            in1 => \N__11728\,
            in2 => \N__13155\,
            in3 => \N__11698\,
            lcout => \this_vga_signals.N_370_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_axb1_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100010110110"
        )
    port map (
            in0 => \N__13790\,
            in1 => \N__13555\,
            in2 => \N__16614\,
            in3 => \N__13020\,
            lcout => \this_vga_signals.mult1_un40_sum_0_axb1_i\,
            ltout => \this_vga_signals.mult1_un40_sum_0_axb1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x1_1_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110010101"
        )
    port map (
            in0 => \N__13293\,
            in1 => \N__16588\,
            in2 => \N__11543\,
            in3 => \N__13792\,
            lcout => \this_vga_signals.mult1_un40_sum_m_x1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_axbxc2_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011010011100"
        )
    port map (
            in0 => \N__11768\,
            in1 => \N__11754\,
            in2 => \N__13314\,
            in3 => \N__13675\,
            lcout => \this_vga_signals.mult1_un40_sum1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_0_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010110011001"
        )
    port map (
            in0 => \N__13016\,
            in1 => \N__11726\,
            in2 => \N__13153\,
            in3 => \N__11696\,
            lcout => \this_vga_signals.N_330_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI8MCG1_9_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__13354\,
            in1 => \N__16612\,
            in2 => \_gnd_net_\,
            in3 => \N__14128\,
            lcout => \this_vga_signals.vsync_1_0_a2_6_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_m11_1_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__14270\,
            in1 => \N__13925\,
            in2 => \_gnd_net_\,
            in3 => \N__13207\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m11_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_m11_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011100010"
        )
    port map (
            in0 => \N__13926\,
            in1 => \N__13310\,
            in2 => \N__11648\,
            in3 => \N__11880\,
            lcout => this_vga_signals_un4_lcounter_if_i3_mux,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_26_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011011101"
        )
    port map (
            in0 => \N__16611\,
            in1 => \N__13800\,
            in2 => \_gnd_net_\,
            in3 => \N__13585\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_sbtinv_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16215\,
            lcout => \this_vga_signals.mult1_un47_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_2_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001000001"
        )
    port map (
            in0 => \N__14344\,
            in1 => \N__11916\,
            in2 => \N__15440\,
            in3 => \N__11969\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_0_x1_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000001100"
        )
    port map (
            in0 => \N__11899\,
            in1 => \N__11829\,
            in2 => \N__11633\,
            in3 => \N__11887\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_1_0_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_0_ns_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17434\,
            in2 => \N__11978\,
            in3 => \N__11929\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_2_1_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__15137\,
            in1 => \N__13924\,
            in2 => \_gnd_net_\,
            in3 => \N__13206\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_2_2_1\,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_2_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_sx_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110111110"
        )
    port map (
            in0 => \N__14343\,
            in1 => \N__15397\,
            in2 => \N__11963\,
            in3 => \N__11918\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14624\,
            in2 => \_gnd_net_\,
            in3 => \N__11953\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_4_tz_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__12942\,
            in1 => \N__11917\,
            in2 => \_gnd_net_\,
            in3 => \N__13847\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_2_4_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__11906\,
            in1 => \N__11900\,
            in2 => \_gnd_net_\,
            in3 => \N__11888\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_c2_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001101"
        )
    port map (
            in0 => \N__14531\,
            in1 => \N__14347\,
            in2 => \N__11861\,
            in3 => \N__11853\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_4_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11774\,
            lcout => \M_this_delay_clk_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25013\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_3_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11780\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25013\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_16_x1_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110000011100"
        )
    port map (
            in0 => \N__14573\,
            in1 => \N__14379\,
            in2 => \N__11995\,
            in3 => \N__12357\,
            lcout => \this_vga_signals.g0_16_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIU9QNGC_4_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15431\,
            in1 => \N__12299\,
            in2 => \_gnd_net_\,
            in3 => \N__12287\,
            lcout => \this_vga_signals.N_57_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__12587\,
            in1 => \N__12281\,
            in2 => \N__12476\,
            in3 => \N__12269\,
            lcout => \this_vga_signals.if_i3_mux_0_1\,
            ltout => \this_vga_signals.if_i3_mux_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_17_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000011111"
        )
    port map (
            in0 => \N__12235\,
            in1 => \N__14131\,
            in2 => \N__12257\,
            in3 => \N__14562\,
            lcout => \this_vga_signals.if_N_6_mux_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_2_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011010011100"
        )
    port map (
            in0 => \N__14563\,
            in1 => \N__12254\,
            in2 => \N__12248\,
            in3 => \N__12236\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_18_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__12227\,
            in1 => \N__12221\,
            in2 => \N__12215\,
            in3 => \N__12212\,
            lcout => \this_vga_signals.g2_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_7_i_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15428\,
            in2 => \N__12192\,
            in3 => \N__12061\,
            lcout => \this_vga_signals.N_5_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_10_1_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__14367\,
            in1 => \N__15141\,
            in2 => \N__15441\,
            in3 => \N__12551\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_10_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_10_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000011000000"
        )
    port map (
            in0 => \N__15143\,
            in1 => \N__12662\,
            in2 => \N__12647\,
            in3 => \N__12640\,
            lcout => \this_vga_signals.if_N_18_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI9OGF9_0_5_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15142\,
            in2 => \_gnd_net_\,
            in3 => \N__12552\,
            lcout => \this_vga_signals.m48_i_x4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g4_1_0_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011111111"
        )
    port map (
            in0 => \N__12553\,
            in1 => \N__15402\,
            in2 => \N__15154\,
            in3 => \N__14368\,
            lcout => \this_vga_signals.g4_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_0_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000111100"
        )
    port map (
            in0 => \N__12833\,
            in1 => \N__12902\,
            in2 => \N__12743\,
            in3 => \N__12410\,
            lcout => \this_vga_signals.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_cry_0_c_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17903\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \this_vga_signals.mult1_un68_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_cry_1_s_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14630\,
            in2 => \N__12890\,
            in3 => \N__12443\,
            lcout => \this_vga_signals.mult1_un68_sum_cry_1_s\,
            ltout => OPEN,
            carryin => \this_vga_signals.mult1_un68_sum_cry_0\,
            carryout => \this_vga_signals.mult1_un68_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_axb_3_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15639\,
            in1 => \N__12440\,
            in2 => \N__12866\,
            in3 => \N__12428\,
            lcout => \this_vga_signals.mult1_un75_sum_axb_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.mult1_un68_sum_cry_1\,
            carryout => \this_vga_signals.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_s_3_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12425\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12413\,
            lcout => \this_vga_signals.mult1_un68_sum_s_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_24_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110101111000"
        )
    port map (
            in0 => \N__12406\,
            in1 => \N__12829\,
            in2 => \N__13382\,
            in3 => \N__12901\,
            lcout => \this_vga_signals.N_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_4_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001111110"
        )
    port map (
            in0 => \N__13683\,
            in1 => \N__13578\,
            in2 => \N__13423\,
            in3 => \N__12857\,
            lcout => \this_vga_signals.g1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_sbtinv_3_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12886\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.mult1_un61_sum_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g6_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111011001001"
        )
    port map (
            in0 => \N__13655\,
            in1 => \N__13568\,
            in2 => \N__13424\,
            in3 => \N__12856\,
            lcout => \this_vga_signals.g6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI1K2D4_7_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__12914\,
            in1 => \N__14723\,
            in2 => \_gnd_net_\,
            in3 => \N__12818\,
            lcout => \M_this_vga_signals_address_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_27_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101100110"
        )
    port map (
            in0 => \N__15092\,
            in1 => \N__13656\,
            in2 => \_gnd_net_\,
            in3 => \N__13927\,
            lcout => \this_vga_signals.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0AS_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011001"
        )
    port map (
            in0 => \N__13798\,
            in1 => \N__12993\,
            in2 => \_gnd_net_\,
            in3 => \N__13567\,
            lcout => \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0ASZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_5_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13045\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24977\,
            ce => \N__15523\,
            sr => \N__15489\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12679\,
            lcout => \this_vga_signals.M_vcounter_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24977\,
            ce => \N__15523\,
            sr => \N__15489\
        );

    \this_vga_signals.M_vcounter_q_esr_6_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12680\,
            lcout => \this_vga_signals_M_vcounter_q_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24977\,
            ce => \N__15523\,
            sr => \N__15489\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010111011"
        )
    port map (
            in0 => \N__13773\,
            in1 => \N__13545\,
            in2 => \_gnd_net_\,
            in3 => \N__13159\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13178\,
            lcout => \this_vga_signals.M_vcounter_q_9_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24983\,
            ce => \N__15522\,
            sr => \N__15487\
        );

    \this_vga_signals.M_vcounter_q_esr_7_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13112\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24983\,
            ce => \N__15522\,
            sr => \N__15487\
        );

    \this_vga_signals.M_vcounter_q_esr_8_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13085\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24983\,
            ce => \N__15522\,
            sr => \N__15487\
        );

    \this_vga_signals.un5_vaddress_if_m1_0_0_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010010011"
        )
    port map (
            in0 => \N__13885\,
            in1 => \N__13544\,
            in2 => \N__13297\,
            in3 => \N__12992\,
            lcout => \this_vga_signals.vaddress_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13049\,
            lcout => \this_vga_signals.M_vcounter_q_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24983\,
            ce => \N__15522\,
            sr => \N__15487\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__13271\,
            in1 => \N__13884\,
            in2 => \_gnd_net_\,
            in3 => \N__12991\,
            lcout => \this_vga_signals.vaddress_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNINLU91_7_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001100"
        )
    port map (
            in0 => \N__12947\,
            in1 => \N__15984\,
            in2 => \N__13359\,
            in3 => \N__16085\,
            lcout => \this_vga_signals.M_this_vga_ramdac_en_i_o2_0_0\,
            ltout => \this_vga_signals.M_this_vga_ramdac_en_i_o2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIC1F54_7_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__14716\,
            in1 => \_gnd_net_\,
            in2 => \N__12905\,
            in3 => \N__13481\,
            lcout => \N_192_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13554\,
            in2 => \_gnd_net_\,
            in3 => \N__13788\,
            lcout => \N_183_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13292\,
            in2 => \_gnd_net_\,
            in3 => \N__13886\,
            lcout => \this_vga_signals.N_188_0_0_0\,
            ltout => \this_vga_signals.N_188_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_25_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110110111111"
        )
    port map (
            in0 => \N__13394\,
            in1 => \N__13676\,
            in2 => \N__13388\,
            in3 => \N__13789\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_c3_0_1_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_3_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010110000"
        )
    port map (
            in0 => \N__16638\,
            in1 => \N__13793\,
            in2 => \N__13385\,
            in3 => \N__13557\,
            lcout => \this_vga_signals.g1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_d_0_sqmuxa_i_0_0_o2_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__13677\,
            in1 => \N__16637\,
            in2 => \N__13358\,
            in3 => \N__15878\,
            lcout => \N_190_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIGBLD1_7_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13802\,
            in1 => \N__15152\,
            in2 => \N__13586\,
            in3 => \N__15339\,
            lcout => \N_275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x0_1_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010010"
        )
    port map (
            in0 => \N__16639\,
            in1 => \N__13801\,
            in2 => \N__13316\,
            in3 => \N__13232\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_m_x0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_1_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13226\,
            in2 => \N__13220\,
            in3 => \N__13217\,
            lcout => \this_vga_signals.mult1_un40_sum_m_ns_1\,
            ltout => \this_vga_signals.mult1_un40_sum_m_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_a3_1_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15151\,
            in2 => \N__13190\,
            in3 => \N__13923\,
            lcout => \this_vga_signals.if_N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_sbtinv_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16992\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.mult1_un54_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIL9AC2_7_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__13433\,
            in1 => \N__14957\,
            in2 => \N__16102\,
            in3 => \N__14828\,
            lcout => \N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_7_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__16640\,
            in1 => \N__13803\,
            in2 => \N__13701\,
            in3 => \N__13582\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_177_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI0T225_9_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__13439\,
            in1 => \N__14740\,
            in2 => \N__13490\,
            in3 => \N__13487\,
            lcout => \N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNICJJV_0_9_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__15877\,
            in1 => \N__15992\,
            in2 => \N__15791\,
            in3 => \N__16093\,
            lcout => \this_vga_signals.N_269_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNILVSO_6_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__15781\,
            in1 => \_gnd_net_\,
            in2 => \N__16342\,
            in3 => \N__16216\,
            lcout => \this_vga_signals.N_286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17002\,
            in1 => \N__14918\,
            in2 => \_gnd_net_\,
            in3 => \N__14909\,
            lcout => this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1,
            ltout => \this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_1_i_a0_2_9_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__17799\,
            in1 => \N__17888\,
            in2 => \N__13427\,
            in3 => \N__18099\,
            lcout => \this_ppu.sprites_addr_1_i_a0_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_o2_4_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__14687\,
            in1 => \N__14670\,
            in2 => \_gnd_net_\,
            in3 => \N__14645\,
            lcout => \this_vga_signals.N_185_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_o2_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__14672\,
            in1 => \N__14641\,
            in2 => \_gnd_net_\,
            in3 => \N__14685\,
            lcout => \N_175_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__14686\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14671\,
            lcout => \this_start_data_delay_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25006\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_sbtinv_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18100\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.mult1_un61_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axbxc1_0_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__14334\,
            in1 => \N__15236\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.vram_addr_1_i_7_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110000"
        )
    port map (
            in0 => \N__15790\,
            in1 => \N__15991\,
            in2 => \N__23843\,
            in3 => \N__16092\,
            lcout => \N_90_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m11_0_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14471\,
            in2 => \_gnd_net_\,
            in3 => \N__14255\,
            lcout => \N_184_0\,
            ltout => \N_184_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14067\,
            in2 => \N__13991\,
            in3 => \N__13966\,
            lcout => \this_vga_signals.N_272_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_0_c_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17803\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => \this_vga_signals.mult1_un75_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_1_c_inv_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14783\,
            in2 => \N__15661\,
            in3 => \N__17901\,
            lcout => \G_504\,
            ltout => OPEN,
            carryin => \this_vga_signals.mult1_un75_sum_cry_0\,
            carryout => \this_vga_signals.mult1_un75_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14762\,
            in2 => \N__14777\,
            in3 => \N__15657\,
            lcout => \G_503\,
            ltout => OPEN,
            carryin => \this_vga_signals.mult1_un75_sum_cry_1\,
            carryout => \this_vga_signals.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_s_3_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14756\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14747\,
            lcout => \this_vga_signals.N_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_m12_0_o2_381_4_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17897\,
            in1 => \N__16967\,
            in2 => \N__17807\,
            in3 => \N__16197\,
            lcout => OPEN,
            ltout => \this_ppu.M_m12_0_o2_381Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI38322_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__22384\,
            in1 => \N__18066\,
            in2 => \N__14744\,
            in3 => \N__15959\,
            lcout => OPEN,
            ltout => \this_ppu.M_m12_0_o2_381_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIIL1T5_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14945\,
            in1 => \N__14741\,
            in2 => \N__14726\,
            in3 => \N__14715\,
            lcout => \this_ppu.M_m12_0_o2_381_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNIPK611_0_6_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010111010111"
        )
    port map (
            in0 => \N__15938\,
            in1 => \N__15844\,
            in2 => \N__16063\,
            in3 => \N__14843\,
            lcout => \this_vga_signals.SUM_7_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_6_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15806\,
            lcout => \this_vga_signals.M_hcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24988\,
            ce => \N__15706\,
            sr => \N__17057\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNIPK611_6_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100101101100"
        )
    port map (
            in0 => \N__15845\,
            in1 => \N__14844\,
            in2 => \N__16064\,
            in3 => \N__15939\,
            lcout => \this_vga_signals.N_336_0\,
            ltout => \this_vga_signals.N_336_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_1_0_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000100010"
        )
    port map (
            in0 => \N__14845\,
            in1 => \N__16284\,
            in2 => \N__14849\,
            in3 => \N__14801\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_fast_esr_RNI21GQ_6_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__16168\,
            in1 => \_gnd_net_\,
            in2 => \N__16314\,
            in3 => \N__14846\,
            lcout => \this_vga_signals.N_287\,
            ltout => \this_vga_signals.N_287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111001010101"
        )
    port map (
            in0 => \N__14804\,
            in1 => \N__16170\,
            in2 => \N__14822\,
            in3 => \N__14819\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14890\,
            in2 => \N__14813\,
            in3 => \N__14863\,
            lcout => this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3,
            ltout => \this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_c3_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011011111"
        )
    port map (
            in0 => \N__16955\,
            in1 => \N__16171\,
            in2 => \N__14810\,
            in3 => \N__15685\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0_1\,
            ltout => \this_vga_signals.mult1_un68_sum_c3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_x0_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001001001011"
        )
    port map (
            in0 => \N__16291\,
            in1 => \N__16207\,
            in2 => \N__14807\,
            in3 => \N__16867\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010011111100"
        )
    port map (
            in0 => \N__14803\,
            in1 => \N__16285\,
            in2 => \N__15766\,
            in3 => \N__16167\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un54_sum_c3_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100110001"
        )
    port map (
            in0 => \N__16286\,
            in1 => \N__14862\,
            in2 => \N__15767\,
            in3 => \N__14802\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16290\,
            in2 => \N__14786\,
            in3 => \N__16169\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_1_i_2_1_9_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__16816\,
            in1 => \N__17979\,
            in2 => \_gnd_net_\,
            in3 => \N__18098\,
            lcout => \this_ppu.sprites_addr_1_i_2_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un54_sum_axb1_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101100000"
        )
    port map (
            in0 => \N__16065\,
            in1 => \N__15846\,
            in2 => \N__15983\,
            in3 => \N__15768\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_0\,
            ltout => \this_vga_signals.mult1_un54_sum_axb1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101111010010"
        )
    port map (
            in0 => \N__16202\,
            in1 => \N__16853\,
            in2 => \N__14930\,
            in3 => \N__16315\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110000111001"
        )
    port map (
            in0 => \N__16316\,
            in1 => \N__16233\,
            in2 => \N__16868\,
            in3 => \N__16203\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14927\,
            in2 => \N__14921\,
            in3 => \N__16762\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_1\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_ac0_1_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__18097\,
            in1 => \N__16987\,
            in2 => \N__14912\,
            in3 => \N__14908\,
            lcout => \this_vga_signals.mult1_un75_sum_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16860\,
            in1 => \N__16318\,
            in2 => \N__16240\,
            in3 => \N__16763\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_x1_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101111010100"
        )
    port map (
            in0 => \N__16317\,
            in1 => \N__16204\,
            in2 => \N__16869\,
            in3 => \N__14907\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_m1_0_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010011010"
        )
    port map (
            in0 => \N__16205\,
            in1 => \N__14894\,
            in2 => \N__14879\,
            in3 => \N__14867\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.pixel_clk_inferred_clock_RNO_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010001000010"
        )
    port map (
            in0 => \N__17801\,
            in1 => \N__15674\,
            in2 => \N__15665\,
            in3 => \N__17896\,
            lcout => \M_this_vga_signals_pixel_clk_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_4_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15542\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals_M_vcounter_q_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24969\,
            ce => \N__15524\,
            sr => \N__15486\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIFF6A3_5_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15458\,
            in1 => \N__15264\,
            in2 => \N__15203\,
            in3 => \N__15128\,
            lcout => \this_vga_signals.N_455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIGUM81_9_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14944\,
            in1 => \N__15875\,
            in2 => \_gnd_net_\,
            in3 => \N__15976\,
            lcout => \this_vga_signals.N_459\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__15876\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15961\,
            lcout => \this_vga_signals.N_404_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_d_0_sqmuxa_i_0_0_o2_0_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__15774\,
            in1 => \N__16309\,
            in2 => \_gnd_net_\,
            in3 => \N__16056\,
            lcout => \N_204_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIOT0S1_9_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17029\,
            in2 => \_gnd_net_\,
            in3 => \N__17086\,
            lcout => \this_vga_signals.N_517_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_1_i_a3_1_9_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__17788\,
            in1 => \N__17881\,
            in2 => \N__17802\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.N_4_0_1\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17148\,
            in1 => \N__18067\,
            in2 => \_gnd_net_\,
            in3 => \N__14933\,
            lcout => \this_vga_signals_M_hcounter_q_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_1_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_1_cry_2\,
            clk => \N__24984\,
            ce => 'H',
            sr => \N__17056\
        );

    \this_vga_signals.M_hcounter_q_3_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17140\,
            in1 => \N__16996\,
            in2 => \_gnd_net_\,
            in3 => \N__16115\,
            lcout => \this_vga_signals_M_hcounter_q_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_1_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_1_cry_3\,
            clk => \N__24984\,
            ce => 'H',
            sr => \N__17056\
        );

    \this_vga_signals.M_hcounter_q_4_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17149\,
            in1 => \N__16198\,
            in2 => \_gnd_net_\,
            in3 => \N__16112\,
            lcout => \this_vga_signals_M_hcounter_q_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_1_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_1_cry_4\,
            clk => \N__24984\,
            ce => 'H',
            sr => \N__17056\
        );

    \this_vga_signals.M_hcounter_q_5_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17141\,
            in1 => \N__16310\,
            in2 => \_gnd_net_\,
            in3 => \N__16109\,
            lcout => \this_vga_signals_M_hcounter_q_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_1_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_1_cry_5\,
            clk => \N__24984\,
            ce => 'H',
            sr => \N__17056\
        );

    \this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUF_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15765\,
            in2 => \_gnd_net_\,
            in3 => \N__16106\,
            lcout => \this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUFZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_1_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_7_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17142\,
            in1 => \N__16062\,
            in2 => \_gnd_net_\,
            in3 => \N__16007\,
            lcout => \this_vga_signals_M_hcounter_q_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_1_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_1_cry_7\,
            clk => \N__24984\,
            ce => 'H',
            sr => \N__17056\
        );

    \this_vga_signals.M_hcounter_q_8_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17150\,
            in1 => \N__15960\,
            in2 => \_gnd_net_\,
            in3 => \N__15896\,
            lcout => \this_vga_signals_M_hcounter_q_8\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_1_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_1_cry_8\,
            clk => \N__24984\,
            ce => 'H',
            sr => \N__17056\
        );

    \this_vga_signals.M_hcounter_q_esr_9_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15863\,
            in2 => \_gnd_net_\,
            in3 => \N__15893\,
            lcout => \this_vga_signals_M_hcounter_q_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24989\,
            ce => \N__15707\,
            sr => \N__17055\
        );

    \this_vga_signals.M_hcounter_q_esr_6_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15805\,
            lcout => \this_vga_signals_M_hcounter_q_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24989\,
            ce => \N__15707\,
            sr => \N__17055\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010111101"
        )
    port map (
            in0 => \N__16214\,
            in1 => \N__16764\,
            in2 => \N__17000\,
            in3 => \N__15686\,
            lcout => this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_1_i_0_0_9_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__23842\,
            in1 => \N__17953\,
            in2 => \N__16820\,
            in3 => \N__17928\,
            lcout => OPEN,
            ltout => \this_ppu.sprites_addr_1_i_0_0Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_1_i_0_2_9_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000010110000"
        )
    port map (
            in0 => \N__17929\,
            in1 => \N__16508\,
            in2 => \N__16499\,
            in3 => \N__16496\,
            lcout => OPEN,
            ltout => \this_ppu.sprites_addr_1_i_0_2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_1_i_0_9_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000010000"
        )
    port map (
            in0 => \N__16787\,
            in1 => \N__17954\,
            in2 => \N__16484\,
            in3 => \N__16793\,
            lcout => \N_138_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_ns_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16373\,
            in1 => \N__16367\,
            in2 => \_gnd_net_\,
            in3 => \N__16361\,
            lcout => if_generate_plus_mult1_un68_sum_axbxc3_ns,
            ltout => \if_generate_plus_mult1_un68_sum_axbxc3_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011001111001"
        )
    port map (
            in0 => \N__16355\,
            in1 => \N__16986\,
            in2 => \N__16349\,
            in3 => \N__16727\,
            lcout => this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0,
            ltout => \this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_m1_0_x1_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18245\,
            in1 => \N__17190\,
            in2 => \N__16346\,
            in3 => \N__17172\,
            lcout => \this_ppu.sprites_m1_0_xZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_m1_0_x0_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17171\,
            in1 => \N__18244\,
            in2 => \N__17194\,
            in3 => \N__17927\,
            lcout => \this_ppu.sprites_m1_0_xZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_m7_0_x4_0_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101111010010"
        )
    port map (
            in0 => \N__16870\,
            in1 => \N__16319\,
            in2 => \N__16241\,
            in3 => \N__16206\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_8_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_m7_0_m2_0_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110001110"
        )
    port map (
            in0 => \N__18082\,
            in1 => \N__16988\,
            in2 => \N__16730\,
            in3 => \N__16725\,
            lcout => this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_c3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_m7_0_o4_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__18083\,
            in1 => \N__16726\,
            in2 => \N__17902\,
            in3 => \N__17170\,
            lcout => \this_vga_signals.if_N_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_13_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010100110000"
        )
    port map (
            in0 => \N__25212\,
            in1 => \N__21242\,
            in2 => \N__21637\,
            in3 => \N__18911\,
            lcout => \M_this_internal_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25002\,
            ce => 'H',
            sr => \N__24739\
        );

    \M_this_internal_address_q_7_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010100110000"
        )
    port map (
            in0 => \N__25213\,
            in1 => \N__18776\,
            in2 => \N__21638\,
            in3 => \N__18305\,
            lcout => \M_this_internal_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25014\,
            ce => 'H',
            sr => \N__24734\
        );

    \CONSTANT_ONE_LUT4_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI4UBI1_9_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__16662\,
            in1 => \N__16712\,
            in2 => \_gnd_net_\,
            in3 => \N__16702\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNI4UBI1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_1_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__16703\,
            in1 => \N__16888\,
            in2 => \_gnd_net_\,
            in3 => \N__24785\,
            lcout => \this_pixel_clk_M_counter_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24970\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_RNIFKS8_0_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__16700\,
            in1 => \N__16887\,
            in2 => \_gnd_net_\,
            in3 => \N__24784\,
            lcout => \M_counter_q_RNIFKS8_0\,
            ltout => \M_counter_q_RNIFKS8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.G_210_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16706\,
            in3 => \N__16701\,
            lcout => \this_vga_signals.GZ0Z_210\,
            ltout => \this_vga_signals.GZ0Z_210_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIRV75_9_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__16688\,
            in1 => \N__16661\,
            in2 => \N__16646\,
            in3 => \N__16641\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNIIRV75Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_0_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16889\,
            lcout => \this_pixel_clk.M_counter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24974\,
            ce => 'H',
            sr => \N__24742\
        );

    \this_sprites_ram.mem_radreg_11_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__23858\,
            in1 => \N__16778\,
            in2 => \N__16739\,
            in3 => \N__18287\,
            lcout => \this_sprites_ram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIG0MN6_7_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__23857\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16874\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__17200\,
            in1 => \N__17173\,
            in2 => \_gnd_net_\,
            in3 => \N__18247\,
            lcout => if_generate_plus_mult1_un75_sum_axbxc3,
            ltout => \if_generate_plus_mult1_un75_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un5_sprites_addr_1_ac0_1_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001000"
        )
    port map (
            in0 => \N__23830\,
            in1 => \N__17966\,
            in2 => \N__16826\,
            in3 => \N__17933\,
            lcout => \this_ppu.un5_sprites_addr_1_c2\,
            ltout => \this_ppu.un5_sprites_addr_1_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un5_sprites_addr_1_ac0_5_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__16773\,
            in1 => \_gnd_net_\,
            in2 => \N__16823\,
            in3 => \N__18249\,
            lcout => \this_ppu.un5_sprites_addr_1_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_1_i_8_tz_9_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111010101110"
        )
    port map (
            in0 => \N__17996\,
            in1 => \N__16815\,
            in2 => \N__18093\,
            in3 => \N__17935\,
            lcout => \this_ppu.sprites_addr_1_i_7_tz_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_1_i_a7_9_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__17934\,
            in1 => \N__18062\,
            in2 => \_gnd_net_\,
            in3 => \N__17995\,
            lcout => \this_ppu.sprites_addr_1_i_a7Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un5_sprites_addr_1_axbxc3_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000001000000"
        )
    port map (
            in0 => \N__18250\,
            in1 => \N__18268\,
            in2 => \N__23856\,
            in3 => \N__16774\,
            lcout => \this_ppu.un5_sprites_addr1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un82_sum_axb1_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17201\,
            in1 => \N__17174\,
            in2 => \N__18107\,
            in3 => \N__18248\,
            lcout => this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axb1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_1_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__17775\,
            in1 => \N__17119\,
            in2 => \_gnd_net_\,
            in3 => \N__17871\,
            lcout => \this_vga_signals_M_hcounter_q_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24990\,
            ce => 'H',
            sr => \N__17054\
        );

    \this_vga_signals.M_hcounter_q_0_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17118\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17774\,
            lcout => \this_vga_signals_M_hcounter_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24990\,
            ce => 'H',
            sr => \N__17054\
        );

    \this_vga_signals.un3_haddress_if_m7_0_m2_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100100111"
        )
    port map (
            in0 => \N__17001\,
            in1 => \N__16916\,
            in2 => \N__18101\,
            in3 => \N__18246\,
            lcout => this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3,
            ltout => \this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_m1_0_ns_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16910\,
            in2 => \N__16904\,
            in3 => \N__16901\,
            lcout => \this_ppu_sprites_N_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_0_2_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__21212\,
            in1 => \N__18471\,
            in2 => \N__22759\,
            in3 => \N__21975\,
            lcout => \M_this_internal_address_q_3_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_0_9_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100100111"
        )
    port map (
            in0 => \N__21977\,
            in1 => \N__22754\,
            in2 => \N__19093\,
            in3 => \N__21214\,
            lcout => \M_this_internal_address_q_3_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_0_8_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011011111"
        )
    port map (
            in0 => \N__21976\,
            in1 => \N__21213\,
            in2 => \N__21035\,
            in3 => \N__19215\,
            lcout => \M_this_internal_address_q_3_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_2_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011101000100"
        )
    port map (
            in0 => \N__16895\,
            in1 => \N__21601\,
            in2 => \N__25252\,
            in3 => \N__18452\,
            lcout => \M_this_internal_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24997\,
            ce => 'H',
            sr => \N__24737\
        );

    \M_this_internal_address_q_9_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__17225\,
            in1 => \N__25215\,
            in2 => \N__21626\,
            in3 => \N__19067\,
            lcout => \M_this_internal_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24997\,
            ce => 'H',
            sr => \N__24737\
        );

    \M_this_internal_address_q_RNO_0_3_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__21224\,
            in1 => \N__18342\,
            in2 => \N__23198\,
            in3 => \N__22021\,
            lcout => OPEN,
            ltout => \M_this_internal_address_q_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_3_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101100001010"
        )
    port map (
            in0 => \N__21602\,
            in1 => \N__25214\,
            in2 => \N__17219\,
            in3 => \N__18323\,
            lcout => \M_this_internal_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24997\,
            ce => 'H',
            sr => \N__24737\
        );

    \M_this_internal_address_q_8_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000110000"
        )
    port map (
            in0 => \N__21225\,
            in1 => \N__17216\,
            in2 => \N__21625\,
            in3 => \N__19196\,
            lcout => \M_this_internal_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24997\,
            ce => 'H',
            sr => \N__24737\
        );

    \M_this_state_q_RNI20CE_0_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25197\,
            in2 => \_gnd_net_\,
            in3 => \N__24798\,
            lcout => \M_this_state_q_RNI20CEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_0_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19556\,
            in2 => \N__23545\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \un1_M_this_data_count_q_cry_0\,
            clk => \N__25007\,
            ce => 'H',
            sr => \N__17696\
        );

    \M_this_data_count_q_1_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23522\,
            in2 => \N__19388\,
            in3 => \N__17210\,
            lcout => \M_this_data_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_0\,
            carryout => \un1_M_this_data_count_q_cry_1\,
            clk => \N__25007\,
            ce => 'H',
            sr => \N__17696\
        );

    \M_this_data_count_q_2_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19415\,
            in2 => \N__23546\,
            in3 => \N__17207\,
            lcout => \M_this_data_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_1\,
            carryout => \un1_M_this_data_count_q_cry_2\,
            clk => \N__25007\,
            ce => 'H',
            sr => \N__17696\
        );

    \M_this_data_count_q_3_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23526\,
            in2 => \N__19430\,
            in3 => \N__17204\,
            lcout => \M_this_data_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_2\,
            carryout => \un1_M_this_data_count_q_cry_3\,
            clk => \N__25007\,
            ce => 'H',
            sr => \N__17696\
        );

    \M_this_data_count_q_4_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19442\,
            in2 => \N__23547\,
            in3 => \N__17252\,
            lcout => \M_this_data_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_3\,
            carryout => \un1_M_this_data_count_q_cry_4\,
            clk => \N__25007\,
            ce => 'H',
            sr => \N__17696\
        );

    \M_this_data_count_q_5_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23530\,
            in2 => \N__19475\,
            in3 => \N__17249\,
            lcout => \M_this_data_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_4\,
            carryout => \un1_M_this_data_count_q_cry_5\,
            clk => \N__25007\,
            ce => 'H',
            sr => \N__17696\
        );

    \M_this_data_count_q_6_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19487\,
            in2 => \N__23548\,
            in3 => \N__17246\,
            lcout => \M_this_data_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_5\,
            carryout => \un1_M_this_data_count_q_cry_6\,
            clk => \N__25007\,
            ce => 'H',
            sr => \N__17696\
        );

    \M_this_data_count_q_7_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23534\,
            in2 => \N__19460\,
            in3 => \N__17243\,
            lcout => \M_this_data_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_6\,
            carryout => \un1_M_this_data_count_q_cry_7\,
            clk => \N__25007\,
            ce => 'H',
            sr => \N__17696\
        );

    \M_this_data_count_q_8_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19513\,
            in2 => \N__23540\,
            in3 => \N__17240\,
            lcout => \M_this_data_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => \un1_M_this_data_count_q_cry_8\,
            clk => \N__25015\,
            ce => 'H',
            sr => \N__17695\
        );

    \M_this_data_count_q_9_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23505\,
            in2 => \N__19529\,
            in3 => \N__17237\,
            lcout => \M_this_data_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_8\,
            carryout => \un1_M_this_data_count_q_cry_9\,
            clk => \N__25015\,
            ce => 'H',
            sr => \N__17695\
        );

    \M_this_data_count_q_10_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19402\,
            in2 => \N__23541\,
            in3 => \N__17234\,
            lcout => \M_this_data_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_9\,
            carryout => \un1_M_this_data_count_q_cry_10\,
            clk => \N__25015\,
            ce => 'H',
            sr => \N__17695\
        );

    \M_this_data_count_q_11_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23509\,
            in2 => \N__19544\,
            in3 => \N__17231\,
            lcout => \M_this_data_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_10\,
            carryout => \un1_M_this_data_count_q_cry_11\,
            clk => \N__25015\,
            ce => 'H',
            sr => \N__17695\
        );

    \M_this_data_count_q_12_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19499\,
            in2 => \N__23542\,
            in3 => \N__17228\,
            lcout => \M_this_data_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_11\,
            carryout => \un1_M_this_data_count_q_cry_12\,
            clk => \N__25015\,
            ce => 'H',
            sr => \N__17695\
        );

    \un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17346\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_12\,
            carryout => \un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17348\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO\,
            carryout => \un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17347\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO\,
            carryout => \un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_13_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__25251\,
            in1 => \N__23543\,
            in2 => \N__19571\,
            in3 => \N__17318\,
            lcout => \M_this_data_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25017\,
            ce => 'H',
            sr => \N__24731\
        );

    \this_reset_cond.M_stage_q_3_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__19352\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17315\,
            lcout => \M_this_state_q_nss_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24965\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19351\,
            in2 => \_gnd_net_\,
            in3 => \N__19319\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24965\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_13_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__18286\,
            in1 => \N__17273\,
            in2 => \N__17302\,
            in3 => \N__17264\,
            lcout => \this_sprites_ram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24973\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_12_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__17272\,
            in1 => \N__17263\,
            in2 => \_gnd_net_\,
            in3 => \N__18285\,
            lcout => \this_sprites_ram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24973\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_ac0_3_0_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101110001001"
        )
    port map (
            in0 => \N__17870\,
            in1 => \N__17714\,
            in2 => \N__17795\,
            in3 => \N__19755\,
            lcout => this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_c3_0,
            ltout => \this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__19756\,
            in1 => \_gnd_net_\,
            in2 => \N__18290\,
            in3 => \N__23691\,
            lcout => if_generate_plus_mult1_un89_sum_axbxc3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_m6_0_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101101110110"
        )
    port map (
            in0 => \N__17869\,
            in1 => \N__17712\,
            in2 => \N__17800\,
            in3 => \N__19754\,
            lcout => OPEN,
            ltout => \this_ppu.sprites_N_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_m7_0_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18272\,
            in3 => \N__23690\,
            lcout => OPEN,
            ltout => \this_ppu.sprites_m7Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.N_140_i_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010100010"
        )
    port map (
            in0 => \N__23859\,
            in1 => \N__18269\,
            in2 => \N__18257\,
            in3 => \N__18254\,
            lcout => \N_140_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010000101011"
        )
    port map (
            in0 => \N__17952\,
            in1 => \N__18105\,
            in2 => \N__17889\,
            in3 => \N__17994\,
            lcout => this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_m1_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17965\,
            in1 => \N__17951\,
            in2 => \_gnd_net_\,
            in3 => \N__17936\,
            lcout => OPEN,
            ltout => \this_ppu.sprites_mZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_m5_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111101000"
        )
    port map (
            in0 => \N__17865\,
            in1 => \N__17773\,
            in2 => \N__17717\,
            in3 => \N__17713\,
            lcout => \this_ppu.sprites_N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_0_10_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011101010101"
        )
    port map (
            in0 => \N__18951\,
            in1 => \N__21215\,
            in2 => \N__23194\,
            in3 => \N__22003\,
            lcout => OPEN,
            ltout => \M_this_internal_address_q_3_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_10_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001110100001100"
        )
    port map (
            in0 => \N__25152\,
            in1 => \N__21583\,
            in2 => \N__17699\,
            in3 => \N__18932\,
            lcout => \M_this_internal_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24985\,
            ce => 'H',
            sr => \N__24736\
        );

    \M_this_internal_address_q_RNO_1_0_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20011\,
            in2 => \N__20141\,
            in3 => \N__20140\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_21_0_\,
            carryout => \un1_M_this_internal_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_1_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19861\,
            in2 => \_gnd_net_\,
            in3 => \N__18578\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_0\,
            carryout => \un1_M_this_internal_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_2_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18472\,
            in2 => \_gnd_net_\,
            in3 => \N__18446\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_1\,
            carryout => \un1_M_this_internal_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_3_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18346\,
            in2 => \_gnd_net_\,
            in3 => \N__18317\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_2\,
            carryout => \un1_M_this_internal_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_4_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20269\,
            in2 => \_gnd_net_\,
            in3 => \N__18314\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_3\,
            carryout => \un1_M_this_internal_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_5_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21406\,
            in2 => \_gnd_net_\,
            in3 => \N__18311\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_4\,
            carryout => \un1_M_this_internal_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_6_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21279\,
            in2 => \_gnd_net_\,
            in3 => \N__18308\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_5\,
            carryout => \un1_M_this_internal_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_7_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18808\,
            in2 => \_gnd_net_\,
            in3 => \N__18293\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_6\,
            carryout => \un1_M_this_internal_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_8_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19216\,
            in2 => \_gnd_net_\,
            in3 => \N__19190\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_16_22_0_\,
            carryout => \un1_M_this_internal_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_9_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19086\,
            in2 => \_gnd_net_\,
            in3 => \N__19061\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_8\,
            carryout => \un1_M_this_internal_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_10_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18958\,
            in2 => \_gnd_net_\,
            in3 => \N__18923\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_9\,
            carryout => \un1_M_this_internal_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_11_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24079\,
            in2 => \_gnd_net_\,
            in3 => \N__18920\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_10\,
            carryout => \un1_M_this_internal_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_12_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24169\,
            in2 => \_gnd_net_\,
            in3 => \N__18917\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_internal_address_q_cry_11\,
            carryout => \un1_M_this_internal_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_1_13_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24030\,
            in2 => \_gnd_net_\,
            in3 => \N__18914\,
            lcout => \M_this_internal_address_q_RNO_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_0_7_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100110011"
        )
    port map (
            in0 => \N__21233\,
            in1 => \N__18801\,
            in2 => \N__20874\,
            in3 => \N__22028\,
            lcout => \M_this_internal_address_q_3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_0_0_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__21232\,
            in1 => \N__20004\,
            in2 => \N__20873\,
            in3 => \N__22027\,
            lcout => \M_this_internal_address_q_3_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \N_235_0_sbtinv_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20192\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_235_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIEOD9_13_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__19567\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19555\,
            lcout => \M_this_state_q_srsts_0_a2_1_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIAVRI_11_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19540\,
            in1 => \N__19525\,
            in2 => \N__19514\,
            in3 => \N__19498\,
            lcout => \M_this_state_q_srsts_0_a2_1_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIAQQL_4_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19486\,
            in1 => \N__19471\,
            in2 => \N__19459\,
            in3 => \N__19441\,
            lcout => \M_this_state_q_srsts_0_a2_1_9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIBTAK_10_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19426\,
            in1 => \N__19414\,
            in2 => \N__19403\,
            in3 => \N__19384\,
            lcout => OPEN,
            ltout => \M_this_state_q_srsts_0_a2_1_8_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIDFF62_10_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19373\,
            in1 => \N__19367\,
            in2 => \N__19361\,
            in3 => \N__19358\,
            lcout => \N_240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19344\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19345\,
            in2 => \_gnd_net_\,
            in3 => \N__19325\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_i_i_a2_0_3_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20448\,
            in2 => \_gnd_net_\,
            in3 => \N__22022\,
            lcout => \N_476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_i_o4_1_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__19799\,
            in1 => \N__20626\,
            in2 => \_gnd_net_\,
            in3 => \N__19828\,
            lcout => \this_vga_signals.N_224_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_addr_1_i_7_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__23692\,
            in1 => \N__19766\,
            in2 => \N__23861\,
            in3 => \N__19760\,
            lcout => \N_134_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_1_4_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__20487\,
            in1 => \N__19628\,
            in2 => \N__20549\,
            in3 => \N__19613\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_i_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_1_4_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__23430\,
            in1 => \N__20449\,
            in2 => \N__20589\,
            in3 => \N__24790\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_4\,
            ltout => \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_4_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011111111"
        )
    port map (
            in0 => \N__24599\,
            in1 => \N__20600\,
            in2 => \N__19622\,
            in3 => \N__19619\,
            lcout => \M_this_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24991\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_0_4_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__19821\,
            in1 => \N__20147\,
            in2 => \N__19802\,
            in3 => \N__24788\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_i_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_1_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__24789\,
            in1 => \N__25153\,
            in2 => \N__19607\,
            in3 => \N__23431\,
            lcout => \M_this_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_0_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19598\,
            lcout => \M_this_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.port_nmib_i_o2_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__23407\,
            in1 => \N__19794\,
            in2 => \_gnd_net_\,
            in3 => \N__20447\,
            lcout => \N_235_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_0_1_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__21223\,
            in1 => \N__19860\,
            in2 => \N__21043\,
            in3 => \N__22042\,
            lcout => \M_this_internal_address_q_3_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_a2_2_4_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__22041\,
            in1 => \N__20167\,
            in2 => \N__25196\,
            in3 => \N__24786\,
            lcout => \this_vga_signals.N_319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un19_i_i_i_a2_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__19798\,
            in1 => \N__22072\,
            in2 => \N__20591\,
            in3 => \N__22040\,
            lcout => un19_i_i_i_a2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_11_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__20390\,
            in1 => \N__25159\,
            in2 => \N__21636\,
            in3 => \N__20126\,
            lcout => \M_this_internal_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25003\,
            ce => 'H',
            sr => \N__24735\
        );

    \M_this_internal_address_q_0_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001011100"
        )
    port map (
            in0 => \N__20120\,
            in1 => \N__20114\,
            in2 => \N__21633\,
            in3 => \N__25161\,
            lcout => \M_this_internal_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25008\,
            ce => 'H',
            sr => \N__24732\
        );

    \M_this_internal_address_q_1_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__19985\,
            in1 => \N__25160\,
            in2 => \N__21634\,
            in3 => \N__19976\,
            lcout => \M_this_internal_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25008\,
            ce => 'H',
            sr => \N__24732\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_1_a2_1_0_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19835\,
            in2 => \_gnd_net_\,
            in3 => \N__21114\,
            lcout => \this_vga_signals.N_479\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_i_a2_2_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__20446\,
            in1 => \N__19800\,
            in2 => \N__20630\,
            in3 => \N__19829\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_343_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_2_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__19801\,
            in1 => \N__22053\,
            in2 => \N__19769\,
            in3 => \N__24799\,
            lcout => \M_this_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24996\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_a4_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__21113\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20445\,
            lcout => \this_vga_signals.N_483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_3_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20450\,
            in2 => \_gnd_net_\,
            in3 => \N__22031\,
            lcout => \M_this_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24998\,
            ce => 'H',
            sr => \N__24741\
        );

    \M_this_internal_address_q_5_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000110000"
        )
    port map (
            in0 => \N__21196\,
            in1 => \N__21380\,
            in2 => \N__21566\,
            in3 => \N__20417\,
            lcout => \M_this_internal_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25004\,
            ce => 'H',
            sr => \N__24740\
        );

    \M_this_internal_address_q_6_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000001100"
        )
    port map (
            in0 => \N__21197\,
            in1 => \N__21541\,
            in2 => \N__21251\,
            in3 => \N__20408\,
            lcout => \M_this_internal_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25004\,
            ce => 'H',
            sr => \N__24740\
        );

    \M_this_internal_address_q_12_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__21122\,
            in1 => \N__25220\,
            in2 => \N__21612\,
            in3 => \N__20399\,
            lcout => \M_this_internal_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25009\,
            ce => 'H',
            sr => \N__24738\
        );

    \M_this_internal_address_q_RNO_0_4_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110110011"
        )
    port map (
            in0 => \N__22036\,
            in1 => \N__20259\,
            in2 => \N__21231\,
            in3 => \N__20823\,
            lcout => \M_this_internal_address_q_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_0_11_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011101010101"
        )
    port map (
            in0 => \N__24080\,
            in1 => \N__21219\,
            in2 => \N__20827\,
            in3 => \N__22035\,
            lcout => \M_this_internal_address_q_3_ns_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_4_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__20384\,
            in1 => \N__25219\,
            in2 => \N__21635\,
            in3 => \N__20378\,
            lcout => \M_this_internal_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25018\,
            ce => 'H',
            sr => \N__24733\
        );

    \this_vga_signals.M_this_vram_write_data_0_i_1_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__23500\,
            in1 => \N__21752\,
            in2 => \N__21042\,
            in3 => \N__22404\,
            lcout => \M_this_vram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_o4_4_4_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__20699\,
            in1 => \N__20678\,
            in2 => \N__20660\,
            in3 => \N__20625\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_i_o4_4Z0Z_4\,
            ltout => \this_vga_signals.M_this_state_q_srsts_0_i_o4_4Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_2_7_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__24595\,
            in1 => \N__20590\,
            in2 => \N__20561\,
            in3 => \N__24791\,
            lcout => \this_vga_signals.N_490\,
            ltout => \this_vga_signals.N_490_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_0_7_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100000"
        )
    port map (
            in0 => \N__20545\,
            in1 => \N__20507\,
            in2 => \N__20558\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_386_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_7_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__21116\,
            in1 => \N__22052\,
            in2 => \N__20555\,
            in3 => \N__24792\,
            lcout => \M_this_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24999\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_internal_address_q_3_ss0_i_a3_0_a2_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21660\,
            in2 => \_gnd_net_\,
            in3 => \N__25154\,
            lcout => \N_355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_6_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__24794\,
            in1 => \N__21649\,
            in2 => \_gnd_net_\,
            in3 => \N__22030\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_387_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_6_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__20459\,
            in1 => \N__20506\,
            in2 => \N__20552\,
            in3 => \N__20544\,
            lcout => \M_this_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25005\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_5_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__21661\,
            in1 => \N__22029\,
            in2 => \_gnd_net_\,
            in3 => \N__24793\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_391_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_5_LC_19_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__20543\,
            in1 => \N__20505\,
            in2 => \N__20462\,
            in3 => \N__20458\,
            lcout => \M_this_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25005\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_internal_address_q_3s2_i_0_LC_19_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010000"
        )
    port map (
            in0 => \N__25155\,
            in1 => \_gnd_net_\,
            in2 => \N__21665\,
            in3 => \N__21650\,
            lcout => \N_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_0_5_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__21170\,
            in1 => \N__21399\,
            in2 => \N__21091\,
            in3 => \N__22044\,
            lcout => \M_this_internal_address_q_3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_0_6_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011110001111"
        )
    port map (
            in0 => \N__22045\,
            in1 => \N__21171\,
            in2 => \N__21280\,
            in3 => \N__22711\,
            lcout => \M_this_internal_address_q_3_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_0_13_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011101010101"
        )
    port map (
            in0 => \N__23988\,
            in1 => \N__21169\,
            in2 => \N__22712\,
            in3 => \N__22043\,
            lcout => \M_this_internal_address_q_3_ns_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_internal_address_q_RNO_0_12_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011011111"
        )
    port map (
            in0 => \N__22054\,
            in1 => \N__21198\,
            in2 => \N__21092\,
            in3 => \N__24160\,
            lcout => \M_this_internal_address_q_3_ns_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_1_a2_2_0_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22026\,
            in2 => \_gnd_net_\,
            in3 => \N__21115\,
            lcout => \this_vga_signals.N_481\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_1_i_1_LC_21_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__21078\,
            in1 => \N__22779\,
            in2 => \N__21047\,
            in3 => \N__24344\,
            lcout => \M_this_sprites_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_1_i_0_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__20881\,
            in1 => \N__22788\,
            in2 => \N__20831\,
            in3 => \N__24354\,
            lcout => \M_this_sprites_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_vram_write_data_0_i_2_LC_22_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__23536\,
            in1 => \N__21761\,
            in2 => \N__22766\,
            in3 => \N__22411\,
            lcout => \M_this_vram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_22_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__22270\,
            in1 => \N__22124\,
            in2 => \N__22212\,
            in3 => \N__21671\,
            lcout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_23_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22910\,
            in1 => \N__21800\,
            in2 => \_gnd_net_\,
            in3 => \N__21779\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_23_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__22211\,
            in1 => \N__22268\,
            in2 => \N__21767\,
            in3 => \N__22544\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_23_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__22484\,
            in1 => \N__22269\,
            in2 => \N__21764\,
            in3 => \N__22610\,
            lcout => \M_this_sprites_ram_read_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_23_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__22298\,
            in1 => \N__22421\,
            in2 => \N__22217\,
            in3 => \N__22577\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_23_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__22299\,
            in1 => \N__22454\,
            in2 => \N__21755\,
            in3 => \N__21710\,
            lcout => \M_this_sprites_ram_read_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_23_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22907\,
            in1 => \N__21743\,
            in2 => \_gnd_net_\,
            in3 => \N__21728\,
            lcout => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22855\,
            in1 => \N__21704\,
            in2 => \_gnd_net_\,
            in3 => \N__21692\,
            lcout => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001100100011"
        )
    port map (
            in0 => \N__23219\,
            in1 => \N__22157\,
            in2 => \N__22300\,
            in3 => \N__23009\,
            lcout => OPEN,
            ltout => \M_this_sprites_ram_read_data_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_vram_write_data_0_i_3_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__23193\,
            in1 => \N__23470\,
            in2 => \N__22415\,
            in3 => \N__22412\,
            lcout => \M_this_vram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__22285\,
            in1 => \N__22949\,
            in2 => \N__22213\,
            in3 => \N__22982\,
            lcout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22895\,
            in1 => \N__22151\,
            in2 => \_gnd_net_\,
            in3 => \N__22139\,
            lcout => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22118\,
            in1 => \N__22106\,
            in2 => \_gnd_net_\,
            in3 => \N__22898\,
            lcout => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_LC_23_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22073\,
            in2 => \_gnd_net_\,
            in3 => \N__22055\,
            lcout => \N_24_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_7_0_wclke_3_LC_23_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24173\,
            in1 => \N__24094\,
            in2 => \N__24041\,
            in3 => \N__23918\,
            lcout => \this_sprites_ram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__24207\,
            in1 => \N__24130\,
            in2 => \N__24051\,
            in3 => \N__23941\,
            lcout => \this_sprites_ram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__23942\,
            in1 => \N__24034\,
            in2 => \N__24134\,
            in3 => \N__24208\,
            lcout => \this_sprites_ram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__24129\,
            in1 => \N__24209\,
            in2 => \N__24052\,
            in3 => \N__23940\,
            lcout => \this_sprites_ram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_24_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22637\,
            in1 => \N__22622\,
            in2 => \_gnd_net_\,
            in3 => \N__22916\,
            lcout => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_24_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22914\,
            in1 => \N__22604\,
            in2 => \_gnd_net_\,
            in3 => \N__22592\,
            lcout => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_24_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22915\,
            in1 => \N__22571\,
            in2 => \_gnd_net_\,
            in3 => \N__22559\,
            lcout => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__24206\,
            in1 => \N__24120\,
            in2 => \N__24053\,
            in3 => \N__23931\,
            lcout => \this_sprites_ram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_24_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22906\,
            in1 => \N__22514\,
            in2 => \_gnd_net_\,
            in3 => \N__22496\,
            lcout => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_24_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22478\,
            in1 => \N__22460\,
            in2 => \_gnd_net_\,
            in3 => \N__22905\,
            lcout => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_24_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22904\,
            in1 => \N__22448\,
            in2 => \_gnd_net_\,
            in3 => \N__22433\,
            lcout => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_24_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22909\,
            in1 => \N__23246\,
            in2 => \_gnd_net_\,
            in3 => \N__23228\,
            lcout => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24194\,
            in1 => \N__24103\,
            in2 => \N__24056\,
            in3 => \N__23919\,
            lcout => \this_sprites_ram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_1_i_3_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__23192\,
            in1 => \N__22795\,
            in2 => \N__23129\,
            in3 => \N__24359\,
            lcout => \M_this_sprites_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_24_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23036\,
            in1 => \N__23024\,
            in2 => \_gnd_net_\,
            in3 => \N__22908\,
            lcout => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_24_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23003\,
            in1 => \N__22894\,
            in2 => \_gnd_net_\,
            in3 => \N__22988\,
            lcout => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22896\,
            in1 => \N__22976\,
            in2 => \_gnd_net_\,
            in3 => \N__22964\,
            lcout => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22943\,
            in1 => \N__22928\,
            in2 => \_gnd_net_\,
            in3 => \N__22897\,
            lcout => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_1_i_2_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__22799\,
            in1 => \N__22755\,
            in2 => \N__22699\,
            in3 => \N__24358\,
            lcout => \M_this_sprites_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__24174\,
            in1 => \N__24095\,
            in2 => \N__24055\,
            in3 => \N__23929\,
            lcout => \this_sprites_ram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__24175\,
            in1 => \N__24096\,
            in2 => \N__24054\,
            in3 => \N__23930\,
            lcout => \this_sprites_ram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.sprites_m7_LC_24_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__23855\,
            in1 => \N__23702\,
            in2 => \_gnd_net_\,
            in3 => \N__23669\,
            lcout => sprites_m7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_0_LC_31_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25253\,
            in1 => \N__23347\,
            in2 => \N__23544\,
            in3 => \N__23535\,
            lcout => \M_this_external_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_31_23_0_\,
            carryout => \un1_M_this_external_address_q_cry_0\,
            clk => \N__25034\,
            ce => 'H',
            sr => \N__24745\
        );

    \M_this_external_address_q_1_LC_31_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25261\,
            in1 => \N__23329\,
            in2 => \_gnd_net_\,
            in3 => \N__23318\,
            lcout => \M_this_external_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_0\,
            carryout => \un1_M_this_external_address_q_cry_1\,
            clk => \N__25034\,
            ce => 'H',
            sr => \N__24745\
        );

    \M_this_external_address_q_2_LC_31_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25254\,
            in1 => \N__23299\,
            in2 => \_gnd_net_\,
            in3 => \N__23288\,
            lcout => \M_this_external_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_1\,
            carryout => \un1_M_this_external_address_q_cry_2\,
            clk => \N__25034\,
            ce => 'H',
            sr => \N__24745\
        );

    \M_this_external_address_q_3_LC_31_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25262\,
            in1 => \N__23275\,
            in2 => \_gnd_net_\,
            in3 => \N__23264\,
            lcout => \M_this_external_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_2\,
            carryout => \un1_M_this_external_address_q_cry_3\,
            clk => \N__25034\,
            ce => 'H',
            sr => \N__24745\
        );

    \M_this_external_address_q_4_LC_31_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25255\,
            in1 => \N__23257\,
            in2 => \_gnd_net_\,
            in3 => \N__24566\,
            lcout => \M_this_external_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_3\,
            carryout => \un1_M_this_external_address_q_cry_4\,
            clk => \N__25034\,
            ce => 'H',
            sr => \N__24745\
        );

    \M_this_external_address_q_5_LC_31_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25263\,
            in1 => \N__24556\,
            in2 => \_gnd_net_\,
            in3 => \N__24545\,
            lcout => \M_this_external_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_4\,
            carryout => \un1_M_this_external_address_q_cry_5\,
            clk => \N__25034\,
            ce => 'H',
            sr => \N__24745\
        );

    \M_this_external_address_q_6_LC_31_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25256\,
            in1 => \N__24535\,
            in2 => \_gnd_net_\,
            in3 => \N__24524\,
            lcout => \M_this_external_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_5\,
            carryout => \un1_M_this_external_address_q_cry_6\,
            clk => \N__25034\,
            ce => 'H',
            sr => \N__24745\
        );

    \M_this_external_address_q_7_LC_31_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25264\,
            in1 => \N__24508\,
            in2 => \_gnd_net_\,
            in3 => \N__24497\,
            lcout => \M_this_external_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_6\,
            carryout => \un1_M_this_external_address_q_cry_7\,
            clk => \N__25034\,
            ce => 'H',
            sr => \N__24745\
        );

    \M_this_external_address_q_8_LC_31_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25260\,
            in1 => \N__24478\,
            in2 => \_gnd_net_\,
            in3 => \N__24467\,
            lcout => \M_this_external_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_31_24_0_\,
            carryout => \un1_M_this_external_address_q_cry_8\,
            clk => \N__25035\,
            ce => 'H',
            sr => \N__24744\
        );

    \M_this_external_address_q_9_LC_31_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25276\,
            in1 => \N__24448\,
            in2 => \_gnd_net_\,
            in3 => \N__24437\,
            lcout => \M_this_external_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_8\,
            carryout => \un1_M_this_external_address_q_cry_9\,
            clk => \N__25035\,
            ce => 'H',
            sr => \N__24744\
        );

    \M_this_external_address_q_10_LC_31_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25257\,
            in1 => \N__24418\,
            in2 => \_gnd_net_\,
            in3 => \N__24407\,
            lcout => \M_this_external_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_9\,
            carryout => \un1_M_this_external_address_q_cry_10\,
            clk => \N__25035\,
            ce => 'H',
            sr => \N__24744\
        );

    \M_this_external_address_q_11_LC_31_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25274\,
            in1 => \N__24391\,
            in2 => \_gnd_net_\,
            in3 => \N__24380\,
            lcout => \M_this_external_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_10\,
            carryout => \un1_M_this_external_address_q_cry_11\,
            clk => \N__25035\,
            ce => 'H',
            sr => \N__24744\
        );

    \M_this_external_address_q_12_LC_31_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25258\,
            in1 => \N__24373\,
            in2 => \_gnd_net_\,
            in3 => \N__24362\,
            lcout => \M_this_external_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_11\,
            carryout => \un1_M_this_external_address_q_cry_12\,
            clk => \N__25035\,
            ce => 'H',
            sr => \N__24744\
        );

    \M_this_external_address_q_13_LC_31_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111101110"
        )
    port map (
            in0 => \N__25275\,
            in1 => \N__25315\,
            in2 => \_gnd_net_\,
            in3 => \N__25304\,
            lcout => \M_this_external_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_12\,
            carryout => \un1_M_this_external_address_q_cry_13\,
            clk => \N__25035\,
            ce => 'H',
            sr => \N__24744\
        );

    \M_this_external_address_q_14_LC_31_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25259\,
            in1 => \N__25291\,
            in2 => \_gnd_net_\,
            in3 => \N__25280\,
            lcout => \M_this_external_address_qZ0Z_14\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_13\,
            carryout => \un1_M_this_external_address_q_cry_14\,
            clk => \N__25035\,
            ce => 'H',
            sr => \N__24744\
        );

    \M_this_external_address_q_15_LC_31_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111101110"
        )
    port map (
            in0 => \N__25277\,
            in1 => \N__25048\,
            in2 => \_gnd_net_\,
            in3 => \N__25064\,
            lcout => \M_this_external_address_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25035\,
            ce => 'H',
            sr => \N__24744\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_o4_5_4_LC_32_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24644\,
            in1 => \N__24632\,
            in2 => \N__24620\,
            in3 => \N__24611\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_i_o4_5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
