-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     May 28 2022 12:21:16

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : inout std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    debug : out std_logic_vector(1 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    led : out std_logic_vector(7 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : inout std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__37833\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37279\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal port_data_rw_i_i : std_logic;
signal port_nmib_0_i : std_logic;
signal this_vga_signals_vvisibility_i : std_logic;
signal rgb_c_2 : std_logic;
signal rgb_c_1 : std_logic;
signal rgb_c_4 : std_logic;
signal \M_this_map_ram_write_data_4\ : std_logic;
signal \N_393_0\ : std_logic;
signal rgb_c_3 : std_logic;
signal \M_this_map_address_qZ0Z_0\ : std_logic;
signal \bfn_10_27_0_\ : std_logic;
signal \M_this_map_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_map_address_q_cry_0\ : std_logic;
signal \M_this_map_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_map_address_q_cry_1\ : std_logic;
signal \M_this_map_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_map_address_q_cry_2\ : std_logic;
signal \M_this_map_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_map_address_q_cry_3\ : std_logic;
signal \M_this_map_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_map_address_q_cry_4\ : std_logic;
signal \M_this_map_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_5\ : std_logic;
signal \M_this_map_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_map_address_q_cry_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_7\ : std_logic;
signal \M_this_map_address_qZ0Z_8\ : std_logic;
signal \bfn_10_28_0_\ : std_logic;
signal \un1_M_this_map_address_q_cry_8\ : std_logic;
signal \M_this_map_address_qZ0Z_9\ : std_logic;
signal rgb_c_0 : std_logic;
signal \this_vga_ramdac.i2_mux_cascade_\ : std_logic;
signal \this_vga_ramdac.N_3300_reto\ : std_logic;
signal \this_vga_ramdac.m6_cascade_\ : std_logic;
signal \this_vga_ramdac.N_3299_reto\ : std_logic;
signal rgb_c_5 : std_logic;
signal \this_vga_signals.N_729\ : std_logic;
signal \N_495\ : std_logic;
signal \this_vga_signals.un2_vsynclt8_cascade_\ : std_logic;
signal this_vga_signals_vsync_1_i : std_logic;
signal \this_vga_signals.vsync_1_2\ : std_logic;
signal \this_vga_signals.vsync_1_3\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_1_1_0_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_5_0_6\ : std_logic;
signal \this_vga_signals.N_5\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_0\ : std_logic;
signal \this_vga_signals.g2_5\ : std_logic;
signal \this_vga_signals.N_18_0\ : std_logic;
signal \this_vga_signals.g0_7_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0_0\ : std_logic;
signal \this_vga_signals.N_4_0_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_1\ : std_logic;
signal \this_vga_signals.if_N_5_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_1_1_0\ : std_logic;
signal \this_vga_ramdac.N_3301_reto\ : std_logic;
signal \this_vga_signals.vvisibility_1_cascade_\ : std_logic;
signal \this_vga_ramdac.m16\ : std_logic;
signal \this_vga_ramdac.m19_cascade_\ : std_logic;
signal \this_vga_ramdac.N_3302_reto\ : std_logic;
signal \this_vga_ramdac.N_3303_reto\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \this_vga_ramdac.i2_mux_0\ : std_logic;
signal \this_pixel_clk_M_counter_q_i_1\ : std_logic;
signal \this_pixel_clk_M_counter_q_0\ : std_logic;
signal \this_vga_ramdac.N_880_i_reto\ : std_logic;
signal \N_880_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal port_clk_c : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_0\ : std_logic;
signal \M_this_map_ram_write_data_1\ : std_logic;
signal \M_this_map_ram_write_data_5\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_0\ : std_logic;
signal \this_vga_signals.if_i1_mux_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \this_vga_signals.N_5_i_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3\ : std_logic;
signal \this_vga_signals.N_3_2_0_1\ : std_logic;
signal \this_vga_signals.g0_i_x4_0_0_cascade_\ : std_logic;
signal \this_vga_signals.N_3_3_0_0\ : std_logic;
signal \this_vga_signals.g0_0_2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_6_2\ : std_logic;
signal \this_vga_signals.g1_1_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.N_5_i_1_0_0\ : std_logic;
signal \this_vga_signals.g0_2_1_cascade_\ : std_logic;
signal \this_vga_signals.N_5_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_x1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_x0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_ns_cascade_\ : std_logic;
signal \this_vga_signals.g0_31_N_4L6\ : std_logic;
signal \this_vga_signals.g0_31_N_2L1_cascade_\ : std_logic;
signal \this_vga_signals.g0_31_N_5L8\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_0_cascade_\ : std_logic;
signal \this_vga_signals.N_2_0_cascade_\ : std_logic;
signal \this_vga_signals.M_this_vga_signals_pixel_clk_0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lt3_cascade_\ : std_logic;
signal \this_vga_ramdac.N_24_mux\ : std_logic;
signal \M_pcounter_q_ret_2_RNIH7PG8\ : std_logic;
signal \this_vga_ramdac.N_3298_reto\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_1_cascade_\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_0\ : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_axbxc3_1_cascade_\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \N_880_0\ : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0_2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1\ : std_logic;
signal \M_this_oam_ram_read_data_4\ : std_logic;
signal \M_this_map_ram_read_data_4\ : std_logic;
signal \M_this_ppu_sprites_addr_10\ : std_logic;
signal \M_this_map_ram_write_data_0\ : std_logic;
signal \M_this_map_ram_write_data_7\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.N_1_4_1_cascade_\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_2_3_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_8_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\ : std_logic;
signal \this_vga_signals.g0_0_0_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_3_0_0\ : std_logic;
signal \this_vga_signals.if_i2_mux\ : std_logic;
signal \this_vga_signals.g0_1_1_x0_cascade_\ : std_logic;
signal \this_vga_signals.g0_1_1_cascade_\ : std_logic;
signal \this_vga_signals.N_4_0_0_0\ : std_logic;
signal \this_vga_signals.g0_0_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.g1_5_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0_x1\ : std_logic;
signal \this_vga_signals.g1_2\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_ns\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c2_0\ : std_logic;
signal \this_vga_signals.N_3_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_3_1\ : std_logic;
signal \this_vga_signals.M_lcounter_d_0_sqmuxa_cascade_\ : std_logic;
signal \this_vga_signals.N_2_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_3_0\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lt7_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_d7_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0_1_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c2_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_9_1\ : std_logic;
signal \this_vga_signals.if_m7_0_x4_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0_2\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3\ : std_logic;
signal \this_vga_signals.SUM_3_i_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0_1_cascade_\ : std_logic;
signal \this_vga_signals.if_N_8_i_0\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lto7_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0\ : std_logic;
signal \M_hcounter_q_esr_RNIR18F4_9\ : std_logic;
signal \this_vga_signals.N_473_0_cascade_\ : std_logic;
signal \this_vga_signals.N_554\ : std_logic;
signal \this_vga_signals.SUM_3_i_1_0\ : std_logic;
signal \this_vga_signals.N_735_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_2_cascade_\ : std_logic;
signal \this_vga_signals.N_735_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_0_3\ : std_logic;
signal \this_vga_signals.hsync_1_i_0_1\ : std_logic;
signal \this_vga_signals.N_507_0\ : std_logic;
signal \M_this_map_ram_write_data_6\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_lcounter_d_0_sqmuxa\ : std_logic;
signal \this_vga_signals.M_hcounter_d7_0\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_7_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\ : std_logic;
signal \this_vga_signals.N_966_0\ : std_logic;
signal \this_vga_signals.N_1332_g\ : std_logic;
signal \this_vga_signals.g1_0_0_0_0\ : std_logic;
signal \this_vga_signals.g0_2_2_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i_2\ : std_logic;
signal \this_vga_signals.vaddress_3_6\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_2\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_2_cascade_\ : std_logic;
signal \this_vga_signals.g0_1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.vaddress_6_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_i\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_654_x0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_654_x1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_654_ns_cascade_\ : std_logic;
signal \this_vga_signals.if_m1_3\ : std_logic;
signal \this_vga_signals.if_m1_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x1\ : std_logic;
signal \this_vga_signals.vaddress_0_6\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_1_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3\ : std_logic;
signal \this_vga_signals.g1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3\ : std_logic;
signal \this_vga_signals.g0_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0_0_1\ : std_logic;
signal \this_vga_signals.N_3_1_0\ : std_logic;
signal \this_vga_signals.N_11_0_0_cascade_\ : std_logic;
signal \this_vga_signals.N_4_1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1\ : std_logic;
signal \this_vga_signals.if_m5_s\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lto8_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lto4_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_0\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.N_966_1\ : std_logic;
signal \this_sprites_ram.mem_WE_8\ : std_logic;
signal \M_this_map_ram_write_data_2\ : std_logic;
signal \this_vga_signals.vaddress_c2\ : std_logic;
signal \this_vga_signals.g0_0_0_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.g2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.g0_2_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_0\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_0_3\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_2_3\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_repZ0Z1\ : std_logic;
signal \this_vga_signals.vaddress_0_0_6_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_654_ns\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_x1\ : std_logic;
signal \this_vga_signals.g0_i_i_a5_1_0_0_0\ : std_logic;
signal \this_vga_signals.g0_i_i_0_0_0\ : std_logic;
signal \this_vga_signals.vaddress_2_6_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_0_0\ : std_logic;
signal \this_vga_signals.vaddress_6\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i_0_0\ : std_logic;
signal \this_vga_signals.N_7_1_0\ : std_logic;
signal \this_vga_signals.vaddress_5\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0\ : std_logic;
signal \this_vga_signals.vaddress_0_0_6\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1\ : std_logic;
signal \this_vga_signals.g0_0_0\ : std_logic;
signal \this_ppu.un13_0_cascade_\ : std_logic;
signal \this_ppu.M_line_clk_out_0_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lt9_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.un4_lvisibility_1\ : std_logic;
signal \this_vga_signals.line_clk_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.un4_lvisibility_1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_7\ : std_logic;
signal \M_this_vga_signals_line_clk_0_cascade_\ : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_0_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_1_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_2_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_3_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_4_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_5_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_6_s1\ : std_logic;
signal \this_ppu.M_count_q_RNO_0Z0Z_7\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_2\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_4\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.GZ0Z_394\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_501_0\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_1\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_2\ : std_logic;
signal \this_sprites_ram.mem_WE_10\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_7_cascade_\ : std_logic;
signal \N_597_cascade_\ : std_logic;
signal \M_this_sprites_address_qc_7_0\ : std_logic;
signal \N_1298_tz_0\ : std_logic;
signal \N_1294_tz_0\ : std_logic;
signal \N_602_cascade_\ : std_logic;
signal \M_this_sprites_address_qc_8_0\ : std_logic;
signal \M_this_map_ram_write_data_3\ : std_logic;
signal \M_this_oam_ram_read_data_2\ : std_logic;
signal \M_this_map_ram_read_data_2\ : std_logic;
signal \M_this_ppu_sprites_addr_8\ : std_logic;
signal \M_this_ppu_sprites_addr_5\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \M_this_ppu_sprites_addr_4\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \this_ppu.M_state_q_srsts_i_2_1_cascade_\ : std_logic;
signal \this_ppu.M_count_qZ0Z_6\ : std_logic;
signal \this_ppu.M_count_qZ0Z_7\ : std_logic;
signal \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_5_cascade_\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_5\ : std_logic;
signal \this_ppu.M_count_qZ0Z_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_8\ : std_logic;
signal \this_ppu.M_state_qZ0Z_1\ : std_logic;
signal \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_5\ : std_logic;
signal \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_4\ : std_logic;
signal \this_ppu.M_count_d_0_sqmuxa_1\ : std_logic;
signal \this_ppu.M_count_d_0_sqmuxa_1_cascade_\ : std_logic;
signal \this_ppu.M_line_clk_out_0\ : std_logic;
signal \this_ppu.N_1417_0\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\ : std_logic;
signal \this_ppu.N_1417_0_cascade_\ : std_logic;
signal \this_ppu.un13_0\ : std_logic;
signal \this_ppu.M_count_qZ0Z_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_2\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_3\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_6\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_7\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_4\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_5\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_0\ : std_logic;
signal \M_this_map_ram_read_data_5\ : std_logic;
signal \M_this_oam_ram_read_data_5\ : std_logic;
signal \M_this_map_ram_read_data_7\ : std_logic;
signal \M_this_oam_ram_read_data_7\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_2\ : std_logic;
signal \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0\ : std_logic;
signal \M_this_oam_ram_read_data_3\ : std_logic;
signal \M_this_map_ram_read_data_3\ : std_logic;
signal \M_this_ppu_sprites_addr_9\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_2\ : std_logic;
signal \M_this_substate_q_s_1\ : std_logic;
signal \M_this_sprites_address_q_0_0_i_480_cascade_\ : std_logic;
signal \M_this_sprites_address_qc_4_0\ : std_logic;
signal \N_511_1\ : std_logic;
signal \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_4\ : std_logic;
signal \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_5\ : std_logic;
signal \this_vga_signals.N_659_cascade_\ : std_logic;
signal \N_572_cascade_\ : std_logic;
signal \M_this_sprites_address_qc_2_0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_2\ : std_logic;
signal \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_3\ : std_logic;
signal \M_this_sprites_address_q_0_0_i_484\ : std_logic;
signal \M_this_sprites_address_qc_3_0_cascade_\ : std_logic;
signal \N_1318_tz_0\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_i_16\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0\ : std_logic;
signal \this_ppu.un2_vscroll_cry_0\ : std_logic;
signal \this_ppu.un2_vscroll_cry_1\ : std_logic;
signal \this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0\ : std_logic;
signal \M_this_oam_ram_read_data_i_17\ : std_logic;
signal \this_ppu.N_124\ : std_logic;
signal \this_ppu.N_124_cascade_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_2_c5_cascade_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_2_c5\ : std_logic;
signal \this_ppu.M_last_q\ : std_logic;
signal \this_ppu.M_state_qZ0Z_0\ : std_logic;
signal \M_this_vga_signals_line_clk_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_0\ : std_logic;
signal \this_ppu.vram_en_i_a2Z0Z_0\ : std_logic;
signal \this_ppu.vram_en_i_a2Z0Z_0_cascade_\ : std_logic;
signal \M_this_ppu_vram_en_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_haddress_q_3_c2_cascade_\ : std_logic;
signal \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2\ : std_logic;
signal \M_this_ppu_vram_data_2\ : std_logic;
signal \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0\ : std_logic;
signal \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\ : std_logic;
signal \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0_cascade_\ : std_logic;
signal \M_this_ppu_vram_data_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_2\ : std_logic;
signal \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\ : std_logic;
signal dma_0_i : std_logic;
signal \this_sprites_ram.mem_out_bus4_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_3\ : std_logic;
signal \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\ : std_logic;
signal \M_this_ppu_vram_data_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_3\ : std_logic;
signal \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_3\ : std_logic;
signal \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\ : std_logic;
signal \this_vga_signals.N_419_0_cascade_\ : std_logic;
signal \N_440_0_cascade_\ : std_logic;
signal \this_vga_signals.N_467_0_cascade_\ : std_logic;
signal \this_vga_signals.N_467_0\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0Z0Z_6\ : std_logic;
signal \N_510_0\ : std_logic;
signal \M_this_sprites_address_qc_5_0\ : std_logic;
signal \N_562_cascade_\ : std_logic;
signal \M_this_sprites_address_q_0_0_i_476\ : std_logic;
signal \M_this_sprites_address_q_0_0_i_496_cascade_\ : std_logic;
signal \M_this_sprites_address_qc_0_1\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_0\ : std_logic;
signal \N_773_cascade_\ : std_logic;
signal \M_this_sprites_address_q_0_0_i_492\ : std_logic;
signal \M_this_sprites_address_qc_1_0_cascade_\ : std_logic;
signal \N_896_0\ : std_logic;
signal \N_512_0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_8\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1Z0Z_5\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_11_cascade_\ : std_logic;
signal \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_1\ : std_logic;
signal \M_this_sprites_address_qc_10_0\ : std_logic;
signal \N_1286_tz_0_cascade_\ : std_logic;
signal \N_617\ : std_logic;
signal \M_this_sprites_address_qc_11_0\ : std_logic;
signal \bfn_19_5_0_\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_0\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_1\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_3\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_4\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_5\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_6\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_7\ : std_logic;
signal \bfn_19_6_0_\ : std_logic;
signal \this_ppu.M_this_ppu_vram_addr_i_0\ : std_logic;
signal \bfn_19_7_0_\ : std_logic;
signal \this_ppu.M_this_ppu_vram_addr_i_1\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_0\ : std_logic;
signal \this_ppu.M_this_ppu_vram_addr_i_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_1\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_0\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_2\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_1\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_3\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_4\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_3\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_5\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_4\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_6\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_7\ : std_logic;
signal \bfn_19_8_0_\ : std_logic;
signal \this_ppu.M_state_qZ0Z_2\ : std_logic;
signal \this_ppu.M_state_qZ0Z_3\ : std_logic;
signal \this_ppu.N_122\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_2_c2\ : std_logic;
signal this_vga_signals_vvisibility : std_logic;
signal \this_ppu.M_count_d_0_sqmuxa\ : std_logic;
signal \this_ppu.M_last_q_RNIQRTEB\ : std_logic;
signal \M_this_ppu_map_addr_1\ : std_logic;
signal \this_ppu.un1_M_haddress_q_3_c2\ : std_logic;
signal \M_this_ppu_map_addr_0\ : std_logic;
signal \M_this_ppu_map_addr_4\ : std_logic;
signal \this_ppu.un1_M_haddress_q_3_c5\ : std_logic;
signal \M_this_ppu_map_addr_2\ : std_logic;
signal \M_this_ppu_map_addr_3\ : std_logic;
signal \M_this_ppu_vram_en_0\ : std_logic;
signal \this_ppu.M_last_q_RNI3BB75\ : std_logic;
signal \M_this_oam_ram_read_data_1\ : std_logic;
signal \M_this_map_ram_read_data_1\ : std_logic;
signal \M_this_ppu_sprites_addr_7\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_1\ : std_logic;
signal \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_11\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\ : std_logic;
signal \M_this_ppu_vram_data_1\ : std_logic;
signal \M_this_oam_ram_read_data_6\ : std_logic;
signal \M_this_map_ram_read_data_6\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_12\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_1\ : std_logic;
signal \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_1\ : std_logic;
signal \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_1\ : std_logic;
signal \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_3\ : std_logic;
signal \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\ : std_logic;
signal \this_vga_signals.N_746_cascade_\ : std_logic;
signal \this_vga_signals.N_505\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_i_a4_2Z0Z_0\ : std_logic;
signal \this_vga_signals.N_459_0\ : std_logic;
signal \N_440_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_0\ : std_logic;
signal \un1_M_this_state_q_6_0\ : std_logic;
signal \M_this_sprites_address_q_RNIRO0N6Z0Z_0\ : std_logic;
signal \bfn_19_22_0_\ : std_logic;
signal \M_this_sprites_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_1\ : std_logic;
signal \M_this_sprites_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_2\ : std_logic;
signal \M_this_sprites_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_3\ : std_logic;
signal \M_this_sprites_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_4\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_5\ : std_logic;
signal \M_this_sprites_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_6\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_7\ : std_logic;
signal \M_this_sprites_address_qZ0Z_8\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0\ : std_logic;
signal \bfn_19_23_0_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_8\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_9\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_10\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_11\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_12\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_9\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_13\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\ : std_logic;
signal \N_627\ : std_logic;
signal \N_509_0_cascade_\ : std_logic;
signal \this_vga_signals.N_415_0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0\ : std_logic;
signal \M_this_sprites_address_q_0_0_i_472\ : std_logic;
signal \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_6\ : std_logic;
signal \N_773\ : std_logic;
signal \M_this_sprites_address_qZ0Z_6\ : std_logic;
signal \M_this_sprites_address_qc_6_0\ : std_logic;
signal \N_1282_tz_0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0\ : std_logic;
signal \N_1290_tz_0_cascade_\ : std_logic;
signal \N_607\ : std_logic;
signal \M_this_sprites_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_10_cascade_\ : std_logic;
signal \N_612\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_4\ : std_logic;
signal \bfn_20_6_0_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_0\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_1\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_2\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_3\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_4\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_5\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_6\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_7\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_7_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_7_THRU_CO\ : std_logic;
signal \bfn_20_7_0_\ : std_logic;
signal \this_ppu.vscroll8\ : std_logic;
signal \M_this_oam_ram_read_data_i_11\ : std_logic;
signal \this_ppu.un2_vscroll_axb_0\ : std_logic;
signal \M_this_ppu_sprites_addr_3\ : std_logic;
signal \M_this_state_q_RNI0A0EZ0Z_6\ : std_logic;
signal \M_this_state_q_RNI244K2Z0Z_6_cascade_\ : std_logic;
signal dma_0 : std_logic;
signal \M_this_state_q_fastZ0Z_9\ : std_logic;
signal \N_861\ : std_logic;
signal \N_861_cascade_\ : std_logic;
signal dma_c4_1 : std_logic;
signal this_vga_signals_un20_i_a2_4_a3_0_a4_2_1 : std_logic;
signal \N_460_0_cascade_\ : std_logic;
signal \N_560\ : std_logic;
signal \M_this_map_ram_write_en_0\ : std_logic;
signal \N_888_0_cascade_\ : std_logic;
signal \this_vga_signals.N_779\ : std_logic;
signal \this_start_data_delay_M_last_q\ : std_logic;
signal port_enb_c : std_logic;
signal \M_this_delay_clk_out_0\ : std_logic;
signal \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\ : std_logic;
signal port_address_in_2 : std_logic;
signal port_address_in_7 : std_logic;
signal port_rw_in : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_5LZ0Z8_cascade_\ : std_logic;
signal \M_this_substate_d_0_sqmuxa\ : std_logic;
signal \M_this_substate_d_0_sqmuxa_cascade_\ : std_logic;
signal dma_c4_1_0 : std_logic;
signal \this_vga_signals.N_732\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0\ : std_logic;
signal \N_622_cascade_\ : std_logic;
signal \N_1278_tz_0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_12\ : std_logic;
signal \M_this_sprites_address_qc_12_0\ : std_logic;
signal \this_vga_signals.N_427_0\ : std_logic;
signal \M_this_state_qZ0Z_1\ : std_logic;
signal \this_vga_signals.N_427_0_cascade_\ : std_logic;
signal \N_1274_tz_0\ : std_logic;
signal \M_this_sprites_address_qc_0_2\ : std_logic;
signal \this_vga_signals.N_889_0\ : std_logic;
signal \this_vga_signals.N_889_0_cascade_\ : std_logic;
signal \N_750\ : std_logic;
signal \N_762\ : std_logic;
signal \M_this_sprites_address_qZ0Z_9\ : std_logic;
signal \N_750_cascade_\ : std_logic;
signal \M_this_sprites_address_qc_9_0\ : std_logic;
signal port_address_in_0 : std_logic;
signal \this_vga_signals.N_648\ : std_logic;
signal port_address_in_1 : std_logic;
signal \N_460_0\ : std_logic;
signal \M_this_state_qZ0Z_8\ : std_logic;
signal \M_this_state_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0Z0Z_2\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_0_0_a2Z0Z_1\ : std_logic;
signal \M_this_state_qZ0Z_2\ : std_logic;
signal \N_250\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_3Z0Z_0_cascade_\ : std_logic;
signal \this_vga_signals.N_743\ : std_logic;
signal \N_228\ : std_logic;
signal \N_248\ : std_logic;
signal \M_this_oam_ram_read_data_16\ : std_logic;
signal \M_this_ppu_vram_addr_7\ : std_logic;
signal \this_ppu.M_this_ppu_vram_addr_i_7\ : std_logic;
signal \bfn_21_6_0_\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_1\ : std_logic;
signal \M_this_oam_ram_read_data_17\ : std_logic;
signal \this_ppu.M_vaddress_q_i_1\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_0\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_2\ : std_logic;
signal \M_this_oam_ram_read_data_18\ : std_logic;
signal \this_ppu.M_vaddress_q_i_2\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_1\ : std_logic;
signal \M_this_ppu_map_addr_5\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_5\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_2\ : std_logic;
signal \M_this_ppu_map_addr_6\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_6\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_3\ : std_logic;
signal \M_this_ppu_map_addr_7\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_7\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_4\ : std_logic;
signal \M_this_ppu_map_addr_8\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_8\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_5\ : std_logic;
signal \M_this_ppu_map_addr_9\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_9\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_6\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_7\ : std_logic;
signal \bfn_21_7_0_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO\ : std_logic;
signal \M_this_oam_ram_write_data_16\ : std_logic;
signal \M_this_oam_ram_read_data_i_19\ : std_logic;
signal \M_this_data_tmp_qZ0Z_16\ : std_logic;
signal this_vga_signals_un20_i_a2_0_a3_0_a4_2_2 : std_logic;
signal \this_sprites_ram.mem_out_bus5_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_0\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_13\ : std_logic;
signal \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\ : std_logic;
signal \M_this_state_qZ0Z_10\ : std_logic;
signal \this_vga_signals.N_433_0_cascade_\ : std_logic;
signal \this_vga_signals.N_442_0_cascade_\ : std_logic;
signal \this_vga_signals.N_719_cascade_\ : std_logic;
signal \this_vga_signals_M_this_data_count_q_3_0_a3_0_a4_0_2\ : std_logic;
signal \this_vga_signals_M_this_data_count_q_3_0_a3_0_a4_0_2_cascade_\ : std_logic;
signal \N_307_0_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_5\ : std_logic;
signal \this_vga_signals.N_665_1_cascade_\ : std_logic;
signal \M_this_data_count_q_3_0_13_cascade_\ : std_logic;
signal \N_755\ : std_logic;
signal \bfn_21_22_0_\ : std_logic;
signal \M_this_data_count_q_cry_0\ : std_logic;
signal \M_this_data_count_q_s_2\ : std_logic;
signal \M_this_data_count_q_cry_1\ : std_logic;
signal \M_this_data_count_q_cry_2\ : std_logic;
signal \M_this_data_count_q_cry_3\ : std_logic;
signal \M_this_data_count_q_cry_4\ : std_logic;
signal \M_this_data_count_q_cry_5\ : std_logic;
signal \M_this_data_count_q_cry_6\ : std_logic;
signal \M_this_data_count_q_cry_7\ : std_logic;
signal \M_this_data_count_q_s_8\ : std_logic;
signal \bfn_21_23_0_\ : std_logic;
signal \M_this_data_count_q_s_9\ : std_logic;
signal \M_this_data_count_q_cry_8\ : std_logic;
signal \M_this_data_count_q_cry_9_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_9\ : std_logic;
signal \M_this_data_count_q_s_11\ : std_logic;
signal \M_this_data_count_q_cry_10\ : std_logic;
signal \M_this_data_count_q_s_12\ : std_logic;
signal \M_this_data_count_q_cry_11\ : std_logic;
signal \M_this_data_count_q_cry_12_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_12\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \M_this_data_count_q_s_14\ : std_logic;
signal \M_this_data_count_q_cry_13\ : std_logic;
signal \M_this_data_count_q_cry_14\ : std_logic;
signal \M_this_data_count_q_s_15\ : std_logic;
signal \this_vga_signals.N_431_0\ : std_logic;
signal \this_vga_signals.N_428_0\ : std_logic;
signal \N_226\ : std_logic;
signal \M_this_data_tmp_qZ0Z_6\ : std_logic;
signal \M_this_oam_ram_write_data_6\ : std_logic;
signal \M_this_data_tmp_qZ0Z_2\ : std_logic;
signal \M_this_oam_ram_write_data_2\ : std_logic;
signal \M_this_data_tmp_qZ0Z_1\ : std_logic;
signal \M_this_oam_ram_write_data_1\ : std_logic;
signal \this_ppu.un1_oam_data_c2_cascade_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_6\ : std_logic;
signal \M_this_data_tmp_qZ0Z_23\ : std_logic;
signal \M_this_oam_ram_write_data_23\ : std_logic;
signal \M_this_oam_ram_read_data_22\ : std_logic;
signal \M_this_oam_ram_read_data_23\ : std_logic;
signal \this_ppu.un1_oam_data_c2\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_7\ : std_logic;
signal \M_this_oam_ram_write_data_25\ : std_logic;
signal \M_this_data_tmp_qZ0Z_17\ : std_logic;
signal \M_this_oam_ram_write_data_17\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_4\ : std_logic;
signal \M_this_oam_ram_write_data_24\ : std_logic;
signal \M_this_state_qZ0Z_12\ : std_logic;
signal \M_this_state_qZ0Z_11\ : std_logic;
signal \this_vga_signals.N_469_0_cascade_\ : std_logic;
signal \this_vga_signals.N_506_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_6\ : std_logic;
signal \M_this_data_count_qZ0Z_14\ : std_logic;
signal \M_this_data_count_qZ0Z_13\ : std_logic;
signal \M_this_data_count_qZ0Z_15\ : std_logic;
signal \M_this_data_count_qZ0Z_12\ : std_logic;
signal \this_vga_signals.N_745\ : std_logic;
signal \this_vga_signals.M_this_external_address_qlde_i_0_aZ0Z2\ : std_logic;
signal \this_vga_signals.N_442_0\ : std_logic;
signal \M_this_reset_cond_out_0\ : std_logic;
signal \this_vga_signals.M_this_external_address_qlde_i_0_aZ0Z2_cascade_\ : std_logic;
signal \this_vga_signals.M_this_data_count_qlde_iZ0Z_1\ : std_logic;
signal \M_this_data_count_qZ0Z_2\ : std_logic;
signal \M_this_data_count_qZ0Z_0\ : std_logic;
signal \M_this_state_d62_11\ : std_logic;
signal \M_this_state_d62_8_cascade_\ : std_logic;
signal \un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2\ : std_logic;
signal \M_this_state_d62_cascade_\ : std_logic;
signal \M_this_data_count_qZ0Z_10\ : std_logic;
signal \M_this_data_count_qZ0Z_9\ : std_logic;
signal \M_this_data_count_qZ0Z_11\ : std_logic;
signal \M_this_data_count_qZ0Z_8\ : std_logic;
signal \M_this_state_d62_10\ : std_logic;
signal \M_this_state_d62_9\ : std_logic;
signal \M_this_data_count_q_cry_0_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_1\ : std_logic;
signal \M_this_data_count_q_cry_2_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_3\ : std_logic;
signal \M_this_data_count_q_cry_3_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_4\ : std_logic;
signal \M_this_data_count_q_cry_4_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_5\ : std_logic;
signal \M_this_data_count_q_cry_5_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_6\ : std_logic;
signal \M_this_oam_ram_write_data_4\ : std_logic;
signal \M_this_data_tmp_qZ0Z_7\ : std_logic;
signal \M_this_oam_ram_write_data_7\ : std_logic;
signal \M_this_oam_ram_write_data_8\ : std_logic;
signal \M_this_oam_ram_write_data_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_4\ : std_logic;
signal \M_this_data_tmp_qZ0Z_0\ : std_logic;
signal \N_1412_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_3\ : std_logic;
signal \M_this_oam_ram_write_data_3\ : std_logic;
signal \M_this_oam_ram_write_data_10\ : std_logic;
signal \M_this_data_tmp_qZ0Z_10\ : std_logic;
signal \M_this_oam_ram_write_data_11\ : std_logic;
signal \M_this_oam_address_qZ0Z_5\ : std_logic;
signal \M_this_oam_address_qZ0Z_4\ : std_logic;
signal \M_this_data_tmp_qZ0Z_11\ : std_logic;
signal \M_this_data_tmp_qZ0Z_8\ : std_logic;
signal \N_413_0\ : std_logic;
signal \un1_M_this_oam_address_q_c4\ : std_logic;
signal \M_this_oam_address_qZ0Z_3\ : std_logic;
signal \M_this_oam_address_qZ0Z_2\ : std_logic;
signal \M_this_oam_address_qZ0Z_0\ : std_logic;
signal \M_this_state_qZ0Z_13\ : std_logic;
signal \M_this_oam_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_oam_address_q_c2\ : std_logic;
signal \this_vga_signals.N_461_0\ : std_logic;
signal \this_vga_signals.N_747\ : std_logic;
signal \M_this_state_qZ0Z_9\ : std_logic;
signal \M_this_state_qZ0Z_7\ : std_logic;
signal \this_vga_signals.N_433_0\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_i_1Z0Z_0\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_i_a4_4Z0Z_0\ : std_logic;
signal \M_this_state_d62\ : std_logic;
signal \this_vga_signals.N_746\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0Z0Z_12\ : std_logic;
signal \M_this_oam_address_q_0_i_o3_0_a2_5\ : std_logic;
signal \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0Z0Z_12_cascade_\ : std_logic;
signal led_c_1 : std_logic;
signal \M_this_substate_qZ0\ : std_logic;
signal \this_vga_signals.N_419_0\ : std_logic;
signal \M_this_data_count_q_cry_6_THRU_CO\ : std_logic;
signal \N_716_i\ : std_logic;
signal \M_this_data_count_qZ0Z_7\ : std_logic;
signal \N_364\ : std_logic;
signal port_data_c_0 : std_logic;
signal \M_this_state_qZ0Z_4\ : std_logic;
signal \N_888_0\ : std_logic;
signal \N_760_cascade_\ : std_logic;
signal \M_this_external_address_q_3_0_12\ : std_logic;
signal \this_sprites_ram.mem_WE_4\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_5\ : std_logic;
signal \M_this_oam_ram_write_data_13\ : std_logic;
signal \M_this_oam_ram_write_data_15\ : std_logic;
signal \M_this_oam_ram_read_data_15\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_7\ : std_logic;
signal \M_this_oam_ram_read_data_12\ : std_logic;
signal \M_this_oam_ram_read_data_11\ : std_logic;
signal \this_ppu.un1_oam_data_1_c2\ : std_logic;
signal \M_this_oam_ram_read_data_14\ : std_logic;
signal \this_ppu.un1_oam_data_1_c2_cascade_\ : std_logic;
signal \M_this_oam_ram_read_data_13\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_6\ : std_logic;
signal \M_this_data_tmp_qZ0Z_12\ : std_logic;
signal \M_this_oam_ram_write_data_12\ : std_logic;
signal \M_this_oam_ram_read_data_21\ : std_logic;
signal \M_this_oam_ram_read_data_20\ : std_logic;
signal \M_this_oam_ram_read_data_19\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_5\ : std_logic;
signal \M_this_data_tmp_qZ0Z_5\ : std_logic;
signal \M_this_oam_ram_write_data_5\ : std_logic;
signal \M_this_oam_ram_read_data_9\ : std_logic;
signal \M_this_oam_ram_write_data_9\ : std_logic;
signal \M_this_oam_ram_write_data_18\ : std_logic;
signal \M_this_oam_ram_write_data_20\ : std_logic;
signal \M_this_oam_ram_write_data_29\ : std_logic;
signal \M_this_oam_ram_write_data_30\ : std_logic;
signal \M_this_data_tmp_qZ0Z_22\ : std_logic;
signal \M_this_oam_ram_write_data_22\ : std_logic;
signal \M_this_oam_ram_write_data_31\ : std_logic;
signal \M_this_data_tmp_qZ0Z_18\ : std_logic;
signal \M_this_data_tmp_qZ0Z_20\ : std_logic;
signal port_data_c_4 : std_logic;
signal \M_this_oam_ram_write_data_28\ : std_logic;
signal \M_this_data_tmp_qZ0Z_21\ : std_logic;
signal \M_this_oam_ram_write_data_21\ : std_logic;
signal \M_this_oam_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_oam_address_q_c6\ : std_logic;
signal \M_this_oam_address_qZ0Z_7\ : std_logic;
signal \N_404_g\ : std_logic;
signal \M_this_data_tmp_qZ0Z_9\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_iZ0Z_8\ : std_logic;
signal \bfn_24_11_0_\ : std_logic;
signal \M_this_oam_ram_read_data_i_9\ : std_logic;
signal \this_ppu.un2_hscroll_cry_0\ : std_logic;
signal \M_this_oam_ram_read_data_10\ : std_logic;
signal \this_ppu.un2_hscroll_cry_1\ : std_logic;
signal \M_this_oam_ram_write_data_26\ : std_logic;
signal \M_this_oam_ram_write_data_19\ : std_logic;
signal \M_this_ppu_vram_addr_1\ : std_logic;
signal \this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0\ : std_logic;
signal \M_this_ppu_sprites_addr_1\ : std_logic;
signal \M_this_oam_ram_read_data_8\ : std_logic;
signal \M_this_ppu_vram_addr_2\ : std_logic;
signal \this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0\ : std_logic;
signal \M_this_ppu_sprites_addr_2\ : std_logic;
signal \this_ppu.un2_hscroll_axb_0\ : std_logic;
signal \M_this_ppu_vram_addr_0\ : std_logic;
signal \M_this_ppu_sprites_addr_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_19\ : std_logic;
signal \N_1396_0\ : std_logic;
signal \M_this_oam_ram_read_data_0\ : std_logic;
signal \M_this_map_ram_read_data_0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_4\ : std_logic;
signal \this_ppu.M_state_qZ0Z_5\ : std_logic;
signal \M_this_ppu_sprites_addr_6\ : std_logic;
signal \this_sprites_ram.mem_WE_14\ : std_logic;
signal \this_sprites_ram.mem_WE_12\ : std_logic;
signal \this_sprites_ram.mem_WE_0\ : std_logic;
signal port_data_c_1 : std_logic;
signal \this_vga_signals_M_this_external_address_q_3_i_0_0_15\ : std_logic;
signal \N_661\ : std_logic;
signal \this_sprites_ram.mem_WE_2\ : std_logic;
signal \this_vga_signals.N_665_1\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_3LZ0Z4\ : std_logic;
signal \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_4LZ0Z6\ : std_logic;
signal port_address_in_3 : std_logic;
signal port_address_in_5 : std_logic;
signal port_address_in_6 : std_logic;
signal port_address_in_4 : std_logic;
signal \this_vga_signals.un1_M_this_state_q_19_i_0_o2Z0Z_4\ : std_logic;
signal port_data_c_2 : std_logic;
signal \N_760\ : std_logic;
signal \M_this_sprites_address_qZ0Z_12\ : std_logic;
signal \N_25_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_13\ : std_logic;
signal \M_this_sprites_address_qZ0Z_11\ : std_logic;
signal \this_sprites_ram.mem_WE_6\ : std_logic;
signal \M_this_oam_ram_write_data_14\ : std_logic;
signal port_data_c_7 : std_logic;
signal \M_this_data_tmp_qZ0Z_15\ : std_logic;
signal port_data_c_6 : std_logic;
signal \M_this_data_tmp_qZ0Z_14\ : std_logic;
signal port_data_c_5 : std_logic;
signal \M_this_data_tmp_qZ0Z_13\ : std_logic;
signal \N_1404_0\ : std_logic;
signal \M_this_reset_cond_out_g_0\ : std_logic;
signal port_data_c_3 : std_logic;
signal \M_this_oam_ram_write_data_0_sqmuxa\ : std_logic;
signal \M_this_oam_ram_write_data_27\ : std_logic;
signal \M_this_external_address_q_3_0_13\ : std_logic;
signal \N_312_0\ : std_logic;
signal \M_this_external_address_qZ0Z_0\ : std_logic;
signal \bfn_26_21_0_\ : std_logic;
signal \M_this_external_address_qZ0Z_1\ : std_logic;
signal \M_this_external_address_q_cry_0\ : std_logic;
signal \M_this_external_address_qZ0Z_2\ : std_logic;
signal \M_this_external_address_q_cry_1\ : std_logic;
signal \M_this_external_address_qZ0Z_3\ : std_logic;
signal \M_this_external_address_q_cry_2\ : std_logic;
signal \M_this_external_address_qZ0Z_4\ : std_logic;
signal \M_this_external_address_q_cry_3\ : std_logic;
signal \M_this_external_address_qZ0Z_5\ : std_logic;
signal \M_this_external_address_q_cry_4\ : std_logic;
signal \M_this_external_address_qZ0Z_6\ : std_logic;
signal \M_this_external_address_q_cry_5\ : std_logic;
signal \N_49\ : std_logic;
signal \M_this_external_address_qZ0Z_7\ : std_logic;
signal \M_this_external_address_q_cry_6\ : std_logic;
signal \M_this_external_address_q_cry_7\ : std_logic;
signal clk_0_c_g : std_logic;
signal \N_47\ : std_logic;
signal \M_this_external_address_qZ0Z_8\ : std_logic;
signal \M_this_external_address_q_s_8\ : std_logic;
signal \bfn_26_22_0_\ : std_logic;
signal \M_this_external_address_qZ0Z_9\ : std_logic;
signal \M_this_external_address_q_s_9\ : std_logic;
signal \M_this_external_address_q_cry_8\ : std_logic;
signal \M_this_external_address_qZ0Z_10\ : std_logic;
signal \M_this_external_address_q_s_10\ : std_logic;
signal \M_this_external_address_q_cry_9\ : std_logic;
signal \M_this_external_address_qZ0Z_11\ : std_logic;
signal \M_this_external_address_q_s_11\ : std_logic;
signal \M_this_external_address_q_cry_10\ : std_logic;
signal \M_this_external_address_qZ0Z_12\ : std_logic;
signal \M_this_external_address_q_cry_11_THRU_CO\ : std_logic;
signal \M_this_external_address_q_cry_11\ : std_logic;
signal \M_this_external_address_qZ0Z_13\ : std_logic;
signal \M_this_external_address_q_cry_12_THRU_CO\ : std_logic;
signal \M_this_external_address_q_cry_12\ : std_logic;
signal \M_this_external_address_qZ0Z_14\ : std_logic;
signal \M_this_external_address_q_cry_13_THRU_CO\ : std_logic;
signal \M_this_external_address_q_cry_13\ : std_logic;
signal \M_this_external_address_qZ0Z_15\ : std_logic;
signal \M_this_external_address_q_cry_14\ : std_logic;
signal \M_this_external_address_q_s_15\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic_vector(1 downto 0);
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal led_wire : std_logic_vector(7 downto 0);
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_map_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    led <= led_wire;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \M_this_map_ram_read_data_3\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_2\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_1\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_0\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&\N__27978\&\N__27276\&\N__27342\&\N__27417\&\N__27486\&\N__21303\&\N__21174\&\N__21246\&\N__21447\&\N__21374\;
    \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&\N__11781\&\N__11814\&\N__11844\&\N__11874\&\N__11904\&\N__11934\&\N__11964\&\N__11610\&\N__11640\&\N__11667\;
    \this_map_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&\N__18555\&'0'&'0'&'0'&\N__15723\&'0'&'0'&'0'&\N__12507\&'0'&'0'&'0'&\N__13314\&'0';
    \M_this_map_ram_read_data_7\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_6\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_5\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_4\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&\N__27972\&\N__27269\&\N__27336\&\N__27411\&\N__27480\&\N__21297\&\N__21167\&\N__21236\&\N__21437\&\N__21362\;
    \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&\N__11775\&\N__11808\&\N__11838\&\N__11868\&\N__11898\&\N__11928\&\N__11958\&\N__11604\&\N__11634\&\N__11661\;
    \this_map_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&\N__13305\&'0'&'0'&'0'&\N__13968\&'0'&'0'&'0'&\N__12495\&'0'&'0'&'0'&\N__11709\&'0';
    \M_this_oam_ram_read_data_15\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(15);
    \M_this_oam_ram_read_data_14\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(14);
    \M_this_oam_ram_read_data_13\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_oam_ram_read_data_12\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(12);
    \M_this_oam_ram_read_data_11\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \M_this_oam_ram_read_data_10\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(10);
    \M_this_oam_ram_read_data_9\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_oam_ram_read_data_8\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(8);
    \M_this_oam_ram_read_data_7\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(7);
    \M_this_oam_ram_read_data_6\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(6);
    \M_this_oam_ram_read_data_5\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_oam_ram_read_data_4\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(4);
    \M_this_oam_ram_read_data_3\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_oam_ram_read_data_2\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_oam_ram_read_data_1\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_0\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__32241\&\N__32274\&\N__30120\&\N__30084\&\N__30747\&\N__30708\;
    \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ <= \N__31881\&\N__34590\&\N__31887\&\N__32148\&\N__30132\&\N__30150\&\N__31968\&\N__29859\&\N__29871\&\N__28395\&\N__32007\&\N__29898\&\N__30162\&\N__28371\&\N__28353\&\N__29850\;
    \M_this_oam_ram_read_data_23\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(7);
    \M_this_oam_ram_read_data_22\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(6);
    \M_this_oam_ram_read_data_21\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_oam_ram_read_data_20\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(4);
    \M_this_oam_ram_read_data_19\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \M_this_oam_ram_read_data_18\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(2);
    \M_this_oam_ram_read_data_17\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_16\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__32234\&\N__32268\&\N__30114\&\N__30078\&\N__30741\&\N__30702\;
    \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ <= \N__32466\&\N__31944\&\N__31950\&\N__32298\&\N__35511\&\N__33090\&\N__29172\&\N__29430\&\N__29253\&\N__32475\&\N__32280\&\N__31956\&\N__33078\&\N__31962\&\N__29154\&\N__27894\;
    \this_sprites_ram.mem_out_bus0_1\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_0\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ <= \N__13111\&\N__19232\&\N__18480\&\N__20987\&\N__33601\&\N__18279\&\N__18100\&\N__24773\&\N__32621\&\N__32878\&\N__34135\;
    \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ <= \N__24615\&\N__26076\&\N__23688\&\N__23937\&\N__24232\&\N__22110\&\N__22358\&\N__22608\&\N__22857\&\N__23087\&\N__23351\;
    \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26754\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28493\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus0_3\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_2\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ <= \N__13125\&\N__19233\&\N__18459\&\N__20997\&\N__33600\&\N__18194\&\N__18101\&\N__24802\&\N__32566\&\N__32842\&\N__34085\;
    \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ <= \N__24605\&\N__26072\&\N__23683\&\N__23961\&\N__24233\&\N__22106\&\N__22367\&\N__22604\&\N__22800\&\N__23110\&\N__23330\;
    \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26883\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__26653\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_1\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_0\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ <= \N__13107\&\N__19182\&\N__18460\&\N__20961\&\N__33550\&\N__18274\&\N__18024\&\N__24772\&\N__32534\&\N__32843\&\N__34062\;
    \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ <= \N__24589\&\N__26065\&\N__23682\&\N__23893\&\N__24205\&\N__22099\&\N__22368\&\N__22603\&\N__22858\&\N__23109\&\N__23329\;
    \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26753\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28485\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_3\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_2\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ <= \N__13105\&\N__19228\&\N__18491\&\N__20992\&\N__33524\&\N__18275\&\N__18099\&\N__24768\&\N__32567\&\N__32882\&\N__34111\;
    \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ <= \N__24588\&\N__26055\&\N__23667\&\N__23970\&\N__24206\&\N__22088\&\N__22345\&\N__22592\&\N__22859\&\N__23094\&\N__23328\;
    \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26879\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__26662\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_1\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_0\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ <= \N__13081\&\N__19146\&\N__18481\&\N__20993\&\N__33646\&\N__18316\&\N__18102\&\N__24809\&\N__32648\&\N__32971\&\N__34203\;
    \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ <= \N__24627\&\N__26019\&\N__23687\&\N__23963\&\N__24240\&\N__22046\&\N__22357\&\N__22557\&\N__22856\&\N__23111\&\N__23355\;
    \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26744\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28494\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_3\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_2\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ <= \N__13036\&\N__19230\&\N__18505\&\N__20995\&\N__33658\&\N__18328\&\N__18113\&\N__24810\&\N__32649\&\N__32983\&\N__34213\;
    \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ <= \N__24623\&\N__26018\&\N__23677\&\N__23942\&\N__24237\&\N__22041\&\N__22352\&\N__22556\&\N__22855\&\N__23011\&\N__23317\;
    \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26854\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__26664\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_1\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_0\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ <= \N__13082\&\N__19231\&\N__18506\&\N__20988\&\N__33665\&\N__18329\&\N__18114\&\N__24811\&\N__32650\&\N__32984\&\N__34214\;
    \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ <= \N__24616\&\N__25980\&\N__23654\&\N__23906\&\N__24238\&\N__22042\&\N__22356\&\N__22554\&\N__22853\&\N__23101\&\N__23353\;
    \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26745\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28489\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_3\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_2\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ <= \N__13112\&\N__19183\&\N__18510\&\N__20994\&\N__33666\&\N__18333\&\N__18112\&\N__24812\&\N__32651\&\N__32988\&\N__34215\;
    \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ <= \N__24593\&\N__26017\&\N__23681\&\N__23946\&\N__24236\&\N__22070\&\N__22366\&\N__22555\&\N__22854\&\N__23112\&\N__23354\;
    \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26855\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__26663\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_1\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_0\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ <= \N__13127\&\N__19214\&\N__18494\&\N__20957\&\N__33656\&\N__18326\&\N__18117\&\N__24808\&\N__32660\&\N__32981\&\N__34175\;
    \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ <= \N__24582\&\N__26042\&\N__23665\&\N__23968\&\N__24222\&\N__22084\&\N__22279\&\N__22587\&\N__22863\&\N__23089\&\N__23335\;
    \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26748\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28460\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_3\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_2\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ <= \N__13131\&\N__19193\&\N__18495\&\N__20956\&\N__33657\&\N__18327\&\N__18116\&\N__24813\&\N__32661\&\N__32982\&\N__34190\;
    \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ <= \N__24583\&\N__26041\&\N__23653\&\N__23969\&\N__24223\&\N__22098\&\N__22348\&\N__22602\&\N__22817\&\N__23108\&\N__23336\;
    \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26877\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__26660\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_1\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_0\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ <= \N__13106\&\N__19213\&\N__18493\&\N__20916\&\N__33639\&\N__18312\&\N__18106\&\N__24804\&\N__32653\&\N__32964\&\N__34174\;
    \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ <= \N__24581\&\N__26020\&\N__23664\&\N__23954\&\N__24224\&\N__22083\&\N__22365\&\N__22586\&\N__22869\&\N__23088\&\N__23334\;
    \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26749\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28445\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_3\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_2\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ <= \N__13118\&\N__19181\&\N__18492\&\N__20980\&\N__33638\&\N__18308\&\N__18110\&\N__24780\&\N__32652\&\N__32963\&\N__34157\;
    \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ <= \N__24580\&\N__26024\&\N__23629\&\N__23883\&\N__24225\&\N__22060\&\N__22335\&\N__22559\&\N__22864\&\N__23055\&\N__23352\;
    \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26856\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__26651\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_1\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_0\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ <= \N__13117\&\N__19215\&\N__18467\&\N__20976\&\N__33613\&\N__18288\&\N__18111\&\N__24803\&\N__32635\&\N__32938\&\N__34156\;
    \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ <= \N__24584\&\N__25990\&\N__23628\&\N__23947\&\N__24149\&\N__22059\&\N__22334\&\N__22558\&\N__22801\&\N__23054\&\N__23337\;
    \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26747\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28444\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_3\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_2\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ <= \N__13086\&\N__19212\&\N__18466\&\N__20996\&\N__33612\&\N__18281\&\N__18115\&\N__24776\&\N__32634\&\N__32937\&\N__34137\;
    \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ <= \N__24585\&\N__26028\&\N__23636\&\N__23938\&\N__24239\&\N__22014\&\N__22347\&\N__22569\&\N__22845\&\N__22974\&\N__23307\;
    \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26853\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__26652\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_1\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_0\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ <= \N__13113\&\N__19165\&\N__18465\&\N__20972\&\N__33582\&\N__18280\&\N__18094\&\N__24775\&\N__32603\&\N__32909\&\N__34136\;
    \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ <= \N__24586\&\N__26029\&\N__23637\&\N__23964\&\N__24235\&\N__22047\&\N__22346\&\N__22570\&\N__22852\&\N__23065\&\N__23341\;
    \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26746\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28461\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_3\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_2\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ <= \N__13126\&\N__19229\&\N__18464\&\N__20962\&\N__33581\&\N__18307\&\N__18098\&\N__24774\&\N__32602\&\N__32908\&\N__34112\;
    \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ <= \N__24587\&\N__26043\&\N__23666\&\N__23962\&\N__24234\&\N__22071\&\N__22309\&\N__22591\&\N__22868\&\N__23093\&\N__23327\;
    \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__26878\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__26661\&'0'&'0'&'0';
    \M_this_vram_read_data_3\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_vram_read_data_2\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_vram_read_data_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_vram_read_data_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__12696\&\N__11700\&\N__12570\&\N__12540\&\N__12555\&\N__13236\&\N__12807\&\N__12786\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__27824\&\N__21170\&\N__21245\&\N__21446\&\N__21375\&\N__32754\&\N__33065\&\N__34314\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20013\&\N__19803\&\N__21720\&\N__19758\;

    \this_map_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36969\,
            RE => \N__28934\,
            WCLKE => \N__25299\,
            WCLK => \N__36970\,
            WE => \N__28851\
        );

    \this_map_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36973\,
            RE => \N__28935\,
            WCLKE => \N__25292\,
            WCLK => \N__36974\,
            WE => \N__28852\
        );

    \this_oam_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36859\,
            RE => \N__29117\,
            WCLKE => \N__35709\,
            WCLK => \N__36860\,
            WE => \N__29102\
        );

    \this_oam_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36874\,
            RE => \N__29081\,
            WCLKE => \N__35708\,
            WCLK => \N__36875\,
            WE => \N__29098\
        );

    \this_sprites_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36891\,
            RE => \N__29068\,
            WCLKE => \N__33483\,
            WCLK => \N__36890\,
            WE => \N__29025\
        );

    \this_sprites_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36901\,
            RE => \N__29023\,
            WCLKE => \N__33482\,
            WCLK => \N__36902\,
            WE => \N__29024\
        );

    \this_sprites_ram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36917\,
            RE => \N__29011\,
            WCLKE => \N__33458\,
            WCLK => \N__36918\,
            WE => \N__28939\
        );

    \this_sprites_ram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36929\,
            RE => \N__28937\,
            WCLKE => \N__33459\,
            WCLK => \N__36930\,
            WE => \N__28938\
        );

    \this_sprites_ram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36945\,
            RE => \N__28717\,
            WCLKE => \N__17450\,
            WCLK => \N__36946\,
            WE => \N__28778\
        );

    \this_sprites_ram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36952\,
            RE => \N__28736\,
            WCLKE => \N__17451\,
            WCLK => \N__36953\,
            WE => \N__28779\
        );

    \this_sprites_ram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36959\,
            RE => \N__28737\,
            WCLKE => \N__15753\,
            WCLK => \N__36960\,
            WE => \N__28842\
        );

    \this_sprites_ram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36964\,
            RE => \N__28850\,
            WCLKE => \N__15752\,
            WCLK => \N__36965\,
            WE => \N__28843\
        );

    \this_sprites_ram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36975\,
            RE => \N__29121\,
            WCLKE => \N__34607\,
            WCLK => \N__36976\,
            WE => \N__29122\
        );

    \this_sprites_ram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36977\,
            RE => \N__28936\,
            WCLKE => \N__34608\,
            WCLK => \N__36978\,
            WE => \N__29123\
        );

    \this_sprites_ram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36971\,
            RE => \N__28853\,
            WCLKE => \N__31929\,
            WCLK => \N__36972\,
            WE => \N__29107\
        );

    \this_sprites_ram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36967\,
            RE => \N__29061\,
            WCLKE => \N__31925\,
            WCLK => \N__36968\,
            WE => \N__29106\
        );

    \this_sprites_ram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36961\,
            RE => \N__29082\,
            WCLKE => \N__33174\,
            WCLK => \N__36962\,
            WE => \N__29083\
        );

    \this_sprites_ram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36955\,
            RE => \N__29066\,
            WCLKE => \N__33170\,
            WCLK => \N__36956\,
            WE => \N__29067\
        );

    \this_sprites_ram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36949\,
            RE => \N__29042\,
            WCLKE => \N__33432\,
            WCLK => \N__36950\,
            WE => \N__29016\
        );

    \this_sprites_ram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36939\,
            RE => \N__29065\,
            WCLKE => \N__33428\,
            WCLK => \N__36940\,
            WE => \N__29015\
        );

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__36934\,
            RE => \N__28652\,
            WCLKE => \N__21102\,
            WCLK => \N__36935\,
            WE => \N__28660\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__37831\,
            GLOBALBUFFEROUTPUT => clk_0_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37833\,
            DIN => \N__37832\,
            DOUT => \N__37831\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37833\,
            PADOUT => \N__37832\,
            PADIN => \N__37831\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37822\,
            DIN => \N__37821\,
            DOUT => \N__37820\,
            PACKAGEPIN => debug_wire(0)
        );

    \debug_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37822\,
            PADOUT => \N__37821\,
            PADIN => \N__37820\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37813\,
            DIN => \N__37812\,
            DOUT => \N__37811\,
            PACKAGEPIN => debug_wire(1)
        );

    \debug_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37813\,
            PADOUT => \N__37812\,
            PADIN => \N__37811\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37804\,
            DIN => \N__37803\,
            DOUT => \N__37802\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37804\,
            PADOUT => \N__37803\,
            PADIN => \N__37802\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12114\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37795\,
            DIN => \N__37794\,
            DOUT => \N__37793\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37795\,
            PADOUT => \N__37794\,
            PADIN => \N__37793\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13743\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37786\,
            DIN => \N__37785\,
            DOUT => \N__37784\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37786\,
            PADOUT => \N__37785\,
            PADIN => \N__37784\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__29124\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37777\,
            DIN => \N__37776\,
            DOUT => \N__37775\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37777\,
            PADOUT => \N__37776\,
            PADIN => \N__37775\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__31653\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37768\,
            DIN => \N__37767\,
            DOUT => \N__37766\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37768\,
            PADOUT => \N__37767\,
            PADIN => \N__37766\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37759\,
            DIN => \N__37758\,
            DOUT => \N__37757\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37759\,
            PADOUT => \N__37758\,
            PADIN => \N__37757\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37750\,
            DIN => \N__37749\,
            DOUT => \N__37748\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37750\,
            PADOUT => \N__37749\,
            PADIN => \N__37748\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37741\,
            DIN => \N__37740\,
            DOUT => \N__37739\,
            PACKAGEPIN => led_wire(5)
        );

    \led_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37741\,
            PADOUT => \N__37740\,
            PADIN => \N__37739\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37732\,
            DIN => \N__37731\,
            DOUT => \N__37730\,
            PACKAGEPIN => led_wire(6)
        );

    \led_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37732\,
            PADOUT => \N__37731\,
            PADIN => \N__37730\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37723\,
            DIN => \N__37722\,
            DOUT => \N__37721\,
            PACKAGEPIN => led_wire(7)
        );

    \led_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37723\,
            PADOUT => \N__37722\,
            PADIN => \N__37721\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37714\,
            DIN => \N__37713\,
            DOUT => \N__37712\,
            PACKAGEPIN => port_address(0)
        );

    \port_address_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37714\,
            PADOUT => \N__37713\,
            PADIN => \N__37712\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__35484\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20157\
        );

    \port_address_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37705\,
            DIN => \N__37704\,
            DOUT => \N__37703\,
            PACKAGEPIN => port_address(1)
        );

    \port_address_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37705\,
            PADOUT => \N__37704\,
            PADIN => \N__37703\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__35457\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20211\
        );

    \port_address_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37696\,
            DIN => \N__37695\,
            DOUT => \N__37694\,
            PACKAGEPIN => port_address(2)
        );

    \port_address_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37696\,
            PADOUT => \N__37695\,
            PADIN => \N__37694\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__35436\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20187\
        );

    \port_address_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37687\,
            DIN => \N__37686\,
            DOUT => \N__37685\,
            PACKAGEPIN => port_address(3)
        );

    \port_address_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37687\,
            PADOUT => \N__37686\,
            PADIN => \N__37685\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__35409\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20155\
        );

    \port_address_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37678\,
            DIN => \N__37677\,
            DOUT => \N__37676\,
            PACKAGEPIN => port_address(4)
        );

    \port_address_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37678\,
            PADOUT => \N__37677\,
            PADIN => \N__37676\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__35382\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20214\
        );

    \port_address_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37669\,
            DIN => \N__37668\,
            DOUT => \N__37667\,
            PACKAGEPIN => port_address(5)
        );

    \port_address_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37669\,
            PADOUT => \N__37668\,
            PADIN => \N__37667\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__37158\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20212\
        );

    \port_address_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37660\,
            DIN => \N__37659\,
            DOUT => \N__37658\,
            PACKAGEPIN => port_address(6)
        );

    \port_address_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37660\,
            PADOUT => \N__37659\,
            PADIN => \N__37658\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__37140\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20192\
        );

    \port_address_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37651\,
            DIN => \N__37650\,
            DOUT => \N__37649\,
            PACKAGEPIN => port_address(7)
        );

    \port_address_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37651\,
            PADOUT => \N__37650\,
            PADIN => \N__37649\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__37008\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20229\
        );

    \port_address_obuft_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37642\,
            DIN => \N__37641\,
            DOUT => \N__37640\,
            PACKAGEPIN => port_address(10)
        );

    \port_address_obuft_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37642\,
            PADOUT => \N__37641\,
            PADIN => \N__37640\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__36438\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20159\
        );

    \port_address_obuft_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37633\,
            DIN => \N__37632\,
            DOUT => \N__37631\,
            PACKAGEPIN => port_address(11)
        );

    \port_address_obuft_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37633\,
            PADOUT => \N__37632\,
            PADIN => \N__37631\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__36399\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20156\
        );

    \port_address_obuft_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37624\,
            DIN => \N__37623\,
            DOUT => \N__37622\,
            PACKAGEPIN => port_address(12)
        );

    \port_address_obuft_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37624\,
            PADOUT => \N__37623\,
            PADIN => \N__37622\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37353\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20215\
        );

    \port_address_obuft_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37615\,
            DIN => \N__37614\,
            DOUT => \N__37613\,
            PACKAGEPIN => port_address(13)
        );

    \port_address_obuft_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37615\,
            PADOUT => \N__37614\,
            PADIN => \N__37613\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37305\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20213\
        );

    \port_address_obuft_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37606\,
            DIN => \N__37605\,
            DOUT => \N__37604\,
            PACKAGEPIN => port_address(14)
        );

    \port_address_obuft_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37606\,
            PADOUT => \N__37605\,
            PADIN => \N__37604\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37260\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20151\
        );

    \port_address_obuft_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37597\,
            DIN => \N__37596\,
            DOUT => \N__37595\,
            PACKAGEPIN => port_address(15)
        );

    \port_address_obuft_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37597\,
            PADOUT => \N__37596\,
            PADIN => \N__37595\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37215\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20228\
        );

    \port_address_obuft_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37588\,
            DIN => \N__37587\,
            DOUT => \N__37586\,
            PACKAGEPIN => port_address(8)
        );

    \port_address_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37588\,
            PADOUT => \N__37587\,
            PADIN => \N__37586\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__36525\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20158\
        );

    \port_address_obuft_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37579\,
            DIN => \N__37578\,
            DOUT => \N__37577\,
            PACKAGEPIN => port_address(9)
        );

    \port_address_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37579\,
            PADOUT => \N__37578\,
            PADIN => \N__37577\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__36483\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20188\
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37570\,
            DIN => \N__37569\,
            DOUT => \N__37568\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37570\,
            PADOUT => \N__37569\,
            PADIN => \N__37568\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37561\,
            DIN => \N__37560\,
            DOUT => \N__37559\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37561\,
            PADOUT => \N__37560\,
            PADIN => \N__37559\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37552\,
            DIN => \N__37551\,
            DOUT => \N__37550\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37552\,
            PADOUT => \N__37551\,
            PADIN => \N__37550\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37543\,
            DIN => \N__37542\,
            DOUT => \N__37541\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37543\,
            PADOUT => \N__37542\,
            PADIN => \N__37541\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37534\,
            DIN => \N__37533\,
            DOUT => \N__37532\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37534\,
            PADOUT => \N__37533\,
            PADIN => \N__37532\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37525\,
            DIN => \N__37524\,
            DOUT => \N__37523\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37525\,
            PADOUT => \N__37524\,
            PADIN => \N__37523\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37516\,
            DIN => \N__37515\,
            DOUT => \N__37514\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37516\,
            PADOUT => \N__37515\,
            PADIN => \N__37514\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37507\,
            DIN => \N__37506\,
            DOUT => \N__37505\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37507\,
            PADOUT => \N__37506\,
            PADIN => \N__37505\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37498\,
            DIN => \N__37497\,
            DOUT => \N__37496\,
            PACKAGEPIN => port_data_wire(7)
        );

    \port_data_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37498\,
            PADOUT => \N__37497\,
            PADIN => \N__37496\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37489\,
            DIN => \N__37488\,
            DOUT => \N__37487\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37489\,
            PADOUT => \N__37488\,
            PADIN => \N__37487\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11583\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37480\,
            DIN => \N__37479\,
            DOUT => \N__37478\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37480\,
            PADOUT => \N__37479\,
            PADIN => \N__37478\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__24984\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37471\,
            DIN => \N__37470\,
            DOUT => \N__37469\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37471\,
            PADOUT => \N__37470\,
            PADIN => \N__37469\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37462\,
            DIN => \N__37461\,
            DOUT => \N__37460\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37462\,
            PADOUT => \N__37461\,
            PADIN => \N__37460\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11577\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37453\,
            DIN => \N__37452\,
            DOUT => \N__37451\,
            PACKAGEPIN => port_rw
        );

    \port_rw_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__37453\,
            PADOUT => \N__37452\,
            PADIN => \N__37451\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_in,
            DIN1 => OPEN,
            DOUT0 => \N__28777\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__20221\
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37444\,
            DIN => \N__37443\,
            DOUT => \N__37442\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37444\,
            PADOUT => \N__37443\,
            PADIN => \N__37442\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12051\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37435\,
            DIN => \N__37434\,
            DOUT => \N__37433\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37435\,
            PADOUT => \N__37434\,
            PADIN => \N__37433\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11742\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37426\,
            DIN => \N__37425\,
            DOUT => \N__37424\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37426\,
            PADOUT => \N__37425\,
            PADIN => \N__37424\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11754\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37417\,
            DIN => \N__37416\,
            DOUT => \N__37415\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37417\,
            PADOUT => \N__37416\,
            PADIN => \N__37415\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11688\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37408\,
            DIN => \N__37407\,
            DOUT => \N__37406\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37408\,
            PADOUT => \N__37407\,
            PADIN => \N__37406\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11733\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37399\,
            DIN => \N__37398\,
            DOUT => \N__37397\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37399\,
            PADOUT => \N__37398\,
            PADIN => \N__37397\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12000\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37390\,
            DIN => \N__37389\,
            DOUT => \N__37388\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37390\,
            PADOUT => \N__37389\,
            PADIN => \N__37388\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37381\,
            DIN => \N__37380\,
            DOUT => \N__37379\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37381\,
            PADOUT => \N__37380\,
            PADIN => \N__37379\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11568\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37372\,
            DIN => \N__37371\,
            DOUT => \N__37370\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37372\,
            PADOUT => \N__37371\,
            PADIN => \N__37370\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12090\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__9454\ : IoInMux
    port map (
            O => \N__37353\,
            I => \N__37350\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__37350\,
            I => \N__37347\
        );

    \I__9452\ : Span4Mux_s1_h
    port map (
            O => \N__37347\,
            I => \N__37344\
        );

    \I__9451\ : Span4Mux_h
    port map (
            O => \N__37344\,
            I => \N__37339\
        );

    \I__9450\ : CascadeMux
    port map (
            O => \N__37343\,
            I => \N__37336\
        );

    \I__9449\ : InMux
    port map (
            O => \N__37342\,
            I => \N__37333\
        );

    \I__9448\ : Span4Mux_h
    port map (
            O => \N__37339\,
            I => \N__37330\
        );

    \I__9447\ : InMux
    port map (
            O => \N__37336\,
            I => \N__37327\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__37333\,
            I => \N__37324\
        );

    \I__9445\ : Odrv4
    port map (
            O => \N__37330\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__37327\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__9443\ : Odrv12
    port map (
            O => \N__37324\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__9442\ : InMux
    port map (
            O => \N__37317\,
            I => \N__37314\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__37314\,
            I => \N__37311\
        );

    \I__9440\ : Odrv4
    port map (
            O => \N__37311\,
            I => \M_this_external_address_q_cry_11_THRU_CO\
        );

    \I__9439\ : InMux
    port map (
            O => \N__37308\,
            I => \M_this_external_address_q_cry_11\
        );

    \I__9438\ : IoInMux
    port map (
            O => \N__37305\,
            I => \N__37302\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__37302\,
            I => \N__37299\
        );

    \I__9436\ : IoSpan4Mux
    port map (
            O => \N__37299\,
            I => \N__37294\
        );

    \I__9435\ : CascadeMux
    port map (
            O => \N__37298\,
            I => \N__37291\
        );

    \I__9434\ : InMux
    port map (
            O => \N__37297\,
            I => \N__37288\
        );

    \I__9433\ : Sp12to4
    port map (
            O => \N__37294\,
            I => \N__37285\
        );

    \I__9432\ : InMux
    port map (
            O => \N__37291\,
            I => \N__37282\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__37288\,
            I => \N__37279\
        );

    \I__9430\ : Odrv12
    port map (
            O => \N__37285\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__37282\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__9428\ : Odrv12
    port map (
            O => \N__37279\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__9427\ : InMux
    port map (
            O => \N__37272\,
            I => \N__37269\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__37269\,
            I => \N__37266\
        );

    \I__9425\ : Odrv4
    port map (
            O => \N__37266\,
            I => \M_this_external_address_q_cry_12_THRU_CO\
        );

    \I__9424\ : InMux
    port map (
            O => \N__37263\,
            I => \M_this_external_address_q_cry_12\
        );

    \I__9423\ : IoInMux
    port map (
            O => \N__37260\,
            I => \N__37257\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__37257\,
            I => \N__37254\
        );

    \I__9421\ : Span4Mux_s3_h
    port map (
            O => \N__37254\,
            I => \N__37249\
        );

    \I__9420\ : CascadeMux
    port map (
            O => \N__37253\,
            I => \N__37246\
        );

    \I__9419\ : InMux
    port map (
            O => \N__37252\,
            I => \N__37243\
        );

    \I__9418\ : Span4Mux_v
    port map (
            O => \N__37249\,
            I => \N__37240\
        );

    \I__9417\ : InMux
    port map (
            O => \N__37246\,
            I => \N__37237\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__37243\,
            I => \N__37234\
        );

    \I__9415\ : Odrv4
    port map (
            O => \N__37240\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__37237\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__9413\ : Odrv4
    port map (
            O => \N__37234\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__9412\ : InMux
    port map (
            O => \N__37227\,
            I => \N__37224\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__37224\,
            I => \N__37221\
        );

    \I__9410\ : Odrv4
    port map (
            O => \N__37221\,
            I => \M_this_external_address_q_cry_13_THRU_CO\
        );

    \I__9409\ : InMux
    port map (
            O => \N__37218\,
            I => \M_this_external_address_q_cry_13\
        );

    \I__9408\ : IoInMux
    port map (
            O => \N__37215\,
            I => \N__37212\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__37212\,
            I => \N__37209\
        );

    \I__9406\ : IoSpan4Mux
    port map (
            O => \N__37209\,
            I => \N__37206\
        );

    \I__9405\ : Span4Mux_s3_h
    port map (
            O => \N__37206\,
            I => \N__37203\
        );

    \I__9404\ : Span4Mux_v
    port map (
            O => \N__37203\,
            I => \N__37199\
        );

    \I__9403\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37196\
        );

    \I__9402\ : Span4Mux_v
    port map (
            O => \N__37199\,
            I => \N__37193\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__37196\,
            I => \N__37190\
        );

    \I__9400\ : Span4Mux_h
    port map (
            O => \N__37193\,
            I => \N__37187\
        );

    \I__9399\ : Span4Mux_h
    port map (
            O => \N__37190\,
            I => \N__37184\
        );

    \I__9398\ : Odrv4
    port map (
            O => \N__37187\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__9397\ : Odrv4
    port map (
            O => \N__37184\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__9396\ : InMux
    port map (
            O => \N__37179\,
            I => \M_this_external_address_q_cry_14\
        );

    \I__9395\ : CascadeMux
    port map (
            O => \N__37176\,
            I => \N__37173\
        );

    \I__9394\ : InMux
    port map (
            O => \N__37173\,
            I => \N__37170\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__37170\,
            I => \N__37167\
        );

    \I__9392\ : Span4Mux_h
    port map (
            O => \N__37167\,
            I => \N__37164\
        );

    \I__9391\ : Odrv4
    port map (
            O => \N__37164\,
            I => \M_this_external_address_q_s_15\
        );

    \I__9390\ : InMux
    port map (
            O => \N__37161\,
            I => \M_this_external_address_q_cry_3\
        );

    \I__9389\ : IoInMux
    port map (
            O => \N__37158\,
            I => \N__37155\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__37155\,
            I => \N__37151\
        );

    \I__9387\ : InMux
    port map (
            O => \N__37154\,
            I => \N__37148\
        );

    \I__9386\ : Odrv12
    port map (
            O => \N__37151\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__37148\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__9384\ : InMux
    port map (
            O => \N__37143\,
            I => \M_this_external_address_q_cry_4\
        );

    \I__9383\ : IoInMux
    port map (
            O => \N__37140\,
            I => \N__37137\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__37137\,
            I => \N__37134\
        );

    \I__9381\ : Span4Mux_s3_h
    port map (
            O => \N__37134\,
            I => \N__37131\
        );

    \I__9380\ : Span4Mux_v
    port map (
            O => \N__37131\,
            I => \N__37127\
        );

    \I__9379\ : InMux
    port map (
            O => \N__37130\,
            I => \N__37124\
        );

    \I__9378\ : Odrv4
    port map (
            O => \N__37127\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__37124\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__9376\ : InMux
    port map (
            O => \N__37119\,
            I => \M_this_external_address_q_cry_5\
        );

    \I__9375\ : InMux
    port map (
            O => \N__37116\,
            I => \N__37100\
        );

    \I__9374\ : InMux
    port map (
            O => \N__37115\,
            I => \N__37100\
        );

    \I__9373\ : InMux
    port map (
            O => \N__37114\,
            I => \N__37097\
        );

    \I__9372\ : InMux
    port map (
            O => \N__37113\,
            I => \N__37092\
        );

    \I__9371\ : InMux
    port map (
            O => \N__37112\,
            I => \N__37092\
        );

    \I__9370\ : InMux
    port map (
            O => \N__37111\,
            I => \N__37083\
        );

    \I__9369\ : InMux
    port map (
            O => \N__37110\,
            I => \N__37083\
        );

    \I__9368\ : InMux
    port map (
            O => \N__37109\,
            I => \N__37083\
        );

    \I__9367\ : InMux
    port map (
            O => \N__37108\,
            I => \N__37083\
        );

    \I__9366\ : InMux
    port map (
            O => \N__37107\,
            I => \N__37072\
        );

    \I__9365\ : InMux
    port map (
            O => \N__37106\,
            I => \N__37072\
        );

    \I__9364\ : InMux
    port map (
            O => \N__37105\,
            I => \N__37072\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__37100\,
            I => \N__37069\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__37097\,
            I => \N__37066\
        );

    \I__9361\ : LocalMux
    port map (
            O => \N__37092\,
            I => \N__37063\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__37083\,
            I => \N__37060\
        );

    \I__9359\ : InMux
    port map (
            O => \N__37082\,
            I => \N__37051\
        );

    \I__9358\ : InMux
    port map (
            O => \N__37081\,
            I => \N__37051\
        );

    \I__9357\ : InMux
    port map (
            O => \N__37080\,
            I => \N__37051\
        );

    \I__9356\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37051\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__37072\,
            I => \N__37048\
        );

    \I__9354\ : Span4Mux_v
    port map (
            O => \N__37069\,
            I => \N__37045\
        );

    \I__9353\ : Span4Mux_v
    port map (
            O => \N__37066\,
            I => \N__37042\
        );

    \I__9352\ : Span4Mux_h
    port map (
            O => \N__37063\,
            I => \N__37039\
        );

    \I__9351\ : Span4Mux_v
    port map (
            O => \N__37060\,
            I => \N__37034\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__37051\,
            I => \N__37034\
        );

    \I__9349\ : Span4Mux_h
    port map (
            O => \N__37048\,
            I => \N__37031\
        );

    \I__9348\ : Span4Mux_h
    port map (
            O => \N__37045\,
            I => \N__37024\
        );

    \I__9347\ : Span4Mux_h
    port map (
            O => \N__37042\,
            I => \N__37024\
        );

    \I__9346\ : Span4Mux_h
    port map (
            O => \N__37039\,
            I => \N__37024\
        );

    \I__9345\ : Sp12to4
    port map (
            O => \N__37034\,
            I => \N__37021\
        );

    \I__9344\ : Span4Mux_h
    port map (
            O => \N__37031\,
            I => \N__37018\
        );

    \I__9343\ : Span4Mux_h
    port map (
            O => \N__37024\,
            I => \N__37015\
        );

    \I__9342\ : Odrv12
    port map (
            O => \N__37021\,
            I => \N_49\
        );

    \I__9341\ : Odrv4
    port map (
            O => \N__37018\,
            I => \N_49\
        );

    \I__9340\ : Odrv4
    port map (
            O => \N__37015\,
            I => \N_49\
        );

    \I__9339\ : IoInMux
    port map (
            O => \N__37008\,
            I => \N__37005\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__37005\,
            I => \N__37002\
        );

    \I__9337\ : Span4Mux_s2_h
    port map (
            O => \N__37002\,
            I => \N__36999\
        );

    \I__9336\ : Span4Mux_h
    port map (
            O => \N__36999\,
            I => \N__36996\
        );

    \I__9335\ : Sp12to4
    port map (
            O => \N__36996\,
            I => \N__36993\
        );

    \I__9334\ : Span12Mux_v
    port map (
            O => \N__36993\,
            I => \N__36989\
        );

    \I__9333\ : InMux
    port map (
            O => \N__36992\,
            I => \N__36986\
        );

    \I__9332\ : Odrv12
    port map (
            O => \N__36989\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__36986\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__9330\ : InMux
    port map (
            O => \N__36981\,
            I => \M_this_external_address_q_cry_6\
        );

    \I__9329\ : ClkMux
    port map (
            O => \N__36978\,
            I => \N__36582\
        );

    \I__9328\ : ClkMux
    port map (
            O => \N__36977\,
            I => \N__36582\
        );

    \I__9327\ : ClkMux
    port map (
            O => \N__36976\,
            I => \N__36582\
        );

    \I__9326\ : ClkMux
    port map (
            O => \N__36975\,
            I => \N__36582\
        );

    \I__9325\ : ClkMux
    port map (
            O => \N__36974\,
            I => \N__36582\
        );

    \I__9324\ : ClkMux
    port map (
            O => \N__36973\,
            I => \N__36582\
        );

    \I__9323\ : ClkMux
    port map (
            O => \N__36972\,
            I => \N__36582\
        );

    \I__9322\ : ClkMux
    port map (
            O => \N__36971\,
            I => \N__36582\
        );

    \I__9321\ : ClkMux
    port map (
            O => \N__36970\,
            I => \N__36582\
        );

    \I__9320\ : ClkMux
    port map (
            O => \N__36969\,
            I => \N__36582\
        );

    \I__9319\ : ClkMux
    port map (
            O => \N__36968\,
            I => \N__36582\
        );

    \I__9318\ : ClkMux
    port map (
            O => \N__36967\,
            I => \N__36582\
        );

    \I__9317\ : ClkMux
    port map (
            O => \N__36966\,
            I => \N__36582\
        );

    \I__9316\ : ClkMux
    port map (
            O => \N__36965\,
            I => \N__36582\
        );

    \I__9315\ : ClkMux
    port map (
            O => \N__36964\,
            I => \N__36582\
        );

    \I__9314\ : ClkMux
    port map (
            O => \N__36963\,
            I => \N__36582\
        );

    \I__9313\ : ClkMux
    port map (
            O => \N__36962\,
            I => \N__36582\
        );

    \I__9312\ : ClkMux
    port map (
            O => \N__36961\,
            I => \N__36582\
        );

    \I__9311\ : ClkMux
    port map (
            O => \N__36960\,
            I => \N__36582\
        );

    \I__9310\ : ClkMux
    port map (
            O => \N__36959\,
            I => \N__36582\
        );

    \I__9309\ : ClkMux
    port map (
            O => \N__36958\,
            I => \N__36582\
        );

    \I__9308\ : ClkMux
    port map (
            O => \N__36957\,
            I => \N__36582\
        );

    \I__9307\ : ClkMux
    port map (
            O => \N__36956\,
            I => \N__36582\
        );

    \I__9306\ : ClkMux
    port map (
            O => \N__36955\,
            I => \N__36582\
        );

    \I__9305\ : ClkMux
    port map (
            O => \N__36954\,
            I => \N__36582\
        );

    \I__9304\ : ClkMux
    port map (
            O => \N__36953\,
            I => \N__36582\
        );

    \I__9303\ : ClkMux
    port map (
            O => \N__36952\,
            I => \N__36582\
        );

    \I__9302\ : ClkMux
    port map (
            O => \N__36951\,
            I => \N__36582\
        );

    \I__9301\ : ClkMux
    port map (
            O => \N__36950\,
            I => \N__36582\
        );

    \I__9300\ : ClkMux
    port map (
            O => \N__36949\,
            I => \N__36582\
        );

    \I__9299\ : ClkMux
    port map (
            O => \N__36948\,
            I => \N__36582\
        );

    \I__9298\ : ClkMux
    port map (
            O => \N__36947\,
            I => \N__36582\
        );

    \I__9297\ : ClkMux
    port map (
            O => \N__36946\,
            I => \N__36582\
        );

    \I__9296\ : ClkMux
    port map (
            O => \N__36945\,
            I => \N__36582\
        );

    \I__9295\ : ClkMux
    port map (
            O => \N__36944\,
            I => \N__36582\
        );

    \I__9294\ : ClkMux
    port map (
            O => \N__36943\,
            I => \N__36582\
        );

    \I__9293\ : ClkMux
    port map (
            O => \N__36942\,
            I => \N__36582\
        );

    \I__9292\ : ClkMux
    port map (
            O => \N__36941\,
            I => \N__36582\
        );

    \I__9291\ : ClkMux
    port map (
            O => \N__36940\,
            I => \N__36582\
        );

    \I__9290\ : ClkMux
    port map (
            O => \N__36939\,
            I => \N__36582\
        );

    \I__9289\ : ClkMux
    port map (
            O => \N__36938\,
            I => \N__36582\
        );

    \I__9288\ : ClkMux
    port map (
            O => \N__36937\,
            I => \N__36582\
        );

    \I__9287\ : ClkMux
    port map (
            O => \N__36936\,
            I => \N__36582\
        );

    \I__9286\ : ClkMux
    port map (
            O => \N__36935\,
            I => \N__36582\
        );

    \I__9285\ : ClkMux
    port map (
            O => \N__36934\,
            I => \N__36582\
        );

    \I__9284\ : ClkMux
    port map (
            O => \N__36933\,
            I => \N__36582\
        );

    \I__9283\ : ClkMux
    port map (
            O => \N__36932\,
            I => \N__36582\
        );

    \I__9282\ : ClkMux
    port map (
            O => \N__36931\,
            I => \N__36582\
        );

    \I__9281\ : ClkMux
    port map (
            O => \N__36930\,
            I => \N__36582\
        );

    \I__9280\ : ClkMux
    port map (
            O => \N__36929\,
            I => \N__36582\
        );

    \I__9279\ : ClkMux
    port map (
            O => \N__36928\,
            I => \N__36582\
        );

    \I__9278\ : ClkMux
    port map (
            O => \N__36927\,
            I => \N__36582\
        );

    \I__9277\ : ClkMux
    port map (
            O => \N__36926\,
            I => \N__36582\
        );

    \I__9276\ : ClkMux
    port map (
            O => \N__36925\,
            I => \N__36582\
        );

    \I__9275\ : ClkMux
    port map (
            O => \N__36924\,
            I => \N__36582\
        );

    \I__9274\ : ClkMux
    port map (
            O => \N__36923\,
            I => \N__36582\
        );

    \I__9273\ : ClkMux
    port map (
            O => \N__36922\,
            I => \N__36582\
        );

    \I__9272\ : ClkMux
    port map (
            O => \N__36921\,
            I => \N__36582\
        );

    \I__9271\ : ClkMux
    port map (
            O => \N__36920\,
            I => \N__36582\
        );

    \I__9270\ : ClkMux
    port map (
            O => \N__36919\,
            I => \N__36582\
        );

    \I__9269\ : ClkMux
    port map (
            O => \N__36918\,
            I => \N__36582\
        );

    \I__9268\ : ClkMux
    port map (
            O => \N__36917\,
            I => \N__36582\
        );

    \I__9267\ : ClkMux
    port map (
            O => \N__36916\,
            I => \N__36582\
        );

    \I__9266\ : ClkMux
    port map (
            O => \N__36915\,
            I => \N__36582\
        );

    \I__9265\ : ClkMux
    port map (
            O => \N__36914\,
            I => \N__36582\
        );

    \I__9264\ : ClkMux
    port map (
            O => \N__36913\,
            I => \N__36582\
        );

    \I__9263\ : ClkMux
    port map (
            O => \N__36912\,
            I => \N__36582\
        );

    \I__9262\ : ClkMux
    port map (
            O => \N__36911\,
            I => \N__36582\
        );

    \I__9261\ : ClkMux
    port map (
            O => \N__36910\,
            I => \N__36582\
        );

    \I__9260\ : ClkMux
    port map (
            O => \N__36909\,
            I => \N__36582\
        );

    \I__9259\ : ClkMux
    port map (
            O => \N__36908\,
            I => \N__36582\
        );

    \I__9258\ : ClkMux
    port map (
            O => \N__36907\,
            I => \N__36582\
        );

    \I__9257\ : ClkMux
    port map (
            O => \N__36906\,
            I => \N__36582\
        );

    \I__9256\ : ClkMux
    port map (
            O => \N__36905\,
            I => \N__36582\
        );

    \I__9255\ : ClkMux
    port map (
            O => \N__36904\,
            I => \N__36582\
        );

    \I__9254\ : ClkMux
    port map (
            O => \N__36903\,
            I => \N__36582\
        );

    \I__9253\ : ClkMux
    port map (
            O => \N__36902\,
            I => \N__36582\
        );

    \I__9252\ : ClkMux
    port map (
            O => \N__36901\,
            I => \N__36582\
        );

    \I__9251\ : ClkMux
    port map (
            O => \N__36900\,
            I => \N__36582\
        );

    \I__9250\ : ClkMux
    port map (
            O => \N__36899\,
            I => \N__36582\
        );

    \I__9249\ : ClkMux
    port map (
            O => \N__36898\,
            I => \N__36582\
        );

    \I__9248\ : ClkMux
    port map (
            O => \N__36897\,
            I => \N__36582\
        );

    \I__9247\ : ClkMux
    port map (
            O => \N__36896\,
            I => \N__36582\
        );

    \I__9246\ : ClkMux
    port map (
            O => \N__36895\,
            I => \N__36582\
        );

    \I__9245\ : ClkMux
    port map (
            O => \N__36894\,
            I => \N__36582\
        );

    \I__9244\ : ClkMux
    port map (
            O => \N__36893\,
            I => \N__36582\
        );

    \I__9243\ : ClkMux
    port map (
            O => \N__36892\,
            I => \N__36582\
        );

    \I__9242\ : ClkMux
    port map (
            O => \N__36891\,
            I => \N__36582\
        );

    \I__9241\ : ClkMux
    port map (
            O => \N__36890\,
            I => \N__36582\
        );

    \I__9240\ : ClkMux
    port map (
            O => \N__36889\,
            I => \N__36582\
        );

    \I__9239\ : ClkMux
    port map (
            O => \N__36888\,
            I => \N__36582\
        );

    \I__9238\ : ClkMux
    port map (
            O => \N__36887\,
            I => \N__36582\
        );

    \I__9237\ : ClkMux
    port map (
            O => \N__36886\,
            I => \N__36582\
        );

    \I__9236\ : ClkMux
    port map (
            O => \N__36885\,
            I => \N__36582\
        );

    \I__9235\ : ClkMux
    port map (
            O => \N__36884\,
            I => \N__36582\
        );

    \I__9234\ : ClkMux
    port map (
            O => \N__36883\,
            I => \N__36582\
        );

    \I__9233\ : ClkMux
    port map (
            O => \N__36882\,
            I => \N__36582\
        );

    \I__9232\ : ClkMux
    port map (
            O => \N__36881\,
            I => \N__36582\
        );

    \I__9231\ : ClkMux
    port map (
            O => \N__36880\,
            I => \N__36582\
        );

    \I__9230\ : ClkMux
    port map (
            O => \N__36879\,
            I => \N__36582\
        );

    \I__9229\ : ClkMux
    port map (
            O => \N__36878\,
            I => \N__36582\
        );

    \I__9228\ : ClkMux
    port map (
            O => \N__36877\,
            I => \N__36582\
        );

    \I__9227\ : ClkMux
    port map (
            O => \N__36876\,
            I => \N__36582\
        );

    \I__9226\ : ClkMux
    port map (
            O => \N__36875\,
            I => \N__36582\
        );

    \I__9225\ : ClkMux
    port map (
            O => \N__36874\,
            I => \N__36582\
        );

    \I__9224\ : ClkMux
    port map (
            O => \N__36873\,
            I => \N__36582\
        );

    \I__9223\ : ClkMux
    port map (
            O => \N__36872\,
            I => \N__36582\
        );

    \I__9222\ : ClkMux
    port map (
            O => \N__36871\,
            I => \N__36582\
        );

    \I__9221\ : ClkMux
    port map (
            O => \N__36870\,
            I => \N__36582\
        );

    \I__9220\ : ClkMux
    port map (
            O => \N__36869\,
            I => \N__36582\
        );

    \I__9219\ : ClkMux
    port map (
            O => \N__36868\,
            I => \N__36582\
        );

    \I__9218\ : ClkMux
    port map (
            O => \N__36867\,
            I => \N__36582\
        );

    \I__9217\ : ClkMux
    port map (
            O => \N__36866\,
            I => \N__36582\
        );

    \I__9216\ : ClkMux
    port map (
            O => \N__36865\,
            I => \N__36582\
        );

    \I__9215\ : ClkMux
    port map (
            O => \N__36864\,
            I => \N__36582\
        );

    \I__9214\ : ClkMux
    port map (
            O => \N__36863\,
            I => \N__36582\
        );

    \I__9213\ : ClkMux
    port map (
            O => \N__36862\,
            I => \N__36582\
        );

    \I__9212\ : ClkMux
    port map (
            O => \N__36861\,
            I => \N__36582\
        );

    \I__9211\ : ClkMux
    port map (
            O => \N__36860\,
            I => \N__36582\
        );

    \I__9210\ : ClkMux
    port map (
            O => \N__36859\,
            I => \N__36582\
        );

    \I__9209\ : ClkMux
    port map (
            O => \N__36858\,
            I => \N__36582\
        );

    \I__9208\ : ClkMux
    port map (
            O => \N__36857\,
            I => \N__36582\
        );

    \I__9207\ : ClkMux
    port map (
            O => \N__36856\,
            I => \N__36582\
        );

    \I__9206\ : ClkMux
    port map (
            O => \N__36855\,
            I => \N__36582\
        );

    \I__9205\ : ClkMux
    port map (
            O => \N__36854\,
            I => \N__36582\
        );

    \I__9204\ : ClkMux
    port map (
            O => \N__36853\,
            I => \N__36582\
        );

    \I__9203\ : ClkMux
    port map (
            O => \N__36852\,
            I => \N__36582\
        );

    \I__9202\ : ClkMux
    port map (
            O => \N__36851\,
            I => \N__36582\
        );

    \I__9201\ : ClkMux
    port map (
            O => \N__36850\,
            I => \N__36582\
        );

    \I__9200\ : ClkMux
    port map (
            O => \N__36849\,
            I => \N__36582\
        );

    \I__9199\ : ClkMux
    port map (
            O => \N__36848\,
            I => \N__36582\
        );

    \I__9198\ : ClkMux
    port map (
            O => \N__36847\,
            I => \N__36582\
        );

    \I__9197\ : GlobalMux
    port map (
            O => \N__36582\,
            I => \N__36579\
        );

    \I__9196\ : gio2CtrlBuf
    port map (
            O => \N__36579\,
            I => clk_0_c_g
        );

    \I__9195\ : CEMux
    port map (
            O => \N__36576\,
            I => \N__36571\
        );

    \I__9194\ : CEMux
    port map (
            O => \N__36575\,
            I => \N__36568\
        );

    \I__9193\ : CEMux
    port map (
            O => \N__36574\,
            I => \N__36565\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__36571\,
            I => \N__36562\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__36568\,
            I => \N__36557\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__36565\,
            I => \N__36554\
        );

    \I__9189\ : Span4Mux_h
    port map (
            O => \N__36562\,
            I => \N__36551\
        );

    \I__9188\ : CEMux
    port map (
            O => \N__36561\,
            I => \N__36548\
        );

    \I__9187\ : CEMux
    port map (
            O => \N__36560\,
            I => \N__36545\
        );

    \I__9186\ : Span4Mux_v
    port map (
            O => \N__36557\,
            I => \N__36540\
        );

    \I__9185\ : Span4Mux_v
    port map (
            O => \N__36554\,
            I => \N__36540\
        );

    \I__9184\ : Span4Mux_h
    port map (
            O => \N__36551\,
            I => \N__36535\
        );

    \I__9183\ : LocalMux
    port map (
            O => \N__36548\,
            I => \N__36535\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__36545\,
            I => \N__36532\
        );

    \I__9181\ : Odrv4
    port map (
            O => \N__36540\,
            I => \N_47\
        );

    \I__9180\ : Odrv4
    port map (
            O => \N__36535\,
            I => \N_47\
        );

    \I__9179\ : Odrv12
    port map (
            O => \N__36532\,
            I => \N_47\
        );

    \I__9178\ : IoInMux
    port map (
            O => \N__36525\,
            I => \N__36522\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__36522\,
            I => \N__36519\
        );

    \I__9176\ : IoSpan4Mux
    port map (
            O => \N__36519\,
            I => \N__36516\
        );

    \I__9175\ : Span4Mux_s3_v
    port map (
            O => \N__36516\,
            I => \N__36513\
        );

    \I__9174\ : Span4Mux_h
    port map (
            O => \N__36513\,
            I => \N__36509\
        );

    \I__9173\ : InMux
    port map (
            O => \N__36512\,
            I => \N__36506\
        );

    \I__9172\ : Span4Mux_v
    port map (
            O => \N__36509\,
            I => \N__36503\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__36506\,
            I => \N__36500\
        );

    \I__9170\ : Odrv4
    port map (
            O => \N__36503\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__9169\ : Odrv4
    port map (
            O => \N__36500\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__9168\ : InMux
    port map (
            O => \N__36495\,
            I => \N__36492\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__36492\,
            I => \N__36489\
        );

    \I__9166\ : Odrv12
    port map (
            O => \N__36489\,
            I => \M_this_external_address_q_s_8\
        );

    \I__9165\ : InMux
    port map (
            O => \N__36486\,
            I => \bfn_26_22_0_\
        );

    \I__9164\ : IoInMux
    port map (
            O => \N__36483\,
            I => \N__36480\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__36480\,
            I => \N__36477\
        );

    \I__9162\ : IoSpan4Mux
    port map (
            O => \N__36477\,
            I => \N__36473\
        );

    \I__9161\ : InMux
    port map (
            O => \N__36476\,
            I => \N__36470\
        );

    \I__9160\ : Span4Mux_s1_v
    port map (
            O => \N__36473\,
            I => \N__36467\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__36470\,
            I => \N__36464\
        );

    \I__9158\ : Sp12to4
    port map (
            O => \N__36467\,
            I => \N__36461\
        );

    \I__9157\ : Span4Mux_h
    port map (
            O => \N__36464\,
            I => \N__36458\
        );

    \I__9156\ : Odrv12
    port map (
            O => \N__36461\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__9155\ : Odrv4
    port map (
            O => \N__36458\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__9154\ : InMux
    port map (
            O => \N__36453\,
            I => \N__36450\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__36450\,
            I => \N__36447\
        );

    \I__9152\ : Span4Mux_h
    port map (
            O => \N__36447\,
            I => \N__36444\
        );

    \I__9151\ : Odrv4
    port map (
            O => \N__36444\,
            I => \M_this_external_address_q_s_9\
        );

    \I__9150\ : InMux
    port map (
            O => \N__36441\,
            I => \M_this_external_address_q_cry_8\
        );

    \I__9149\ : IoInMux
    port map (
            O => \N__36438\,
            I => \N__36435\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__36435\,
            I => \N__36432\
        );

    \I__9147\ : IoSpan4Mux
    port map (
            O => \N__36432\,
            I => \N__36429\
        );

    \I__9146\ : Span4Mux_s3_v
    port map (
            O => \N__36429\,
            I => \N__36425\
        );

    \I__9145\ : InMux
    port map (
            O => \N__36428\,
            I => \N__36422\
        );

    \I__9144\ : Span4Mux_v
    port map (
            O => \N__36425\,
            I => \N__36419\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__36422\,
            I => \N__36416\
        );

    \I__9142\ : Odrv4
    port map (
            O => \N__36419\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__9141\ : Odrv4
    port map (
            O => \N__36416\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__9140\ : InMux
    port map (
            O => \N__36411\,
            I => \N__36408\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__36408\,
            I => \N__36405\
        );

    \I__9138\ : Odrv4
    port map (
            O => \N__36405\,
            I => \M_this_external_address_q_s_10\
        );

    \I__9137\ : InMux
    port map (
            O => \N__36402\,
            I => \M_this_external_address_q_cry_9\
        );

    \I__9136\ : IoInMux
    port map (
            O => \N__36399\,
            I => \N__36396\
        );

    \I__9135\ : LocalMux
    port map (
            O => \N__36396\,
            I => \N__36393\
        );

    \I__9134\ : Span4Mux_s2_v
    port map (
            O => \N__36393\,
            I => \N__36390\
        );

    \I__9133\ : Span4Mux_v
    port map (
            O => \N__36390\,
            I => \N__36387\
        );

    \I__9132\ : Span4Mux_v
    port map (
            O => \N__36387\,
            I => \N__36383\
        );

    \I__9131\ : InMux
    port map (
            O => \N__36386\,
            I => \N__36380\
        );

    \I__9130\ : Sp12to4
    port map (
            O => \N__36383\,
            I => \N__36375\
        );

    \I__9129\ : LocalMux
    port map (
            O => \N__36380\,
            I => \N__36375\
        );

    \I__9128\ : Odrv12
    port map (
            O => \N__36375\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__9127\ : InMux
    port map (
            O => \N__36372\,
            I => \N__36369\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__36369\,
            I => \N__36366\
        );

    \I__9125\ : Odrv4
    port map (
            O => \N__36366\,
            I => \M_this_external_address_q_s_11\
        );

    \I__9124\ : InMux
    port map (
            O => \N__36363\,
            I => \M_this_external_address_q_cry_10\
        );

    \I__9123\ : InMux
    port map (
            O => \N__36360\,
            I => \N__36357\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__36357\,
            I => \N__36352\
        );

    \I__9121\ : CascadeMux
    port map (
            O => \N__36356\,
            I => \N__36349\
        );

    \I__9120\ : InMux
    port map (
            O => \N__36355\,
            I => \N__36345\
        );

    \I__9119\ : Span4Mux_v
    port map (
            O => \N__36352\,
            I => \N__36341\
        );

    \I__9118\ : InMux
    port map (
            O => \N__36349\,
            I => \N__36338\
        );

    \I__9117\ : CascadeMux
    port map (
            O => \N__36348\,
            I => \N__36335\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__36345\,
            I => \N__36329\
        );

    \I__9115\ : InMux
    port map (
            O => \N__36344\,
            I => \N__36326\
        );

    \I__9114\ : Span4Mux_h
    port map (
            O => \N__36341\,
            I => \N__36318\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__36338\,
            I => \N__36318\
        );

    \I__9112\ : InMux
    port map (
            O => \N__36335\,
            I => \N__36315\
        );

    \I__9111\ : InMux
    port map (
            O => \N__36334\,
            I => \N__36310\
        );

    \I__9110\ : InMux
    port map (
            O => \N__36333\,
            I => \N__36307\
        );

    \I__9109\ : CascadeMux
    port map (
            O => \N__36332\,
            I => \N__36304\
        );

    \I__9108\ : Span4Mux_v
    port map (
            O => \N__36329\,
            I => \N__36297\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__36326\,
            I => \N__36294\
        );

    \I__9106\ : InMux
    port map (
            O => \N__36325\,
            I => \N__36291\
        );

    \I__9105\ : InMux
    port map (
            O => \N__36324\,
            I => \N__36288\
        );

    \I__9104\ : InMux
    port map (
            O => \N__36323\,
            I => \N__36285\
        );

    \I__9103\ : Span4Mux_v
    port map (
            O => \N__36318\,
            I => \N__36281\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__36315\,
            I => \N__36278\
        );

    \I__9101\ : InMux
    port map (
            O => \N__36314\,
            I => \N__36275\
        );

    \I__9100\ : InMux
    port map (
            O => \N__36313\,
            I => \N__36272\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__36310\,
            I => \N__36267\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__36307\,
            I => \N__36267\
        );

    \I__9097\ : InMux
    port map (
            O => \N__36304\,
            I => \N__36260\
        );

    \I__9096\ : InMux
    port map (
            O => \N__36303\,
            I => \N__36260\
        );

    \I__9095\ : InMux
    port map (
            O => \N__36302\,
            I => \N__36260\
        );

    \I__9094\ : InMux
    port map (
            O => \N__36301\,
            I => \N__36256\
        );

    \I__9093\ : InMux
    port map (
            O => \N__36300\,
            I => \N__36253\
        );

    \I__9092\ : Span4Mux_v
    port map (
            O => \N__36297\,
            I => \N__36249\
        );

    \I__9091\ : Span4Mux_v
    port map (
            O => \N__36294\,
            I => \N__36244\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__36291\,
            I => \N__36244\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__36288\,
            I => \N__36241\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__36285\,
            I => \N__36238\
        );

    \I__9087\ : InMux
    port map (
            O => \N__36284\,
            I => \N__36235\
        );

    \I__9086\ : Span4Mux_h
    port map (
            O => \N__36281\,
            I => \N__36222\
        );

    \I__9085\ : Span4Mux_v
    port map (
            O => \N__36278\,
            I => \N__36222\
        );

    \I__9084\ : LocalMux
    port map (
            O => \N__36275\,
            I => \N__36222\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__36272\,
            I => \N__36222\
        );

    \I__9082\ : Span4Mux_v
    port map (
            O => \N__36267\,
            I => \N__36222\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__36260\,
            I => \N__36222\
        );

    \I__9080\ : InMux
    port map (
            O => \N__36259\,
            I => \N__36219\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__36256\,
            I => \N__36214\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__36253\,
            I => \N__36214\
        );

    \I__9077\ : InMux
    port map (
            O => \N__36252\,
            I => \N__36211\
        );

    \I__9076\ : Span4Mux_v
    port map (
            O => \N__36249\,
            I => \N__36204\
        );

    \I__9075\ : Span4Mux_v
    port map (
            O => \N__36244\,
            I => \N__36204\
        );

    \I__9074\ : Span4Mux_v
    port map (
            O => \N__36241\,
            I => \N__36204\
        );

    \I__9073\ : Span4Mux_h
    port map (
            O => \N__36238\,
            I => \N__36199\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__36235\,
            I => \N__36199\
        );

    \I__9071\ : Span4Mux_v
    port map (
            O => \N__36222\,
            I => \N__36196\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__36219\,
            I => \N__36193\
        );

    \I__9069\ : Span12Mux_h
    port map (
            O => \N__36214\,
            I => \N__36190\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__36211\,
            I => \N__36187\
        );

    \I__9067\ : Span4Mux_h
    port map (
            O => \N__36204\,
            I => \N__36182\
        );

    \I__9066\ : Span4Mux_v
    port map (
            O => \N__36199\,
            I => \N__36182\
        );

    \I__9065\ : Span4Mux_h
    port map (
            O => \N__36196\,
            I => \N__36177\
        );

    \I__9064\ : Span4Mux_v
    port map (
            O => \N__36193\,
            I => \N__36177\
        );

    \I__9063\ : Span12Mux_v
    port map (
            O => \N__36190\,
            I => \N__36174\
        );

    \I__9062\ : Span12Mux_v
    port map (
            O => \N__36187\,
            I => \N__36169\
        );

    \I__9061\ : Sp12to4
    port map (
            O => \N__36182\,
            I => \N__36169\
        );

    \I__9060\ : Span4Mux_h
    port map (
            O => \N__36177\,
            I => \N__36166\
        );

    \I__9059\ : Odrv12
    port map (
            O => \N__36174\,
            I => port_data_c_5
        );

    \I__9058\ : Odrv12
    port map (
            O => \N__36169\,
            I => port_data_c_5
        );

    \I__9057\ : Odrv4
    port map (
            O => \N__36166\,
            I => port_data_c_5
        );

    \I__9056\ : InMux
    port map (
            O => \N__36159\,
            I => \N__36156\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__36156\,
            I => \N__36153\
        );

    \I__9054\ : Span4Mux_h
    port map (
            O => \N__36153\,
            I => \N__36150\
        );

    \I__9053\ : Odrv4
    port map (
            O => \N__36150\,
            I => \M_this_data_tmp_qZ0Z_13\
        );

    \I__9052\ : CEMux
    port map (
            O => \N__36147\,
            I => \N__36144\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__36144\,
            I => \N__36138\
        );

    \I__9050\ : CEMux
    port map (
            O => \N__36143\,
            I => \N__36135\
        );

    \I__9049\ : CEMux
    port map (
            O => \N__36142\,
            I => \N__36132\
        );

    \I__9048\ : CEMux
    port map (
            O => \N__36141\,
            I => \N__36129\
        );

    \I__9047\ : Span4Mux_h
    port map (
            O => \N__36138\,
            I => \N__36119\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__36135\,
            I => \N__36119\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__36132\,
            I => \N__36119\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__36129\,
            I => \N__36119\
        );

    \I__9043\ : CEMux
    port map (
            O => \N__36128\,
            I => \N__36116\
        );

    \I__9042\ : Span4Mux_v
    port map (
            O => \N__36119\,
            I => \N__36113\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__36116\,
            I => \N__36110\
        );

    \I__9040\ : Odrv4
    port map (
            O => \N__36113\,
            I => \N_1404_0\
        );

    \I__9039\ : Odrv12
    port map (
            O => \N__36110\,
            I => \N_1404_0\
        );

    \I__9038\ : InMux
    port map (
            O => \N__36105\,
            I => \N__36083\
        );

    \I__9037\ : InMux
    port map (
            O => \N__36104\,
            I => \N__36080\
        );

    \I__9036\ : InMux
    port map (
            O => \N__36103\,
            I => \N__36077\
        );

    \I__9035\ : InMux
    port map (
            O => \N__36102\,
            I => \N__36074\
        );

    \I__9034\ : InMux
    port map (
            O => \N__36101\,
            I => \N__36071\
        );

    \I__9033\ : InMux
    port map (
            O => \N__36100\,
            I => \N__36068\
        );

    \I__9032\ : InMux
    port map (
            O => \N__36099\,
            I => \N__36065\
        );

    \I__9031\ : InMux
    port map (
            O => \N__36098\,
            I => \N__36062\
        );

    \I__9030\ : InMux
    port map (
            O => \N__36097\,
            I => \N__36059\
        );

    \I__9029\ : InMux
    port map (
            O => \N__36096\,
            I => \N__36056\
        );

    \I__9028\ : InMux
    port map (
            O => \N__36095\,
            I => \N__36053\
        );

    \I__9027\ : InMux
    port map (
            O => \N__36094\,
            I => \N__36048\
        );

    \I__9026\ : InMux
    port map (
            O => \N__36093\,
            I => \N__36048\
        );

    \I__9025\ : InMux
    port map (
            O => \N__36092\,
            I => \N__36045\
        );

    \I__9024\ : InMux
    port map (
            O => \N__36091\,
            I => \N__36042\
        );

    \I__9023\ : InMux
    port map (
            O => \N__36090\,
            I => \N__36035\
        );

    \I__9022\ : InMux
    port map (
            O => \N__36089\,
            I => \N__36035\
        );

    \I__9021\ : InMux
    port map (
            O => \N__36088\,
            I => \N__36035\
        );

    \I__9020\ : InMux
    port map (
            O => \N__36087\,
            I => \N__36030\
        );

    \I__9019\ : InMux
    port map (
            O => \N__36086\,
            I => \N__36030\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__36083\,
            I => \N__36002\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__36080\,
            I => \N__35999\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__36077\,
            I => \N__35996\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__36074\,
            I => \N__35993\
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__36071\,
            I => \N__35990\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__36068\,
            I => \N__35987\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__36065\,
            I => \N__35984\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__36062\,
            I => \N__35981\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__36059\,
            I => \N__35978\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__36056\,
            I => \N__35975\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__36053\,
            I => \N__35972\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__36048\,
            I => \N__35969\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__36045\,
            I => \N__35966\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__36042\,
            I => \N__35963\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__36035\,
            I => \N__35960\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__36030\,
            I => \N__35957\
        );

    \I__9002\ : SRMux
    port map (
            O => \N__36029\,
            I => \N__35874\
        );

    \I__9001\ : SRMux
    port map (
            O => \N__36028\,
            I => \N__35874\
        );

    \I__9000\ : SRMux
    port map (
            O => \N__36027\,
            I => \N__35874\
        );

    \I__8999\ : SRMux
    port map (
            O => \N__36026\,
            I => \N__35874\
        );

    \I__8998\ : SRMux
    port map (
            O => \N__36025\,
            I => \N__35874\
        );

    \I__8997\ : SRMux
    port map (
            O => \N__36024\,
            I => \N__35874\
        );

    \I__8996\ : SRMux
    port map (
            O => \N__36023\,
            I => \N__35874\
        );

    \I__8995\ : SRMux
    port map (
            O => \N__36022\,
            I => \N__35874\
        );

    \I__8994\ : SRMux
    port map (
            O => \N__36021\,
            I => \N__35874\
        );

    \I__8993\ : SRMux
    port map (
            O => \N__36020\,
            I => \N__35874\
        );

    \I__8992\ : SRMux
    port map (
            O => \N__36019\,
            I => \N__35874\
        );

    \I__8991\ : SRMux
    port map (
            O => \N__36018\,
            I => \N__35874\
        );

    \I__8990\ : SRMux
    port map (
            O => \N__36017\,
            I => \N__35874\
        );

    \I__8989\ : SRMux
    port map (
            O => \N__36016\,
            I => \N__35874\
        );

    \I__8988\ : SRMux
    port map (
            O => \N__36015\,
            I => \N__35874\
        );

    \I__8987\ : SRMux
    port map (
            O => \N__36014\,
            I => \N__35874\
        );

    \I__8986\ : SRMux
    port map (
            O => \N__36013\,
            I => \N__35874\
        );

    \I__8985\ : SRMux
    port map (
            O => \N__36012\,
            I => \N__35874\
        );

    \I__8984\ : SRMux
    port map (
            O => \N__36011\,
            I => \N__35874\
        );

    \I__8983\ : SRMux
    port map (
            O => \N__36010\,
            I => \N__35874\
        );

    \I__8982\ : SRMux
    port map (
            O => \N__36009\,
            I => \N__35874\
        );

    \I__8981\ : SRMux
    port map (
            O => \N__36008\,
            I => \N__35874\
        );

    \I__8980\ : SRMux
    port map (
            O => \N__36007\,
            I => \N__35874\
        );

    \I__8979\ : SRMux
    port map (
            O => \N__36006\,
            I => \N__35874\
        );

    \I__8978\ : SRMux
    port map (
            O => \N__36005\,
            I => \N__35874\
        );

    \I__8977\ : Glb2LocalMux
    port map (
            O => \N__36002\,
            I => \N__35874\
        );

    \I__8976\ : Glb2LocalMux
    port map (
            O => \N__35999\,
            I => \N__35874\
        );

    \I__8975\ : Glb2LocalMux
    port map (
            O => \N__35996\,
            I => \N__35874\
        );

    \I__8974\ : Glb2LocalMux
    port map (
            O => \N__35993\,
            I => \N__35874\
        );

    \I__8973\ : Glb2LocalMux
    port map (
            O => \N__35990\,
            I => \N__35874\
        );

    \I__8972\ : Glb2LocalMux
    port map (
            O => \N__35987\,
            I => \N__35874\
        );

    \I__8971\ : Glb2LocalMux
    port map (
            O => \N__35984\,
            I => \N__35874\
        );

    \I__8970\ : Glb2LocalMux
    port map (
            O => \N__35981\,
            I => \N__35874\
        );

    \I__8969\ : Glb2LocalMux
    port map (
            O => \N__35978\,
            I => \N__35874\
        );

    \I__8968\ : Glb2LocalMux
    port map (
            O => \N__35975\,
            I => \N__35874\
        );

    \I__8967\ : Glb2LocalMux
    port map (
            O => \N__35972\,
            I => \N__35874\
        );

    \I__8966\ : Glb2LocalMux
    port map (
            O => \N__35969\,
            I => \N__35874\
        );

    \I__8965\ : Glb2LocalMux
    port map (
            O => \N__35966\,
            I => \N__35874\
        );

    \I__8964\ : Glb2LocalMux
    port map (
            O => \N__35963\,
            I => \N__35874\
        );

    \I__8963\ : Glb2LocalMux
    port map (
            O => \N__35960\,
            I => \N__35874\
        );

    \I__8962\ : Glb2LocalMux
    port map (
            O => \N__35957\,
            I => \N__35874\
        );

    \I__8961\ : GlobalMux
    port map (
            O => \N__35874\,
            I => \N__35871\
        );

    \I__8960\ : gio2CtrlBuf
    port map (
            O => \N__35871\,
            I => \M_this_reset_cond_out_g_0\
        );

    \I__8959\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35865\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__35865\,
            I => \N__35860\
        );

    \I__8957\ : InMux
    port map (
            O => \N__35864\,
            I => \N__35857\
        );

    \I__8956\ : CascadeMux
    port map (
            O => \N__35863\,
            I => \N__35854\
        );

    \I__8955\ : Span4Mux_h
    port map (
            O => \N__35860\,
            I => \N__35849\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__35857\,
            I => \N__35849\
        );

    \I__8953\ : InMux
    port map (
            O => \N__35854\,
            I => \N__35843\
        );

    \I__8952\ : Span4Mux_h
    port map (
            O => \N__35849\,
            I => \N__35840\
        );

    \I__8951\ : InMux
    port map (
            O => \N__35848\,
            I => \N__35835\
        );

    \I__8950\ : CascadeMux
    port map (
            O => \N__35847\,
            I => \N__35832\
        );

    \I__8949\ : CascadeMux
    port map (
            O => \N__35846\,
            I => \N__35827\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__35843\,
            I => \N__35823\
        );

    \I__8947\ : Span4Mux_v
    port map (
            O => \N__35840\,
            I => \N__35820\
        );

    \I__8946\ : InMux
    port map (
            O => \N__35839\,
            I => \N__35817\
        );

    \I__8945\ : InMux
    port map (
            O => \N__35838\,
            I => \N__35814\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__35835\,
            I => \N__35811\
        );

    \I__8943\ : InMux
    port map (
            O => \N__35832\,
            I => \N__35808\
        );

    \I__8942\ : CascadeMux
    port map (
            O => \N__35831\,
            I => \N__35805\
        );

    \I__8941\ : InMux
    port map (
            O => \N__35830\,
            I => \N__35802\
        );

    \I__8940\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35797\
        );

    \I__8939\ : InMux
    port map (
            O => \N__35826\,
            I => \N__35797\
        );

    \I__8938\ : Span4Mux_v
    port map (
            O => \N__35823\,
            I => \N__35794\
        );

    \I__8937\ : Span4Mux_v
    port map (
            O => \N__35820\,
            I => \N__35791\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__35817\,
            I => \N__35788\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__35814\,
            I => \N__35785\
        );

    \I__8934\ : Span4Mux_v
    port map (
            O => \N__35811\,
            I => \N__35782\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__35808\,
            I => \N__35779\
        );

    \I__8932\ : InMux
    port map (
            O => \N__35805\,
            I => \N__35776\
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__35802\,
            I => \N__35773\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__35797\,
            I => \N__35770\
        );

    \I__8929\ : Span4Mux_h
    port map (
            O => \N__35794\,
            I => \N__35767\
        );

    \I__8928\ : Span4Mux_v
    port map (
            O => \N__35791\,
            I => \N__35762\
        );

    \I__8927\ : Span4Mux_h
    port map (
            O => \N__35788\,
            I => \N__35762\
        );

    \I__8926\ : Span4Mux_h
    port map (
            O => \N__35785\,
            I => \N__35759\
        );

    \I__8925\ : Span4Mux_v
    port map (
            O => \N__35782\,
            I => \N__35754\
        );

    \I__8924\ : Span4Mux_h
    port map (
            O => \N__35779\,
            I => \N__35754\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__35776\,
            I => \N__35751\
        );

    \I__8922\ : Span4Mux_h
    port map (
            O => \N__35773\,
            I => \N__35746\
        );

    \I__8921\ : Span4Mux_v
    port map (
            O => \N__35770\,
            I => \N__35746\
        );

    \I__8920\ : Span4Mux_h
    port map (
            O => \N__35767\,
            I => \N__35741\
        );

    \I__8919\ : Span4Mux_v
    port map (
            O => \N__35762\,
            I => \N__35741\
        );

    \I__8918\ : Sp12to4
    port map (
            O => \N__35759\,
            I => \N__35738\
        );

    \I__8917\ : Span4Mux_h
    port map (
            O => \N__35754\,
            I => \N__35735\
        );

    \I__8916\ : Span12Mux_v
    port map (
            O => \N__35751\,
            I => \N__35730\
        );

    \I__8915\ : Sp12to4
    port map (
            O => \N__35746\,
            I => \N__35730\
        );

    \I__8914\ : Span4Mux_v
    port map (
            O => \N__35741\,
            I => \N__35727\
        );

    \I__8913\ : Span12Mux_v
    port map (
            O => \N__35738\,
            I => \N__35722\
        );

    \I__8912\ : Sp12to4
    port map (
            O => \N__35735\,
            I => \N__35722\
        );

    \I__8911\ : Span12Mux_h
    port map (
            O => \N__35730\,
            I => \N__35719\
        );

    \I__8910\ : IoSpan4Mux
    port map (
            O => \N__35727\,
            I => \N__35716\
        );

    \I__8909\ : Odrv12
    port map (
            O => \N__35722\,
            I => port_data_c_3
        );

    \I__8908\ : Odrv12
    port map (
            O => \N__35719\,
            I => port_data_c_3
        );

    \I__8907\ : Odrv4
    port map (
            O => \N__35716\,
            I => port_data_c_3
        );

    \I__8906\ : CEMux
    port map (
            O => \N__35709\,
            I => \N__35685\
        );

    \I__8905\ : CEMux
    port map (
            O => \N__35708\,
            I => \N__35682\
        );

    \I__8904\ : InMux
    port map (
            O => \N__35707\,
            I => \N__35679\
        );

    \I__8903\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35674\
        );

    \I__8902\ : InMux
    port map (
            O => \N__35705\,
            I => \N__35674\
        );

    \I__8901\ : InMux
    port map (
            O => \N__35704\,
            I => \N__35667\
        );

    \I__8900\ : InMux
    port map (
            O => \N__35703\,
            I => \N__35667\
        );

    \I__8899\ : InMux
    port map (
            O => \N__35702\,
            I => \N__35667\
        );

    \I__8898\ : InMux
    port map (
            O => \N__35701\,
            I => \N__35658\
        );

    \I__8897\ : InMux
    port map (
            O => \N__35700\,
            I => \N__35658\
        );

    \I__8896\ : InMux
    port map (
            O => \N__35699\,
            I => \N__35658\
        );

    \I__8895\ : InMux
    port map (
            O => \N__35698\,
            I => \N__35658\
        );

    \I__8894\ : InMux
    port map (
            O => \N__35697\,
            I => \N__35645\
        );

    \I__8893\ : InMux
    port map (
            O => \N__35696\,
            I => \N__35645\
        );

    \I__8892\ : InMux
    port map (
            O => \N__35695\,
            I => \N__35645\
        );

    \I__8891\ : InMux
    port map (
            O => \N__35694\,
            I => \N__35645\
        );

    \I__8890\ : InMux
    port map (
            O => \N__35693\,
            I => \N__35645\
        );

    \I__8889\ : InMux
    port map (
            O => \N__35692\,
            I => \N__35645\
        );

    \I__8888\ : InMux
    port map (
            O => \N__35691\,
            I => \N__35638\
        );

    \I__8887\ : InMux
    port map (
            O => \N__35690\,
            I => \N__35631\
        );

    \I__8886\ : InMux
    port map (
            O => \N__35689\,
            I => \N__35631\
        );

    \I__8885\ : InMux
    port map (
            O => \N__35688\,
            I => \N__35631\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__35685\,
            I => \N__35622\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__35682\,
            I => \N__35619\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__35679\,
            I => \N__35616\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__35674\,
            I => \N__35609\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__35667\,
            I => \N__35609\
        );

    \I__8879\ : LocalMux
    port map (
            O => \N__35658\,
            I => \N__35609\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__35645\,
            I => \N__35606\
        );

    \I__8877\ : InMux
    port map (
            O => \N__35644\,
            I => \N__35601\
        );

    \I__8876\ : InMux
    port map (
            O => \N__35643\,
            I => \N__35601\
        );

    \I__8875\ : InMux
    port map (
            O => \N__35642\,
            I => \N__35598\
        );

    \I__8874\ : InMux
    port map (
            O => \N__35641\,
            I => \N__35595\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__35638\,
            I => \N__35592\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__35631\,
            I => \N__35589\
        );

    \I__8871\ : InMux
    port map (
            O => \N__35630\,
            I => \N__35584\
        );

    \I__8870\ : InMux
    port map (
            O => \N__35629\,
            I => \N__35584\
        );

    \I__8869\ : InMux
    port map (
            O => \N__35628\,
            I => \N__35577\
        );

    \I__8868\ : InMux
    port map (
            O => \N__35627\,
            I => \N__35577\
        );

    \I__8867\ : InMux
    port map (
            O => \N__35626\,
            I => \N__35577\
        );

    \I__8866\ : InMux
    port map (
            O => \N__35625\,
            I => \N__35574\
        );

    \I__8865\ : Span4Mux_v
    port map (
            O => \N__35622\,
            I => \N__35571\
        );

    \I__8864\ : Span4Mux_h
    port map (
            O => \N__35619\,
            I => \N__35568\
        );

    \I__8863\ : Span4Mux_h
    port map (
            O => \N__35616\,
            I => \N__35559\
        );

    \I__8862\ : Span4Mux_v
    port map (
            O => \N__35609\,
            I => \N__35559\
        );

    \I__8861\ : Span4Mux_h
    port map (
            O => \N__35606\,
            I => \N__35559\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__35601\,
            I => \N__35559\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__35598\,
            I => \N__35554\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__35595\,
            I => \N__35554\
        );

    \I__8857\ : Span4Mux_h
    port map (
            O => \N__35592\,
            I => \N__35545\
        );

    \I__8856\ : Span4Mux_h
    port map (
            O => \N__35589\,
            I => \N__35545\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__35584\,
            I => \N__35545\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__35577\,
            I => \N__35545\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__35574\,
            I => \N__35542\
        );

    \I__8852\ : Span4Mux_v
    port map (
            O => \N__35571\,
            I => \N__35535\
        );

    \I__8851\ : Span4Mux_v
    port map (
            O => \N__35568\,
            I => \N__35535\
        );

    \I__8850\ : Span4Mux_v
    port map (
            O => \N__35559\,
            I => \N__35532\
        );

    \I__8849\ : Span4Mux_h
    port map (
            O => \N__35554\,
            I => \N__35525\
        );

    \I__8848\ : Span4Mux_v
    port map (
            O => \N__35545\,
            I => \N__35525\
        );

    \I__8847\ : Span4Mux_h
    port map (
            O => \N__35542\,
            I => \N__35525\
        );

    \I__8846\ : InMux
    port map (
            O => \N__35541\,
            I => \N__35520\
        );

    \I__8845\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35520\
        );

    \I__8844\ : Odrv4
    port map (
            O => \N__35535\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__8843\ : Odrv4
    port map (
            O => \N__35532\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__8842\ : Odrv4
    port map (
            O => \N__35525\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__35520\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__8840\ : InMux
    port map (
            O => \N__35511\,
            I => \N__35508\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__35508\,
            I => \N__35505\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__35505\,
            I => \M_this_oam_ram_write_data_27\
        );

    \I__8837\ : InMux
    port map (
            O => \N__35502\,
            I => \N__35499\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__35499\,
            I => \N__35496\
        );

    \I__8835\ : Odrv4
    port map (
            O => \N__35496\,
            I => \M_this_external_address_q_3_0_13\
        );

    \I__8834\ : InMux
    port map (
            O => \N__35493\,
            I => \N__35490\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__35490\,
            I => \N__35487\
        );

    \I__8832\ : Odrv4
    port map (
            O => \N__35487\,
            I => \N_312_0\
        );

    \I__8831\ : IoInMux
    port map (
            O => \N__35484\,
            I => \N__35481\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__35481\,
            I => \N__35478\
        );

    \I__8829\ : Span4Mux_s3_v
    port map (
            O => \N__35478\,
            I => \N__35475\
        );

    \I__8828\ : Sp12to4
    port map (
            O => \N__35475\,
            I => \N__35472\
        );

    \I__8827\ : Span12Mux_h
    port map (
            O => \N__35472\,
            I => \N__35468\
        );

    \I__8826\ : InMux
    port map (
            O => \N__35471\,
            I => \N__35465\
        );

    \I__8825\ : Odrv12
    port map (
            O => \N__35468\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__35465\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__8823\ : InMux
    port map (
            O => \N__35460\,
            I => \bfn_26_21_0_\
        );

    \I__8822\ : IoInMux
    port map (
            O => \N__35457\,
            I => \N__35454\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__35454\,
            I => \N__35451\
        );

    \I__8820\ : Span12Mux_s2_v
    port map (
            O => \N__35451\,
            I => \N__35447\
        );

    \I__8819\ : InMux
    port map (
            O => \N__35450\,
            I => \N__35444\
        );

    \I__8818\ : Odrv12
    port map (
            O => \N__35447\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__35444\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__8816\ : InMux
    port map (
            O => \N__35439\,
            I => \M_this_external_address_q_cry_0\
        );

    \I__8815\ : IoInMux
    port map (
            O => \N__35436\,
            I => \N__35433\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__35433\,
            I => \N__35430\
        );

    \I__8813\ : Span4Mux_s1_v
    port map (
            O => \N__35430\,
            I => \N__35427\
        );

    \I__8812\ : Span4Mux_h
    port map (
            O => \N__35427\,
            I => \N__35424\
        );

    \I__8811\ : Sp12to4
    port map (
            O => \N__35424\,
            I => \N__35420\
        );

    \I__8810\ : InMux
    port map (
            O => \N__35423\,
            I => \N__35417\
        );

    \I__8809\ : Odrv12
    port map (
            O => \N__35420\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__35417\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__8807\ : InMux
    port map (
            O => \N__35412\,
            I => \M_this_external_address_q_cry_1\
        );

    \I__8806\ : IoInMux
    port map (
            O => \N__35409\,
            I => \N__35406\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__35406\,
            I => \N__35403\
        );

    \I__8804\ : Span4Mux_s2_h
    port map (
            O => \N__35403\,
            I => \N__35400\
        );

    \I__8803\ : Span4Mux_h
    port map (
            O => \N__35400\,
            I => \N__35397\
        );

    \I__8802\ : Span4Mux_v
    port map (
            O => \N__35397\,
            I => \N__35393\
        );

    \I__8801\ : InMux
    port map (
            O => \N__35396\,
            I => \N__35390\
        );

    \I__8800\ : Odrv4
    port map (
            O => \N__35393\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__8799\ : LocalMux
    port map (
            O => \N__35390\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__8798\ : InMux
    port map (
            O => \N__35385\,
            I => \M_this_external_address_q_cry_2\
        );

    \I__8797\ : IoInMux
    port map (
            O => \N__35382\,
            I => \N__35379\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__35379\,
            I => \N__35376\
        );

    \I__8795\ : Span4Mux_s2_h
    port map (
            O => \N__35376\,
            I => \N__35373\
        );

    \I__8794\ : Span4Mux_h
    port map (
            O => \N__35373\,
            I => \N__35369\
        );

    \I__8793\ : InMux
    port map (
            O => \N__35372\,
            I => \N__35366\
        );

    \I__8792\ : Odrv4
    port map (
            O => \N__35369\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__35366\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__8790\ : InMux
    port map (
            O => \N__35361\,
            I => \N__35358\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__35358\,
            I => \N__35355\
        );

    \I__8788\ : Odrv4
    port map (
            O => \N__35355\,
            I => \this_vga_signals.N_665_1\
        );

    \I__8787\ : InMux
    port map (
            O => \N__35352\,
            I => \N__35349\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__35349\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_3LZ0Z4\
        );

    \I__8785\ : InMux
    port map (
            O => \N__35346\,
            I => \N__35343\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__35343\,
            I => \N__35340\
        );

    \I__8783\ : Odrv12
    port map (
            O => \N__35340\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_4LZ0Z6\
        );

    \I__8782\ : InMux
    port map (
            O => \N__35337\,
            I => \N__35334\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__35334\,
            I => \N__35331\
        );

    \I__8780\ : Span4Mux_v
    port map (
            O => \N__35331\,
            I => \N__35328\
        );

    \I__8779\ : Span4Mux_h
    port map (
            O => \N__35328\,
            I => \N__35324\
        );

    \I__8778\ : InMux
    port map (
            O => \N__35327\,
            I => \N__35321\
        );

    \I__8777\ : Span4Mux_v
    port map (
            O => \N__35324\,
            I => \N__35318\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__35321\,
            I => \N__35315\
        );

    \I__8775\ : Sp12to4
    port map (
            O => \N__35318\,
            I => \N__35310\
        );

    \I__8774\ : Span12Mux_v
    port map (
            O => \N__35315\,
            I => \N__35310\
        );

    \I__8773\ : Odrv12
    port map (
            O => \N__35310\,
            I => port_address_in_3
        );

    \I__8772\ : CascadeMux
    port map (
            O => \N__35307\,
            I => \N__35303\
        );

    \I__8771\ : InMux
    port map (
            O => \N__35306\,
            I => \N__35300\
        );

    \I__8770\ : InMux
    port map (
            O => \N__35303\,
            I => \N__35297\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__35300\,
            I => \N__35292\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__35297\,
            I => \N__35292\
        );

    \I__8767\ : Odrv12
    port map (
            O => \N__35292\,
            I => port_address_in_5
        );

    \I__8766\ : CascadeMux
    port map (
            O => \N__35289\,
            I => \N__35286\
        );

    \I__8765\ : InMux
    port map (
            O => \N__35286\,
            I => \N__35280\
        );

    \I__8764\ : InMux
    port map (
            O => \N__35285\,
            I => \N__35280\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__35280\,
            I => \N__35277\
        );

    \I__8762\ : Span12Mux_v
    port map (
            O => \N__35277\,
            I => \N__35274\
        );

    \I__8761\ : Odrv12
    port map (
            O => \N__35274\,
            I => port_address_in_6
        );

    \I__8760\ : InMux
    port map (
            O => \N__35271\,
            I => \N__35265\
        );

    \I__8759\ : InMux
    port map (
            O => \N__35270\,
            I => \N__35265\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__35265\,
            I => \N__35262\
        );

    \I__8757\ : Span4Mux_v
    port map (
            O => \N__35262\,
            I => \N__35259\
        );

    \I__8756\ : Span4Mux_h
    port map (
            O => \N__35259\,
            I => \N__35256\
        );

    \I__8755\ : Odrv4
    port map (
            O => \N__35256\,
            I => port_address_in_4
        );

    \I__8754\ : InMux
    port map (
            O => \N__35253\,
            I => \N__35250\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__35250\,
            I => \N__35247\
        );

    \I__8752\ : Span4Mux_h
    port map (
            O => \N__35247\,
            I => \N__35244\
        );

    \I__8751\ : Span4Mux_h
    port map (
            O => \N__35244\,
            I => \N__35241\
        );

    \I__8750\ : Odrv4
    port map (
            O => \N__35241\,
            I => \this_vga_signals.un1_M_this_state_q_19_i_0_o2Z0Z_4\
        );

    \I__8749\ : CascadeMux
    port map (
            O => \N__35238\,
            I => \N__35235\
        );

    \I__8748\ : InMux
    port map (
            O => \N__35235\,
            I => \N__35230\
        );

    \I__8747\ : InMux
    port map (
            O => \N__35234\,
            I => \N__35225\
        );

    \I__8746\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35221\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__35230\,
            I => \N__35215\
        );

    \I__8744\ : InMux
    port map (
            O => \N__35229\,
            I => \N__35212\
        );

    \I__8743\ : CascadeMux
    port map (
            O => \N__35228\,
            I => \N__35208\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__35225\,
            I => \N__35204\
        );

    \I__8741\ : CascadeMux
    port map (
            O => \N__35224\,
            I => \N__35200\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__35221\,
            I => \N__35197\
        );

    \I__8739\ : InMux
    port map (
            O => \N__35220\,
            I => \N__35194\
        );

    \I__8738\ : InMux
    port map (
            O => \N__35219\,
            I => \N__35189\
        );

    \I__8737\ : InMux
    port map (
            O => \N__35218\,
            I => \N__35189\
        );

    \I__8736\ : Span4Mux_v
    port map (
            O => \N__35215\,
            I => \N__35184\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__35212\,
            I => \N__35184\
        );

    \I__8734\ : InMux
    port map (
            O => \N__35211\,
            I => \N__35179\
        );

    \I__8733\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35179\
        );

    \I__8732\ : CascadeMux
    port map (
            O => \N__35207\,
            I => \N__35176\
        );

    \I__8731\ : Span4Mux_v
    port map (
            O => \N__35204\,
            I => \N__35173\
        );

    \I__8730\ : InMux
    port map (
            O => \N__35203\,
            I => \N__35169\
        );

    \I__8729\ : InMux
    port map (
            O => \N__35200\,
            I => \N__35165\
        );

    \I__8728\ : Span4Mux_v
    port map (
            O => \N__35197\,
            I => \N__35153\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__35194\,
            I => \N__35153\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__35189\,
            I => \N__35153\
        );

    \I__8725\ : Span4Mux_h
    port map (
            O => \N__35184\,
            I => \N__35153\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__35179\,
            I => \N__35153\
        );

    \I__8723\ : InMux
    port map (
            O => \N__35176\,
            I => \N__35150\
        );

    \I__8722\ : Span4Mux_v
    port map (
            O => \N__35173\,
            I => \N__35147\
        );

    \I__8721\ : CascadeMux
    port map (
            O => \N__35172\,
            I => \N__35144\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__35169\,
            I => \N__35141\
        );

    \I__8719\ : InMux
    port map (
            O => \N__35168\,
            I => \N__35138\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__35165\,
            I => \N__35133\
        );

    \I__8717\ : InMux
    port map (
            O => \N__35164\,
            I => \N__35130\
        );

    \I__8716\ : Span4Mux_v
    port map (
            O => \N__35153\,
            I => \N__35125\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__35150\,
            I => \N__35125\
        );

    \I__8714\ : Span4Mux_v
    port map (
            O => \N__35147\,
            I => \N__35122\
        );

    \I__8713\ : InMux
    port map (
            O => \N__35144\,
            I => \N__35119\
        );

    \I__8712\ : Span4Mux_v
    port map (
            O => \N__35141\,
            I => \N__35114\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__35138\,
            I => \N__35114\
        );

    \I__8710\ : InMux
    port map (
            O => \N__35137\,
            I => \N__35111\
        );

    \I__8709\ : InMux
    port map (
            O => \N__35136\,
            I => \N__35108\
        );

    \I__8708\ : Span4Mux_v
    port map (
            O => \N__35133\,
            I => \N__35105\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__35130\,
            I => \N__35102\
        );

    \I__8706\ : Span4Mux_v
    port map (
            O => \N__35125\,
            I => \N__35099\
        );

    \I__8705\ : Span4Mux_v
    port map (
            O => \N__35122\,
            I => \N__35094\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__35119\,
            I => \N__35094\
        );

    \I__8703\ : Span4Mux_h
    port map (
            O => \N__35114\,
            I => \N__35091\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__35111\,
            I => \N__35088\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__35108\,
            I => \N__35085\
        );

    \I__8700\ : Span4Mux_h
    port map (
            O => \N__35105\,
            I => \N__35080\
        );

    \I__8699\ : Span4Mux_v
    port map (
            O => \N__35102\,
            I => \N__35080\
        );

    \I__8698\ : Span4Mux_h
    port map (
            O => \N__35099\,
            I => \N__35075\
        );

    \I__8697\ : Span4Mux_v
    port map (
            O => \N__35094\,
            I => \N__35075\
        );

    \I__8696\ : Sp12to4
    port map (
            O => \N__35091\,
            I => \N__35072\
        );

    \I__8695\ : Span12Mux_s7_v
    port map (
            O => \N__35088\,
            I => \N__35069\
        );

    \I__8694\ : Span12Mux_h
    port map (
            O => \N__35085\,
            I => \N__35066\
        );

    \I__8693\ : Span4Mux_h
    port map (
            O => \N__35080\,
            I => \N__35063\
        );

    \I__8692\ : Span4Mux_v
    port map (
            O => \N__35075\,
            I => \N__35060\
        );

    \I__8691\ : Span12Mux_v
    port map (
            O => \N__35072\,
            I => \N__35055\
        );

    \I__8690\ : Span12Mux_h
    port map (
            O => \N__35069\,
            I => \N__35055\
        );

    \I__8689\ : Span12Mux_v
    port map (
            O => \N__35066\,
            I => \N__35050\
        );

    \I__8688\ : Sp12to4
    port map (
            O => \N__35063\,
            I => \N__35050\
        );

    \I__8687\ : IoSpan4Mux
    port map (
            O => \N__35060\,
            I => \N__35047\
        );

    \I__8686\ : Odrv12
    port map (
            O => \N__35055\,
            I => port_data_c_2
        );

    \I__8685\ : Odrv12
    port map (
            O => \N__35050\,
            I => port_data_c_2
        );

    \I__8684\ : Odrv4
    port map (
            O => \N__35047\,
            I => port_data_c_2
        );

    \I__8683\ : InMux
    port map (
            O => \N__35040\,
            I => \N__35032\
        );

    \I__8682\ : InMux
    port map (
            O => \N__35039\,
            I => \N__35029\
        );

    \I__8681\ : InMux
    port map (
            O => \N__35038\,
            I => \N__35026\
        );

    \I__8680\ : InMux
    port map (
            O => \N__35037\,
            I => \N__35023\
        );

    \I__8679\ : InMux
    port map (
            O => \N__35036\,
            I => \N__35020\
        );

    \I__8678\ : InMux
    port map (
            O => \N__35035\,
            I => \N__35017\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__35032\,
            I => \N__35014\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__35029\,
            I => \N__35007\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__35026\,
            I => \N__35007\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__35023\,
            I => \N__35007\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__35020\,
            I => \N_760\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__35017\,
            I => \N_760\
        );

    \I__8671\ : Odrv4
    port map (
            O => \N__35014\,
            I => \N_760\
        );

    \I__8670\ : Odrv4
    port map (
            O => \N__35007\,
            I => \N_760\
        );

    \I__8669\ : InMux
    port map (
            O => \N__34998\,
            I => \N__34988\
        );

    \I__8668\ : InMux
    port map (
            O => \N__34997\,
            I => \N__34983\
        );

    \I__8667\ : InMux
    port map (
            O => \N__34996\,
            I => \N__34983\
        );

    \I__8666\ : InMux
    port map (
            O => \N__34995\,
            I => \N__34980\
        );

    \I__8665\ : InMux
    port map (
            O => \N__34994\,
            I => \N__34977\
        );

    \I__8664\ : InMux
    port map (
            O => \N__34993\,
            I => \N__34974\
        );

    \I__8663\ : InMux
    port map (
            O => \N__34992\,
            I => \N__34971\
        );

    \I__8662\ : InMux
    port map (
            O => \N__34991\,
            I => \N__34968\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__34988\,
            I => \N__34963\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__34983\,
            I => \N__34963\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__34980\,
            I => \N__34960\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__34977\,
            I => \N__34957\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__34974\,
            I => \N__34948\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__34971\,
            I => \N__34948\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__34968\,
            I => \N__34943\
        );

    \I__8654\ : Span4Mux_v
    port map (
            O => \N__34963\,
            I => \N__34943\
        );

    \I__8653\ : Span4Mux_v
    port map (
            O => \N__34960\,
            I => \N__34938\
        );

    \I__8652\ : Span4Mux_v
    port map (
            O => \N__34957\,
            I => \N__34938\
        );

    \I__8651\ : InMux
    port map (
            O => \N__34956\,
            I => \N__34931\
        );

    \I__8650\ : InMux
    port map (
            O => \N__34955\,
            I => \N__34931\
        );

    \I__8649\ : InMux
    port map (
            O => \N__34954\,
            I => \N__34931\
        );

    \I__8648\ : InMux
    port map (
            O => \N__34953\,
            I => \N__34928\
        );

    \I__8647\ : Span4Mux_v
    port map (
            O => \N__34948\,
            I => \N__34921\
        );

    \I__8646\ : Span4Mux_v
    port map (
            O => \N__34943\,
            I => \N__34921\
        );

    \I__8645\ : Span4Mux_h
    port map (
            O => \N__34938\,
            I => \N__34921\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__34931\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__34928\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__8642\ : Odrv4
    port map (
            O => \N__34921\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__8641\ : InMux
    port map (
            O => \N__34914\,
            I => \N__34907\
        );

    \I__8640\ : CascadeMux
    port map (
            O => \N__34913\,
            I => \N__34902\
        );

    \I__8639\ : InMux
    port map (
            O => \N__34912\,
            I => \N__34899\
        );

    \I__8638\ : InMux
    port map (
            O => \N__34911\,
            I => \N__34896\
        );

    \I__8637\ : InMux
    port map (
            O => \N__34910\,
            I => \N__34893\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__34907\,
            I => \N__34890\
        );

    \I__8635\ : InMux
    port map (
            O => \N__34906\,
            I => \N__34886\
        );

    \I__8634\ : InMux
    port map (
            O => \N__34905\,
            I => \N__34881\
        );

    \I__8633\ : InMux
    port map (
            O => \N__34902\,
            I => \N__34881\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__34899\,
            I => \N__34878\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__34896\,
            I => \N__34873\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__34893\,
            I => \N__34873\
        );

    \I__8629\ : Span4Mux_h
    port map (
            O => \N__34890\,
            I => \N__34870\
        );

    \I__8628\ : InMux
    port map (
            O => \N__34889\,
            I => \N__34867\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__34886\,
            I => \N__34864\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__34881\,
            I => \N__34861\
        );

    \I__8625\ : Span4Mux_h
    port map (
            O => \N__34878\,
            I => \N__34858\
        );

    \I__8624\ : Span4Mux_h
    port map (
            O => \N__34873\,
            I => \N__34853\
        );

    \I__8623\ : Span4Mux_h
    port map (
            O => \N__34870\,
            I => \N__34853\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__34867\,
            I => \N__34850\
        );

    \I__8621\ : Span4Mux_h
    port map (
            O => \N__34864\,
            I => \N__34847\
        );

    \I__8620\ : Span4Mux_h
    port map (
            O => \N__34861\,
            I => \N__34840\
        );

    \I__8619\ : Span4Mux_h
    port map (
            O => \N__34858\,
            I => \N__34840\
        );

    \I__8618\ : Span4Mux_v
    port map (
            O => \N__34853\,
            I => \N__34840\
        );

    \I__8617\ : Odrv12
    port map (
            O => \N__34850\,
            I => \N_25_0\
        );

    \I__8616\ : Odrv4
    port map (
            O => \N__34847\,
            I => \N_25_0\
        );

    \I__8615\ : Odrv4
    port map (
            O => \N__34840\,
            I => \N_25_0\
        );

    \I__8614\ : CascadeMux
    port map (
            O => \N__34833\,
            I => \N__34825\
        );

    \I__8613\ : CascadeMux
    port map (
            O => \N__34832\,
            I => \N__34822\
        );

    \I__8612\ : InMux
    port map (
            O => \N__34831\,
            I => \N__34815\
        );

    \I__8611\ : CascadeMux
    port map (
            O => \N__34830\,
            I => \N__34812\
        );

    \I__8610\ : CascadeMux
    port map (
            O => \N__34829\,
            I => \N__34809\
        );

    \I__8609\ : CascadeMux
    port map (
            O => \N__34828\,
            I => \N__34806\
        );

    \I__8608\ : InMux
    port map (
            O => \N__34825\,
            I => \N__34803\
        );

    \I__8607\ : InMux
    port map (
            O => \N__34822\,
            I => \N__34798\
        );

    \I__8606\ : InMux
    port map (
            O => \N__34821\,
            I => \N__34798\
        );

    \I__8605\ : CascadeMux
    port map (
            O => \N__34820\,
            I => \N__34795\
        );

    \I__8604\ : CascadeMux
    port map (
            O => \N__34819\,
            I => \N__34792\
        );

    \I__8603\ : InMux
    port map (
            O => \N__34818\,
            I => \N__34789\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__34815\,
            I => \N__34786\
        );

    \I__8601\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34783\
        );

    \I__8600\ : InMux
    port map (
            O => \N__34809\,
            I => \N__34780\
        );

    \I__8599\ : InMux
    port map (
            O => \N__34806\,
            I => \N__34777\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__34803\,
            I => \N__34772\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__34798\,
            I => \N__34772\
        );

    \I__8596\ : InMux
    port map (
            O => \N__34795\,
            I => \N__34768\
        );

    \I__8595\ : InMux
    port map (
            O => \N__34792\,
            I => \N__34765\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__34789\,
            I => \N__34762\
        );

    \I__8593\ : Span4Mux_v
    port map (
            O => \N__34786\,
            I => \N__34759\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__34783\,
            I => \N__34754\
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__34780\,
            I => \N__34754\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__34777\,
            I => \N__34749\
        );

    \I__8589\ : Span4Mux_v
    port map (
            O => \N__34772\,
            I => \N__34749\
        );

    \I__8588\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34745\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__34768\,
            I => \N__34742\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__34765\,
            I => \N__34739\
        );

    \I__8585\ : Span4Mux_v
    port map (
            O => \N__34762\,
            I => \N__34730\
        );

    \I__8584\ : Span4Mux_h
    port map (
            O => \N__34759\,
            I => \N__34730\
        );

    \I__8583\ : Span4Mux_v
    port map (
            O => \N__34754\,
            I => \N__34730\
        );

    \I__8582\ : Span4Mux_v
    port map (
            O => \N__34749\,
            I => \N__34730\
        );

    \I__8581\ : InMux
    port map (
            O => \N__34748\,
            I => \N__34727\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__34745\,
            I => \N__34724\
        );

    \I__8579\ : Span4Mux_v
    port map (
            O => \N__34742\,
            I => \N__34717\
        );

    \I__8578\ : Span4Mux_v
    port map (
            O => \N__34739\,
            I => \N__34717\
        );

    \I__8577\ : Span4Mux_h
    port map (
            O => \N__34730\,
            I => \N__34717\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__34727\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__8575\ : Odrv4
    port map (
            O => \N__34724\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__8574\ : Odrv4
    port map (
            O => \N__34717\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__8573\ : InMux
    port map (
            O => \N__34710\,
            I => \N__34703\
        );

    \I__8572\ : InMux
    port map (
            O => \N__34709\,
            I => \N__34703\
        );

    \I__8571\ : InMux
    port map (
            O => \N__34708\,
            I => \N__34700\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__34703\,
            I => \N__34694\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__34700\,
            I => \N__34694\
        );

    \I__8568\ : InMux
    port map (
            O => \N__34699\,
            I => \N__34690\
        );

    \I__8567\ : Span4Mux_v
    port map (
            O => \N__34694\,
            I => \N__34687\
        );

    \I__8566\ : InMux
    port map (
            O => \N__34693\,
            I => \N__34684\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__34690\,
            I => \N__34679\
        );

    \I__8564\ : Sp12to4
    port map (
            O => \N__34687\,
            I => \N__34670\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__34684\,
            I => \N__34670\
        );

    \I__8562\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34667\
        );

    \I__8561\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34664\
        );

    \I__8560\ : Span4Mux_h
    port map (
            O => \N__34679\,
            I => \N__34661\
        );

    \I__8559\ : InMux
    port map (
            O => \N__34678\,
            I => \N__34658\
        );

    \I__8558\ : CascadeMux
    port map (
            O => \N__34677\,
            I => \N__34655\
        );

    \I__8557\ : CascadeMux
    port map (
            O => \N__34676\,
            I => \N__34652\
        );

    \I__8556\ : InMux
    port map (
            O => \N__34675\,
            I => \N__34648\
        );

    \I__8555\ : Span12Mux_h
    port map (
            O => \N__34670\,
            I => \N__34645\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__34667\,
            I => \N__34640\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__34664\,
            I => \N__34640\
        );

    \I__8552\ : Span4Mux_v
    port map (
            O => \N__34661\,
            I => \N__34635\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__34658\,
            I => \N__34635\
        );

    \I__8550\ : InMux
    port map (
            O => \N__34655\,
            I => \N__34632\
        );

    \I__8549\ : InMux
    port map (
            O => \N__34652\,
            I => \N__34629\
        );

    \I__8548\ : InMux
    port map (
            O => \N__34651\,
            I => \N__34626\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__34648\,
            I => \N__34623\
        );

    \I__8546\ : Odrv12
    port map (
            O => \N__34645\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__8545\ : Odrv12
    port map (
            O => \N__34640\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__8544\ : Odrv4
    port map (
            O => \N__34635\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__34632\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__34629\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__34626\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__8540\ : Odrv4
    port map (
            O => \N__34623\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__8539\ : CEMux
    port map (
            O => \N__34608\,
            I => \N__34604\
        );

    \I__8538\ : CEMux
    port map (
            O => \N__34607\,
            I => \N__34601\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__34604\,
            I => \N__34596\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__34601\,
            I => \N__34596\
        );

    \I__8535\ : Span4Mux_v
    port map (
            O => \N__34596\,
            I => \N__34593\
        );

    \I__8534\ : Odrv4
    port map (
            O => \N__34593\,
            I => \this_sprites_ram.mem_WE_6\
        );

    \I__8533\ : InMux
    port map (
            O => \N__34590\,
            I => \N__34587\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__34587\,
            I => \N__34584\
        );

    \I__8531\ : Odrv4
    port map (
            O => \N__34584\,
            I => \M_this_oam_ram_write_data_14\
        );

    \I__8530\ : InMux
    port map (
            O => \N__34581\,
            I => \N__34578\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__34578\,
            I => \N__34574\
        );

    \I__8528\ : CascadeMux
    port map (
            O => \N__34577\,
            I => \N__34570\
        );

    \I__8527\ : Span4Mux_v
    port map (
            O => \N__34574\,
            I => \N__34566\
        );

    \I__8526\ : InMux
    port map (
            O => \N__34573\,
            I => \N__34561\
        );

    \I__8525\ : InMux
    port map (
            O => \N__34570\,
            I => \N__34561\
        );

    \I__8524\ : CascadeMux
    port map (
            O => \N__34569\,
            I => \N__34558\
        );

    \I__8523\ : Span4Mux_h
    port map (
            O => \N__34566\,
            I => \N__34553\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__34561\,
            I => \N__34553\
        );

    \I__8521\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34549\
        );

    \I__8520\ : Span4Mux_h
    port map (
            O => \N__34553\,
            I => \N__34546\
        );

    \I__8519\ : InMux
    port map (
            O => \N__34552\,
            I => \N__34543\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__34549\,
            I => \N__34539\
        );

    \I__8517\ : Span4Mux_h
    port map (
            O => \N__34546\,
            I => \N__34536\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__34543\,
            I => \N__34533\
        );

    \I__8515\ : InMux
    port map (
            O => \N__34542\,
            I => \N__34530\
        );

    \I__8514\ : Span4Mux_v
    port map (
            O => \N__34539\,
            I => \N__34526\
        );

    \I__8513\ : Span4Mux_v
    port map (
            O => \N__34536\,
            I => \N__34521\
        );

    \I__8512\ : Span4Mux_h
    port map (
            O => \N__34533\,
            I => \N__34521\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__34530\,
            I => \N__34518\
        );

    \I__8510\ : InMux
    port map (
            O => \N__34529\,
            I => \N__34515\
        );

    \I__8509\ : Span4Mux_h
    port map (
            O => \N__34526\,
            I => \N__34510\
        );

    \I__8508\ : Span4Mux_v
    port map (
            O => \N__34521\,
            I => \N__34507\
        );

    \I__8507\ : Span4Mux_v
    port map (
            O => \N__34518\,
            I => \N__34504\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__34515\,
            I => \N__34501\
        );

    \I__8505\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34498\
        );

    \I__8504\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34495\
        );

    \I__8503\ : Sp12to4
    port map (
            O => \N__34510\,
            I => \N__34490\
        );

    \I__8502\ : Sp12to4
    port map (
            O => \N__34507\,
            I => \N__34490\
        );

    \I__8501\ : Span4Mux_h
    port map (
            O => \N__34504\,
            I => \N__34485\
        );

    \I__8500\ : Span4Mux_v
    port map (
            O => \N__34501\,
            I => \N__34485\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__34498\,
            I => \N__34482\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__34495\,
            I => \N__34479\
        );

    \I__8497\ : Span12Mux_v
    port map (
            O => \N__34490\,
            I => \N__34470\
        );

    \I__8496\ : Sp12to4
    port map (
            O => \N__34485\,
            I => \N__34470\
        );

    \I__8495\ : Span12Mux_h
    port map (
            O => \N__34482\,
            I => \N__34470\
        );

    \I__8494\ : Span12Mux_s9_v
    port map (
            O => \N__34479\,
            I => \N__34470\
        );

    \I__8493\ : Odrv12
    port map (
            O => \N__34470\,
            I => port_data_c_7
        );

    \I__8492\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34464\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__34464\,
            I => \N__34461\
        );

    \I__8490\ : Span4Mux_h
    port map (
            O => \N__34461\,
            I => \N__34458\
        );

    \I__8489\ : Odrv4
    port map (
            O => \N__34458\,
            I => \M_this_data_tmp_qZ0Z_15\
        );

    \I__8488\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34452\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__34452\,
            I => \N__34449\
        );

    \I__8486\ : Span4Mux_h
    port map (
            O => \N__34449\,
            I => \N__34446\
        );

    \I__8485\ : Span4Mux_h
    port map (
            O => \N__34446\,
            I => \N__34436\
        );

    \I__8484\ : InMux
    port map (
            O => \N__34445\,
            I => \N__34433\
        );

    \I__8483\ : InMux
    port map (
            O => \N__34444\,
            I => \N__34428\
        );

    \I__8482\ : InMux
    port map (
            O => \N__34443\,
            I => \N__34428\
        );

    \I__8481\ : CascadeMux
    port map (
            O => \N__34442\,
            I => \N__34425\
        );

    \I__8480\ : InMux
    port map (
            O => \N__34441\,
            I => \N__34421\
        );

    \I__8479\ : InMux
    port map (
            O => \N__34440\,
            I => \N__34418\
        );

    \I__8478\ : CascadeMux
    port map (
            O => \N__34439\,
            I => \N__34414\
        );

    \I__8477\ : Span4Mux_v
    port map (
            O => \N__34436\,
            I => \N__34407\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__34433\,
            I => \N__34407\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__34428\,
            I => \N__34407\
        );

    \I__8474\ : InMux
    port map (
            O => \N__34425\,
            I => \N__34404\
        );

    \I__8473\ : CascadeMux
    port map (
            O => \N__34424\,
            I => \N__34401\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__34421\,
            I => \N__34398\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__34418\,
            I => \N__34395\
        );

    \I__8470\ : InMux
    port map (
            O => \N__34417\,
            I => \N__34392\
        );

    \I__8469\ : InMux
    port map (
            O => \N__34414\,
            I => \N__34388\
        );

    \I__8468\ : Span4Mux_v
    port map (
            O => \N__34407\,
            I => \N__34385\
        );

    \I__8467\ : LocalMux
    port map (
            O => \N__34404\,
            I => \N__34382\
        );

    \I__8466\ : InMux
    port map (
            O => \N__34401\,
            I => \N__34379\
        );

    \I__8465\ : Span4Mux_v
    port map (
            O => \N__34398\,
            I => \N__34372\
        );

    \I__8464\ : Span4Mux_v
    port map (
            O => \N__34395\,
            I => \N__34372\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__34392\,
            I => \N__34372\
        );

    \I__8462\ : InMux
    port map (
            O => \N__34391\,
            I => \N__34369\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__34388\,
            I => \N__34366\
        );

    \I__8460\ : Span4Mux_h
    port map (
            O => \N__34385\,
            I => \N__34359\
        );

    \I__8459\ : Span4Mux_h
    port map (
            O => \N__34382\,
            I => \N__34359\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__34379\,
            I => \N__34359\
        );

    \I__8457\ : Span4Mux_h
    port map (
            O => \N__34372\,
            I => \N__34354\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__34369\,
            I => \N__34354\
        );

    \I__8455\ : Span12Mux_h
    port map (
            O => \N__34366\,
            I => \N__34351\
        );

    \I__8454\ : Sp12to4
    port map (
            O => \N__34359\,
            I => \N__34348\
        );

    \I__8453\ : Span4Mux_h
    port map (
            O => \N__34354\,
            I => \N__34345\
        );

    \I__8452\ : Span12Mux_v
    port map (
            O => \N__34351\,
            I => \N__34342\
        );

    \I__8451\ : Span12Mux_v
    port map (
            O => \N__34348\,
            I => \N__34339\
        );

    \I__8450\ : Span4Mux_v
    port map (
            O => \N__34345\,
            I => \N__34336\
        );

    \I__8449\ : Odrv12
    port map (
            O => \N__34342\,
            I => port_data_c_6
        );

    \I__8448\ : Odrv12
    port map (
            O => \N__34339\,
            I => port_data_c_6
        );

    \I__8447\ : Odrv4
    port map (
            O => \N__34336\,
            I => port_data_c_6
        );

    \I__8446\ : InMux
    port map (
            O => \N__34329\,
            I => \N__34326\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__34326\,
            I => \N__34323\
        );

    \I__8444\ : Odrv4
    port map (
            O => \N__34323\,
            I => \M_this_data_tmp_qZ0Z_14\
        );

    \I__8443\ : InMux
    port map (
            O => \N__34320\,
            I => \N__34317\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__34317\,
            I => \this_ppu.un2_hscroll_axb_0\
        );

    \I__8441\ : CascadeMux
    port map (
            O => \N__34314\,
            I => \N__34311\
        );

    \I__8440\ : InMux
    port map (
            O => \N__34311\,
            I => \N__34308\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__34308\,
            I => \N__34304\
        );

    \I__8438\ : CascadeMux
    port map (
            O => \N__34307\,
            I => \N__34298\
        );

    \I__8437\ : Span4Mux_v
    port map (
            O => \N__34304\,
            I => \N__34294\
        );

    \I__8436\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34291\
        );

    \I__8435\ : InMux
    port map (
            O => \N__34302\,
            I => \N__34287\
        );

    \I__8434\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34284\
        );

    \I__8433\ : InMux
    port map (
            O => \N__34298\,
            I => \N__34280\
        );

    \I__8432\ : InMux
    port map (
            O => \N__34297\,
            I => \N__34277\
        );

    \I__8431\ : Sp12to4
    port map (
            O => \N__34294\,
            I => \N__34274\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__34291\,
            I => \N__34271\
        );

    \I__8429\ : InMux
    port map (
            O => \N__34290\,
            I => \N__34268\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__34287\,
            I => \N__34264\
        );

    \I__8427\ : LocalMux
    port map (
            O => \N__34284\,
            I => \N__34261\
        );

    \I__8426\ : InMux
    port map (
            O => \N__34283\,
            I => \N__34258\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__34280\,
            I => \N__34255\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__34277\,
            I => \N__34252\
        );

    \I__8423\ : Span12Mux_h
    port map (
            O => \N__34274\,
            I => \N__34249\
        );

    \I__8422\ : Span4Mux_v
    port map (
            O => \N__34271\,
            I => \N__34244\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__34268\,
            I => \N__34244\
        );

    \I__8420\ : InMux
    port map (
            O => \N__34267\,
            I => \N__34241\
        );

    \I__8419\ : Sp12to4
    port map (
            O => \N__34264\,
            I => \N__34236\
        );

    \I__8418\ : Span12Mux_v
    port map (
            O => \N__34261\,
            I => \N__34236\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__34258\,
            I => \N__34231\
        );

    \I__8416\ : Span12Mux_h
    port map (
            O => \N__34255\,
            I => \N__34231\
        );

    \I__8415\ : Span4Mux_v
    port map (
            O => \N__34252\,
            I => \N__34228\
        );

    \I__8414\ : Odrv12
    port map (
            O => \N__34249\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__8413\ : Odrv4
    port map (
            O => \N__34244\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__34241\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__8411\ : Odrv12
    port map (
            O => \N__34236\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__8410\ : Odrv12
    port map (
            O => \N__34231\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__8409\ : Odrv4
    port map (
            O => \N__34228\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__8408\ : CascadeMux
    port map (
            O => \N__34215\,
            I => \N__34210\
        );

    \I__8407\ : CascadeMux
    port map (
            O => \N__34214\,
            I => \N__34207\
        );

    \I__8406\ : CascadeMux
    port map (
            O => \N__34213\,
            I => \N__34204\
        );

    \I__8405\ : InMux
    port map (
            O => \N__34210\,
            I => \N__34200\
        );

    \I__8404\ : InMux
    port map (
            O => \N__34207\,
            I => \N__34197\
        );

    \I__8403\ : InMux
    port map (
            O => \N__34204\,
            I => \N__34194\
        );

    \I__8402\ : CascadeMux
    port map (
            O => \N__34203\,
            I => \N__34191\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__34200\,
            I => \N__34185\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__34197\,
            I => \N__34185\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__34194\,
            I => \N__34182\
        );

    \I__8398\ : InMux
    port map (
            O => \N__34191\,
            I => \N__34179\
        );

    \I__8397\ : CascadeMux
    port map (
            O => \N__34190\,
            I => \N__34176\
        );

    \I__8396\ : Span4Mux_v
    port map (
            O => \N__34185\,
            I => \N__34167\
        );

    \I__8395\ : Span4Mux_h
    port map (
            O => \N__34182\,
            I => \N__34167\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__34179\,
            I => \N__34167\
        );

    \I__8393\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34164\
        );

    \I__8392\ : CascadeMux
    port map (
            O => \N__34175\,
            I => \N__34161\
        );

    \I__8391\ : CascadeMux
    port map (
            O => \N__34174\,
            I => \N__34158\
        );

    \I__8390\ : Span4Mux_v
    port map (
            O => \N__34167\,
            I => \N__34153\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__34164\,
            I => \N__34150\
        );

    \I__8388\ : InMux
    port map (
            O => \N__34161\,
            I => \N__34147\
        );

    \I__8387\ : InMux
    port map (
            O => \N__34158\,
            I => \N__34144\
        );

    \I__8386\ : CascadeMux
    port map (
            O => \N__34157\,
            I => \N__34141\
        );

    \I__8385\ : CascadeMux
    port map (
            O => \N__34156\,
            I => \N__34138\
        );

    \I__8384\ : Span4Mux_h
    port map (
            O => \N__34153\,
            I => \N__34132\
        );

    \I__8383\ : Span4Mux_s3_v
    port map (
            O => \N__34150\,
            I => \N__34125\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__34147\,
            I => \N__34125\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__34144\,
            I => \N__34125\
        );

    \I__8380\ : InMux
    port map (
            O => \N__34141\,
            I => \N__34122\
        );

    \I__8379\ : InMux
    port map (
            O => \N__34138\,
            I => \N__34119\
        );

    \I__8378\ : CascadeMux
    port map (
            O => \N__34137\,
            I => \N__34116\
        );

    \I__8377\ : CascadeMux
    port map (
            O => \N__34136\,
            I => \N__34113\
        );

    \I__8376\ : CascadeMux
    port map (
            O => \N__34135\,
            I => \N__34108\
        );

    \I__8375\ : Span4Mux_h
    port map (
            O => \N__34132\,
            I => \N__34105\
        );

    \I__8374\ : Span4Mux_v
    port map (
            O => \N__34125\,
            I => \N__34098\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__34122\,
            I => \N__34098\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__34119\,
            I => \N__34098\
        );

    \I__8371\ : InMux
    port map (
            O => \N__34116\,
            I => \N__34095\
        );

    \I__8370\ : InMux
    port map (
            O => \N__34113\,
            I => \N__34092\
        );

    \I__8369\ : CascadeMux
    port map (
            O => \N__34112\,
            I => \N__34089\
        );

    \I__8368\ : CascadeMux
    port map (
            O => \N__34111\,
            I => \N__34086\
        );

    \I__8367\ : InMux
    port map (
            O => \N__34108\,
            I => \N__34082\
        );

    \I__8366\ : Span4Mux_h
    port map (
            O => \N__34105\,
            I => \N__34079\
        );

    \I__8365\ : Span4Mux_v
    port map (
            O => \N__34098\,
            I => \N__34072\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__34095\,
            I => \N__34072\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__34092\,
            I => \N__34072\
        );

    \I__8362\ : InMux
    port map (
            O => \N__34089\,
            I => \N__34069\
        );

    \I__8361\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34066\
        );

    \I__8360\ : CascadeMux
    port map (
            O => \N__34085\,
            I => \N__34063\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__34082\,
            I => \N__34059\
        );

    \I__8358\ : Span4Mux_h
    port map (
            O => \N__34079\,
            I => \N__34050\
        );

    \I__8357\ : Span4Mux_v
    port map (
            O => \N__34072\,
            I => \N__34050\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__34069\,
            I => \N__34050\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__34066\,
            I => \N__34050\
        );

    \I__8354\ : InMux
    port map (
            O => \N__34063\,
            I => \N__34047\
        );

    \I__8353\ : CascadeMux
    port map (
            O => \N__34062\,
            I => \N__34044\
        );

    \I__8352\ : Span4Mux_h
    port map (
            O => \N__34059\,
            I => \N__34037\
        );

    \I__8351\ : Span4Mux_v
    port map (
            O => \N__34050\,
            I => \N__34037\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__34047\,
            I => \N__34037\
        );

    \I__8349\ : InMux
    port map (
            O => \N__34044\,
            I => \N__34034\
        );

    \I__8348\ : Odrv4
    port map (
            O => \N__34037\,
            I => \M_this_ppu_sprites_addr_0\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__34034\,
            I => \M_this_ppu_sprites_addr_0\
        );

    \I__8346\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34026\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__34026\,
            I => \N__34023\
        );

    \I__8344\ : Odrv12
    port map (
            O => \N__34023\,
            I => \M_this_data_tmp_qZ0Z_19\
        );

    \I__8343\ : CEMux
    port map (
            O => \N__34020\,
            I => \N__34015\
        );

    \I__8342\ : CEMux
    port map (
            O => \N__34019\,
            I => \N__34012\
        );

    \I__8341\ : CEMux
    port map (
            O => \N__34018\,
            I => \N__34009\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__34015\,
            I => \N__34006\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__34012\,
            I => \N__34002\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__34009\,
            I => \N__33999\
        );

    \I__8337\ : Span4Mux_v
    port map (
            O => \N__34006\,
            I => \N__33996\
        );

    \I__8336\ : CEMux
    port map (
            O => \N__34005\,
            I => \N__33993\
        );

    \I__8335\ : Span4Mux_v
    port map (
            O => \N__34002\,
            I => \N__33990\
        );

    \I__8334\ : Span4Mux_v
    port map (
            O => \N__33999\,
            I => \N__33987\
        );

    \I__8333\ : Span4Mux_v
    port map (
            O => \N__33996\,
            I => \N__33982\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__33993\,
            I => \N__33982\
        );

    \I__8331\ : Odrv4
    port map (
            O => \N__33990\,
            I => \N_1396_0\
        );

    \I__8330\ : Odrv4
    port map (
            O => \N__33987\,
            I => \N_1396_0\
        );

    \I__8329\ : Odrv4
    port map (
            O => \N__33982\,
            I => \N_1396_0\
        );

    \I__8328\ : InMux
    port map (
            O => \N__33975\,
            I => \N__33972\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__33972\,
            I => \N__33969\
        );

    \I__8326\ : Span4Mux_v
    port map (
            O => \N__33969\,
            I => \N__33966\
        );

    \I__8325\ : Span4Mux_v
    port map (
            O => \N__33966\,
            I => \N__33963\
        );

    \I__8324\ : Odrv4
    port map (
            O => \N__33963\,
            I => \M_this_oam_ram_read_data_0\
        );

    \I__8323\ : InMux
    port map (
            O => \N__33960\,
            I => \N__33957\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__33957\,
            I => \N__33954\
        );

    \I__8321\ : Span4Mux_v
    port map (
            O => \N__33954\,
            I => \N__33951\
        );

    \I__8320\ : Sp12to4
    port map (
            O => \N__33951\,
            I => \N__33948\
        );

    \I__8319\ : Span12Mux_h
    port map (
            O => \N__33948\,
            I => \N__33945\
        );

    \I__8318\ : Span12Mux_v
    port map (
            O => \N__33945\,
            I => \N__33942\
        );

    \I__8317\ : Odrv12
    port map (
            O => \N__33942\,
            I => \M_this_map_ram_read_data_0\
        );

    \I__8316\ : CascadeMux
    port map (
            O => \N__33939\,
            I => \N__33936\
        );

    \I__8315\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33928\
        );

    \I__8314\ : CascadeMux
    port map (
            O => \N__33935\,
            I => \N__33924\
        );

    \I__8313\ : CascadeMux
    port map (
            O => \N__33934\,
            I => \N__33921\
        );

    \I__8312\ : CascadeMux
    port map (
            O => \N__33933\,
            I => \N__33918\
        );

    \I__8311\ : CascadeMux
    port map (
            O => \N__33932\,
            I => \N__33914\
        );

    \I__8310\ : CascadeMux
    port map (
            O => \N__33931\,
            I => \N__33911\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__33928\,
            I => \N__33908\
        );

    \I__8308\ : CascadeMux
    port map (
            O => \N__33927\,
            I => \N__33903\
        );

    \I__8307\ : InMux
    port map (
            O => \N__33924\,
            I => \N__33898\
        );

    \I__8306\ : InMux
    port map (
            O => \N__33921\,
            I => \N__33898\
        );

    \I__8305\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33894\
        );

    \I__8304\ : InMux
    port map (
            O => \N__33917\,
            I => \N__33889\
        );

    \I__8303\ : InMux
    port map (
            O => \N__33914\,
            I => \N__33889\
        );

    \I__8302\ : InMux
    port map (
            O => \N__33911\,
            I => \N__33885\
        );

    \I__8301\ : Span4Mux_v
    port map (
            O => \N__33908\,
            I => \N__33882\
        );

    \I__8300\ : InMux
    port map (
            O => \N__33907\,
            I => \N__33875\
        );

    \I__8299\ : InMux
    port map (
            O => \N__33906\,
            I => \N__33875\
        );

    \I__8298\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33875\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__33898\,
            I => \N__33872\
        );

    \I__8296\ : CascadeMux
    port map (
            O => \N__33897\,
            I => \N__33869\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__33894\,
            I => \N__33864\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__33889\,
            I => \N__33864\
        );

    \I__8293\ : CascadeMux
    port map (
            O => \N__33888\,
            I => \N__33860\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__33885\,
            I => \N__33857\
        );

    \I__8291\ : Span4Mux_h
    port map (
            O => \N__33882\,
            I => \N__33850\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__33875\,
            I => \N__33850\
        );

    \I__8289\ : Span4Mux_h
    port map (
            O => \N__33872\,
            I => \N__33850\
        );

    \I__8288\ : InMux
    port map (
            O => \N__33869\,
            I => \N__33847\
        );

    \I__8287\ : Span4Mux_v
    port map (
            O => \N__33864\,
            I => \N__33841\
        );

    \I__8286\ : InMux
    port map (
            O => \N__33863\,
            I => \N__33836\
        );

    \I__8285\ : InMux
    port map (
            O => \N__33860\,
            I => \N__33836\
        );

    \I__8284\ : Span4Mux_h
    port map (
            O => \N__33857\,
            I => \N__33829\
        );

    \I__8283\ : Span4Mux_v
    port map (
            O => \N__33850\,
            I => \N__33829\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__33847\,
            I => \N__33829\
        );

    \I__8281\ : CascadeMux
    port map (
            O => \N__33846\,
            I => \N__33826\
        );

    \I__8280\ : CascadeMux
    port map (
            O => \N__33845\,
            I => \N__33823\
        );

    \I__8279\ : InMux
    port map (
            O => \N__33844\,
            I => \N__33820\
        );

    \I__8278\ : Span4Mux_h
    port map (
            O => \N__33841\,
            I => \N__33817\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__33836\,
            I => \N__33814\
        );

    \I__8276\ : Span4Mux_h
    port map (
            O => \N__33829\,
            I => \N__33811\
        );

    \I__8275\ : InMux
    port map (
            O => \N__33826\,
            I => \N__33808\
        );

    \I__8274\ : InMux
    port map (
            O => \N__33823\,
            I => \N__33805\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__33820\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__8272\ : Odrv4
    port map (
            O => \N__33817\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__8271\ : Odrv4
    port map (
            O => \N__33814\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__8270\ : Odrv4
    port map (
            O => \N__33811\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__33808\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__33805\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__8267\ : InMux
    port map (
            O => \N__33792\,
            I => \N__33787\
        );

    \I__8266\ : InMux
    port map (
            O => \N__33791\,
            I => \N__33781\
        );

    \I__8265\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33778\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__33787\,
            I => \N__33768\
        );

    \I__8263\ : InMux
    port map (
            O => \N__33786\,
            I => \N__33761\
        );

    \I__8262\ : InMux
    port map (
            O => \N__33785\,
            I => \N__33761\
        );

    \I__8261\ : InMux
    port map (
            O => \N__33784\,
            I => \N__33761\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__33781\,
            I => \N__33757\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__33778\,
            I => \N__33754\
        );

    \I__8258\ : InMux
    port map (
            O => \N__33777\,
            I => \N__33749\
        );

    \I__8257\ : InMux
    port map (
            O => \N__33776\,
            I => \N__33749\
        );

    \I__8256\ : InMux
    port map (
            O => \N__33775\,
            I => \N__33743\
        );

    \I__8255\ : InMux
    port map (
            O => \N__33774\,
            I => \N__33743\
        );

    \I__8254\ : InMux
    port map (
            O => \N__33773\,
            I => \N__33738\
        );

    \I__8253\ : InMux
    port map (
            O => \N__33772\,
            I => \N__33738\
        );

    \I__8252\ : InMux
    port map (
            O => \N__33771\,
            I => \N__33735\
        );

    \I__8251\ : Span4Mux_v
    port map (
            O => \N__33768\,
            I => \N__33732\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__33761\,
            I => \N__33729\
        );

    \I__8249\ : InMux
    port map (
            O => \N__33760\,
            I => \N__33726\
        );

    \I__8248\ : Span4Mux_v
    port map (
            O => \N__33757\,
            I => \N__33720\
        );

    \I__8247\ : Span4Mux_h
    port map (
            O => \N__33754\,
            I => \N__33720\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__33749\,
            I => \N__33717\
        );

    \I__8245\ : InMux
    port map (
            O => \N__33748\,
            I => \N__33714\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__33743\,
            I => \N__33710\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__33738\,
            I => \N__33707\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__33735\,
            I => \N__33704\
        );

    \I__8241\ : Span4Mux_h
    port map (
            O => \N__33732\,
            I => \N__33697\
        );

    \I__8240\ : Span4Mux_v
    port map (
            O => \N__33729\,
            I => \N__33697\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__33726\,
            I => \N__33697\
        );

    \I__8238\ : InMux
    port map (
            O => \N__33725\,
            I => \N__33694\
        );

    \I__8237\ : Span4Mux_h
    port map (
            O => \N__33720\,
            I => \N__33687\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__33717\,
            I => \N__33687\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__33714\,
            I => \N__33687\
        );

    \I__8234\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33684\
        );

    \I__8233\ : Span4Mux_h
    port map (
            O => \N__33710\,
            I => \N__33675\
        );

    \I__8232\ : Span4Mux_v
    port map (
            O => \N__33707\,
            I => \N__33675\
        );

    \I__8231\ : Span4Mux_h
    port map (
            O => \N__33704\,
            I => \N__33675\
        );

    \I__8230\ : Span4Mux_v
    port map (
            O => \N__33697\,
            I => \N__33675\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__33694\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__8228\ : Odrv4
    port map (
            O => \N__33687\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__33684\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__8226\ : Odrv4
    port map (
            O => \N__33675\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__8225\ : CascadeMux
    port map (
            O => \N__33666\,
            I => \N__33662\
        );

    \I__8224\ : CascadeMux
    port map (
            O => \N__33665\,
            I => \N__33659\
        );

    \I__8223\ : InMux
    port map (
            O => \N__33662\,
            I => \N__33653\
        );

    \I__8222\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33650\
        );

    \I__8221\ : CascadeMux
    port map (
            O => \N__33658\,
            I => \N__33647\
        );

    \I__8220\ : CascadeMux
    port map (
            O => \N__33657\,
            I => \N__33643\
        );

    \I__8219\ : CascadeMux
    port map (
            O => \N__33656\,
            I => \N__33640\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__33653\,
            I => \N__33635\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__33650\,
            I => \N__33632\
        );

    \I__8216\ : InMux
    port map (
            O => \N__33647\,
            I => \N__33629\
        );

    \I__8215\ : CascadeMux
    port map (
            O => \N__33646\,
            I => \N__33626\
        );

    \I__8214\ : InMux
    port map (
            O => \N__33643\,
            I => \N__33623\
        );

    \I__8213\ : InMux
    port map (
            O => \N__33640\,
            I => \N__33620\
        );

    \I__8212\ : CascadeMux
    port map (
            O => \N__33639\,
            I => \N__33617\
        );

    \I__8211\ : CascadeMux
    port map (
            O => \N__33638\,
            I => \N__33614\
        );

    \I__8210\ : Span4Mux_v
    port map (
            O => \N__33635\,
            I => \N__33605\
        );

    \I__8209\ : Span4Mux_h
    port map (
            O => \N__33632\,
            I => \N__33605\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__33629\,
            I => \N__33605\
        );

    \I__8207\ : InMux
    port map (
            O => \N__33626\,
            I => \N__33602\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__33623\,
            I => \N__33595\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__33620\,
            I => \N__33595\
        );

    \I__8204\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33592\
        );

    \I__8203\ : InMux
    port map (
            O => \N__33614\,
            I => \N__33589\
        );

    \I__8202\ : CascadeMux
    port map (
            O => \N__33613\,
            I => \N__33586\
        );

    \I__8201\ : CascadeMux
    port map (
            O => \N__33612\,
            I => \N__33583\
        );

    \I__8200\ : Span4Mux_v
    port map (
            O => \N__33605\,
            I => \N__33576\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__33602\,
            I => \N__33576\
        );

    \I__8198\ : CascadeMux
    port map (
            O => \N__33601\,
            I => \N__33573\
        );

    \I__8197\ : CascadeMux
    port map (
            O => \N__33600\,
            I => \N__33570\
        );

    \I__8196\ : Span4Mux_v
    port map (
            O => \N__33595\,
            I => \N__33563\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__33592\,
            I => \N__33563\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__33589\,
            I => \N__33563\
        );

    \I__8193\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33560\
        );

    \I__8192\ : InMux
    port map (
            O => \N__33583\,
            I => \N__33557\
        );

    \I__8191\ : CascadeMux
    port map (
            O => \N__33582\,
            I => \N__33554\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__33581\,
            I => \N__33551\
        );

    \I__8189\ : Span4Mux_v
    port map (
            O => \N__33576\,
            I => \N__33547\
        );

    \I__8188\ : InMux
    port map (
            O => \N__33573\,
            I => \N__33544\
        );

    \I__8187\ : InMux
    port map (
            O => \N__33570\,
            I => \N__33541\
        );

    \I__8186\ : Span4Mux_v
    port map (
            O => \N__33563\,
            I => \N__33534\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__33560\,
            I => \N__33534\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__33557\,
            I => \N__33534\
        );

    \I__8183\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33531\
        );

    \I__8182\ : InMux
    port map (
            O => \N__33551\,
            I => \N__33528\
        );

    \I__8181\ : CascadeMux
    port map (
            O => \N__33550\,
            I => \N__33525\
        );

    \I__8180\ : Sp12to4
    port map (
            O => \N__33547\,
            I => \N__33521\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__33544\,
            I => \N__33516\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__33541\,
            I => \N__33516\
        );

    \I__8177\ : Span4Mux_v
    port map (
            O => \N__33534\,
            I => \N__33509\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__33531\,
            I => \N__33509\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__33528\,
            I => \N__33509\
        );

    \I__8174\ : InMux
    port map (
            O => \N__33525\,
            I => \N__33506\
        );

    \I__8173\ : CascadeMux
    port map (
            O => \N__33524\,
            I => \N__33503\
        );

    \I__8172\ : Span12Mux_h
    port map (
            O => \N__33521\,
            I => \N__33500\
        );

    \I__8171\ : Span4Mux_v
    port map (
            O => \N__33516\,
            I => \N__33493\
        );

    \I__8170\ : Span4Mux_v
    port map (
            O => \N__33509\,
            I => \N__33493\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__33506\,
            I => \N__33493\
        );

    \I__8168\ : InMux
    port map (
            O => \N__33503\,
            I => \N__33490\
        );

    \I__8167\ : Odrv12
    port map (
            O => \N__33500\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__8166\ : Odrv4
    port map (
            O => \N__33493\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__33490\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__8164\ : CEMux
    port map (
            O => \N__33483\,
            I => \N__33479\
        );

    \I__8163\ : CEMux
    port map (
            O => \N__33482\,
            I => \N__33476\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__33479\,
            I => \N__33473\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__33476\,
            I => \N__33470\
        );

    \I__8160\ : Span4Mux_v
    port map (
            O => \N__33473\,
            I => \N__33467\
        );

    \I__8159\ : Span4Mux_v
    port map (
            O => \N__33470\,
            I => \N__33464\
        );

    \I__8158\ : Odrv4
    port map (
            O => \N__33467\,
            I => \this_sprites_ram.mem_WE_14\
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__33464\,
            I => \this_sprites_ram.mem_WE_14\
        );

    \I__8156\ : CEMux
    port map (
            O => \N__33459\,
            I => \N__33455\
        );

    \I__8155\ : CEMux
    port map (
            O => \N__33458\,
            I => \N__33452\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__33455\,
            I => \N__33449\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__33452\,
            I => \N__33446\
        );

    \I__8152\ : Span4Mux_v
    port map (
            O => \N__33449\,
            I => \N__33443\
        );

    \I__8151\ : Span4Mux_v
    port map (
            O => \N__33446\,
            I => \N__33440\
        );

    \I__8150\ : Span4Mux_h
    port map (
            O => \N__33443\,
            I => \N__33437\
        );

    \I__8149\ : Odrv4
    port map (
            O => \N__33440\,
            I => \this_sprites_ram.mem_WE_12\
        );

    \I__8148\ : Odrv4
    port map (
            O => \N__33437\,
            I => \this_sprites_ram.mem_WE_12\
        );

    \I__8147\ : CEMux
    port map (
            O => \N__33432\,
            I => \N__33429\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__33429\,
            I => \N__33425\
        );

    \I__8145\ : CEMux
    port map (
            O => \N__33428\,
            I => \N__33422\
        );

    \I__8144\ : Span4Mux_h
    port map (
            O => \N__33425\,
            I => \N__33419\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__33422\,
            I => \N__33416\
        );

    \I__8142\ : Odrv4
    port map (
            O => \N__33419\,
            I => \this_sprites_ram.mem_WE_0\
        );

    \I__8141\ : Odrv4
    port map (
            O => \N__33416\,
            I => \this_sprites_ram.mem_WE_0\
        );

    \I__8140\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33408\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__33408\,
            I => \N__33404\
        );

    \I__8138\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33401\
        );

    \I__8137\ : Span4Mux_v
    port map (
            O => \N__33404\,
            I => \N__33395\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__33401\,
            I => \N__33395\
        );

    \I__8135\ : CascadeMux
    port map (
            O => \N__33400\,
            I => \N__33392\
        );

    \I__8134\ : Span4Mux_v
    port map (
            O => \N__33395\,
            I => \N__33388\
        );

    \I__8133\ : InMux
    port map (
            O => \N__33392\,
            I => \N__33385\
        );

    \I__8132\ : CascadeMux
    port map (
            O => \N__33391\,
            I => \N__33382\
        );

    \I__8131\ : Span4Mux_v
    port map (
            O => \N__33388\,
            I => \N__33379\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__33385\,
            I => \N__33376\
        );

    \I__8129\ : InMux
    port map (
            O => \N__33382\,
            I => \N__33373\
        );

    \I__8128\ : Span4Mux_v
    port map (
            O => \N__33379\,
            I => \N__33364\
        );

    \I__8127\ : Span4Mux_h
    port map (
            O => \N__33376\,
            I => \N__33364\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__33373\,
            I => \N__33364\
        );

    \I__8125\ : CascadeMux
    port map (
            O => \N__33372\,
            I => \N__33361\
        );

    \I__8124\ : InMux
    port map (
            O => \N__33371\,
            I => \N__33356\
        );

    \I__8123\ : Span4Mux_v
    port map (
            O => \N__33364\,
            I => \N__33351\
        );

    \I__8122\ : InMux
    port map (
            O => \N__33361\,
            I => \N__33348\
        );

    \I__8121\ : CascadeMux
    port map (
            O => \N__33360\,
            I => \N__33345\
        );

    \I__8120\ : InMux
    port map (
            O => \N__33359\,
            I => \N__33342\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__33356\,
            I => \N__33339\
        );

    \I__8118\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33334\
        );

    \I__8117\ : InMux
    port map (
            O => \N__33354\,
            I => \N__33334\
        );

    \I__8116\ : Span4Mux_v
    port map (
            O => \N__33351\,
            I => \N__33329\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__33348\,
            I => \N__33329\
        );

    \I__8114\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33326\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__33342\,
            I => \N__33323\
        );

    \I__8112\ : Span4Mux_v
    port map (
            O => \N__33339\,
            I => \N__33320\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__33334\,
            I => \N__33317\
        );

    \I__8110\ : Span4Mux_h
    port map (
            O => \N__33329\,
            I => \N__33312\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__33326\,
            I => \N__33312\
        );

    \I__8108\ : Span12Mux_h
    port map (
            O => \N__33323\,
            I => \N__33308\
        );

    \I__8107\ : Sp12to4
    port map (
            O => \N__33320\,
            I => \N__33305\
        );

    \I__8106\ : Span4Mux_v
    port map (
            O => \N__33317\,
            I => \N__33302\
        );

    \I__8105\ : Span4Mux_v
    port map (
            O => \N__33312\,
            I => \N__33299\
        );

    \I__8104\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33296\
        );

    \I__8103\ : Span12Mux_v
    port map (
            O => \N__33308\,
            I => \N__33293\
        );

    \I__8102\ : Span12Mux_v
    port map (
            O => \N__33305\,
            I => \N__33286\
        );

    \I__8101\ : Sp12to4
    port map (
            O => \N__33302\,
            I => \N__33286\
        );

    \I__8100\ : Sp12to4
    port map (
            O => \N__33299\,
            I => \N__33286\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__33296\,
            I => \N__33283\
        );

    \I__8098\ : Span12Mux_v
    port map (
            O => \N__33293\,
            I => \N__33280\
        );

    \I__8097\ : Span12Mux_h
    port map (
            O => \N__33286\,
            I => \N__33277\
        );

    \I__8096\ : Span4Mux_v
    port map (
            O => \N__33283\,
            I => \N__33274\
        );

    \I__8095\ : Odrv12
    port map (
            O => \N__33280\,
            I => port_data_c_1
        );

    \I__8094\ : Odrv12
    port map (
            O => \N__33277\,
            I => port_data_c_1
        );

    \I__8093\ : Odrv4
    port map (
            O => \N__33274\,
            I => port_data_c_1
        );

    \I__8092\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33264\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__33264\,
            I => \this_vga_signals_M_this_external_address_q_3_i_0_0_15\
        );

    \I__8090\ : CascadeMux
    port map (
            O => \N__33261\,
            I => \N__33258\
        );

    \I__8089\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33252\
        );

    \I__8088\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33252\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__33252\,
            I => \N__33247\
        );

    \I__8086\ : CascadeMux
    port map (
            O => \N__33251\,
            I => \N__33241\
        );

    \I__8085\ : InMux
    port map (
            O => \N__33250\,
            I => \N__33236\
        );

    \I__8084\ : Span4Mux_v
    port map (
            O => \N__33247\,
            I => \N__33233\
        );

    \I__8083\ : InMux
    port map (
            O => \N__33246\,
            I => \N__33228\
        );

    \I__8082\ : InMux
    port map (
            O => \N__33245\,
            I => \N__33228\
        );

    \I__8081\ : InMux
    port map (
            O => \N__33244\,
            I => \N__33224\
        );

    \I__8080\ : InMux
    port map (
            O => \N__33241\,
            I => \N__33219\
        );

    \I__8079\ : InMux
    port map (
            O => \N__33240\,
            I => \N__33219\
        );

    \I__8078\ : InMux
    port map (
            O => \N__33239\,
            I => \N__33216\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__33236\,
            I => \N__33211\
        );

    \I__8076\ : Span4Mux_v
    port map (
            O => \N__33233\,
            I => \N__33211\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__33228\,
            I => \N__33208\
        );

    \I__8074\ : InMux
    port map (
            O => \N__33227\,
            I => \N__33205\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__33224\,
            I => \N__33202\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__33219\,
            I => \N__33199\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__33216\,
            I => \N__33196\
        );

    \I__8070\ : Span4Mux_v
    port map (
            O => \N__33211\,
            I => \N__33193\
        );

    \I__8069\ : Span12Mux_v
    port map (
            O => \N__33208\,
            I => \N__33190\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__33205\,
            I => \N__33183\
        );

    \I__8067\ : Span4Mux_v
    port map (
            O => \N__33202\,
            I => \N__33183\
        );

    \I__8066\ : Span4Mux_v
    port map (
            O => \N__33199\,
            I => \N__33183\
        );

    \I__8065\ : Odrv12
    port map (
            O => \N__33196\,
            I => \N_661\
        );

    \I__8064\ : Odrv4
    port map (
            O => \N__33193\,
            I => \N_661\
        );

    \I__8063\ : Odrv12
    port map (
            O => \N__33190\,
            I => \N_661\
        );

    \I__8062\ : Odrv4
    port map (
            O => \N__33183\,
            I => \N_661\
        );

    \I__8061\ : CEMux
    port map (
            O => \N__33174\,
            I => \N__33171\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__33171\,
            I => \N__33167\
        );

    \I__8059\ : CEMux
    port map (
            O => \N__33170\,
            I => \N__33164\
        );

    \I__8058\ : Span4Mux_v
    port map (
            O => \N__33167\,
            I => \N__33161\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__33164\,
            I => \N__33158\
        );

    \I__8056\ : Odrv4
    port map (
            O => \N__33161\,
            I => \this_sprites_ram.mem_WE_2\
        );

    \I__8055\ : Odrv4
    port map (
            O => \N__33158\,
            I => \this_sprites_ram.mem_WE_2\
        );

    \I__8054\ : InMux
    port map (
            O => \N__33153\,
            I => \N__33150\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__33150\,
            I => \this_ppu.M_this_oam_ram_read_data_iZ0Z_8\
        );

    \I__8052\ : InMux
    port map (
            O => \N__33147\,
            I => \N__33144\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__33144\,
            I => \N__33141\
        );

    \I__8050\ : Odrv12
    port map (
            O => \N__33141\,
            I => \M_this_oam_ram_read_data_i_9\
        );

    \I__8049\ : InMux
    port map (
            O => \N__33138\,
            I => \this_ppu.un2_hscroll_cry_0\
        );

    \I__8048\ : CascadeMux
    port map (
            O => \N__33135\,
            I => \N__33132\
        );

    \I__8047\ : InMux
    port map (
            O => \N__33132\,
            I => \N__33127\
        );

    \I__8046\ : InMux
    port map (
            O => \N__33131\,
            I => \N__33124\
        );

    \I__8045\ : CascadeMux
    port map (
            O => \N__33130\,
            I => \N__33121\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__33127\,
            I => \N__33118\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__33124\,
            I => \N__33115\
        );

    \I__8042\ : InMux
    port map (
            O => \N__33121\,
            I => \N__33112\
        );

    \I__8041\ : Span4Mux_h
    port map (
            O => \N__33118\,
            I => \N__33109\
        );

    \I__8040\ : Span4Mux_v
    port map (
            O => \N__33115\,
            I => \N__33106\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__33112\,
            I => \N__33103\
        );

    \I__8038\ : Span4Mux_h
    port map (
            O => \N__33109\,
            I => \N__33100\
        );

    \I__8037\ : Odrv4
    port map (
            O => \N__33106\,
            I => \M_this_oam_ram_read_data_10\
        );

    \I__8036\ : Odrv12
    port map (
            O => \N__33103\,
            I => \M_this_oam_ram_read_data_10\
        );

    \I__8035\ : Odrv4
    port map (
            O => \N__33100\,
            I => \M_this_oam_ram_read_data_10\
        );

    \I__8034\ : InMux
    port map (
            O => \N__33093\,
            I => \this_ppu.un2_hscroll_cry_1\
        );

    \I__8033\ : InMux
    port map (
            O => \N__33090\,
            I => \N__33087\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__33087\,
            I => \N__33084\
        );

    \I__8031\ : Span4Mux_v
    port map (
            O => \N__33084\,
            I => \N__33081\
        );

    \I__8030\ : Odrv4
    port map (
            O => \N__33081\,
            I => \M_this_oam_ram_write_data_26\
        );

    \I__8029\ : InMux
    port map (
            O => \N__33078\,
            I => \N__33075\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__33075\,
            I => \N__33072\
        );

    \I__8027\ : Span4Mux_h
    port map (
            O => \N__33072\,
            I => \N__33069\
        );

    \I__8026\ : Odrv4
    port map (
            O => \N__33069\,
            I => \M_this_oam_ram_write_data_19\
        );

    \I__8025\ : CascadeMux
    port map (
            O => \N__33066\,
            I => \N__33061\
        );

    \I__8024\ : CascadeMux
    port map (
            O => \N__33065\,
            I => \N__33057\
        );

    \I__8023\ : InMux
    port map (
            O => \N__33064\,
            I => \N__33054\
        );

    \I__8022\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33051\
        );

    \I__8021\ : InMux
    port map (
            O => \N__33060\,
            I => \N__33048\
        );

    \I__8020\ : InMux
    port map (
            O => \N__33057\,
            I => \N__33045\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__33054\,
            I => \N__33040\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__33051\,
            I => \N__33040\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__33048\,
            I => \N__33036\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__33045\,
            I => \N__33033\
        );

    \I__8015\ : Span4Mux_v
    port map (
            O => \N__33040\,
            I => \N__33028\
        );

    \I__8014\ : InMux
    port map (
            O => \N__33039\,
            I => \N__33025\
        );

    \I__8013\ : Span4Mux_v
    port map (
            O => \N__33036\,
            I => \N__33022\
        );

    \I__8012\ : Span12Mux_v
    port map (
            O => \N__33033\,
            I => \N__33019\
        );

    \I__8011\ : InMux
    port map (
            O => \N__33032\,
            I => \N__33016\
        );

    \I__8010\ : InMux
    port map (
            O => \N__33031\,
            I => \N__33013\
        );

    \I__8009\ : Span4Mux_h
    port map (
            O => \N__33028\,
            I => \N__33010\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__33025\,
            I => \N__33005\
        );

    \I__8007\ : Span4Mux_v
    port map (
            O => \N__33022\,
            I => \N__33005\
        );

    \I__8006\ : Odrv12
    port map (
            O => \N__33019\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__33016\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__33013\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__8003\ : Odrv4
    port map (
            O => \N__33010\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__8002\ : Odrv4
    port map (
            O => \N__33005\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__8001\ : InMux
    port map (
            O => \N__32994\,
            I => \N__32991\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__32991\,
            I => \this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0\
        );

    \I__7999\ : CascadeMux
    port map (
            O => \N__32988\,
            I => \N__32985\
        );

    \I__7998\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32978\
        );

    \I__7997\ : CascadeMux
    port map (
            O => \N__32984\,
            I => \N__32975\
        );

    \I__7996\ : CascadeMux
    port map (
            O => \N__32983\,
            I => \N__32972\
        );

    \I__7995\ : CascadeMux
    port map (
            O => \N__32982\,
            I => \N__32968\
        );

    \I__7994\ : CascadeMux
    port map (
            O => \N__32981\,
            I => \N__32965\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__32978\,
            I => \N__32960\
        );

    \I__7992\ : InMux
    port map (
            O => \N__32975\,
            I => \N__32957\
        );

    \I__7991\ : InMux
    port map (
            O => \N__32972\,
            I => \N__32954\
        );

    \I__7990\ : CascadeMux
    port map (
            O => \N__32971\,
            I => \N__32951\
        );

    \I__7989\ : InMux
    port map (
            O => \N__32968\,
            I => \N__32948\
        );

    \I__7988\ : InMux
    port map (
            O => \N__32965\,
            I => \N__32945\
        );

    \I__7987\ : CascadeMux
    port map (
            O => \N__32964\,
            I => \N__32942\
        );

    \I__7986\ : CascadeMux
    port map (
            O => \N__32963\,
            I => \N__32939\
        );

    \I__7985\ : Span4Mux_v
    port map (
            O => \N__32960\,
            I => \N__32930\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__32957\,
            I => \N__32930\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__32954\,
            I => \N__32930\
        );

    \I__7982\ : InMux
    port map (
            O => \N__32951\,
            I => \N__32927\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__32948\,
            I => \N__32922\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__32945\,
            I => \N__32922\
        );

    \I__7979\ : InMux
    port map (
            O => \N__32942\,
            I => \N__32919\
        );

    \I__7978\ : InMux
    port map (
            O => \N__32939\,
            I => \N__32916\
        );

    \I__7977\ : CascadeMux
    port map (
            O => \N__32938\,
            I => \N__32913\
        );

    \I__7976\ : CascadeMux
    port map (
            O => \N__32937\,
            I => \N__32910\
        );

    \I__7975\ : Span4Mux_v
    port map (
            O => \N__32930\,
            I => \N__32903\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__32927\,
            I => \N__32903\
        );

    \I__7973\ : Span4Mux_v
    port map (
            O => \N__32922\,
            I => \N__32900\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__32919\,
            I => \N__32895\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__32916\,
            I => \N__32895\
        );

    \I__7970\ : InMux
    port map (
            O => \N__32913\,
            I => \N__32892\
        );

    \I__7969\ : InMux
    port map (
            O => \N__32910\,
            I => \N__32889\
        );

    \I__7968\ : CascadeMux
    port map (
            O => \N__32909\,
            I => \N__32886\
        );

    \I__7967\ : CascadeMux
    port map (
            O => \N__32908\,
            I => \N__32883\
        );

    \I__7966\ : Span4Mux_v
    port map (
            O => \N__32903\,
            I => \N__32879\
        );

    \I__7965\ : Span4Mux_v
    port map (
            O => \N__32900\,
            I => \N__32869\
        );

    \I__7964\ : Span4Mux_v
    port map (
            O => \N__32895\,
            I => \N__32869\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__32892\,
            I => \N__32869\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__32889\,
            I => \N__32869\
        );

    \I__7961\ : InMux
    port map (
            O => \N__32886\,
            I => \N__32866\
        );

    \I__7960\ : InMux
    port map (
            O => \N__32883\,
            I => \N__32863\
        );

    \I__7959\ : CascadeMux
    port map (
            O => \N__32882\,
            I => \N__32860\
        );

    \I__7958\ : Span4Mux_v
    port map (
            O => \N__32879\,
            I => \N__32857\
        );

    \I__7957\ : CascadeMux
    port map (
            O => \N__32878\,
            I => \N__32854\
        );

    \I__7956\ : Span4Mux_v
    port map (
            O => \N__32869\,
            I => \N__32847\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__32866\,
            I => \N__32847\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__32863\,
            I => \N__32847\
        );

    \I__7953\ : InMux
    port map (
            O => \N__32860\,
            I => \N__32844\
        );

    \I__7952\ : Sp12to4
    port map (
            O => \N__32857\,
            I => \N__32839\
        );

    \I__7951\ : InMux
    port map (
            O => \N__32854\,
            I => \N__32836\
        );

    \I__7950\ : Span4Mux_v
    port map (
            O => \N__32847\,
            I => \N__32831\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__32844\,
            I => \N__32831\
        );

    \I__7948\ : CascadeMux
    port map (
            O => \N__32843\,
            I => \N__32828\
        );

    \I__7947\ : CascadeMux
    port map (
            O => \N__32842\,
            I => \N__32825\
        );

    \I__7946\ : Span12Mux_h
    port map (
            O => \N__32839\,
            I => \N__32822\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__32836\,
            I => \N__32819\
        );

    \I__7944\ : Span4Mux_v
    port map (
            O => \N__32831\,
            I => \N__32816\
        );

    \I__7943\ : InMux
    port map (
            O => \N__32828\,
            I => \N__32813\
        );

    \I__7942\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32810\
        );

    \I__7941\ : Odrv12
    port map (
            O => \N__32822\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__7940\ : Odrv4
    port map (
            O => \N__32819\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__7939\ : Odrv4
    port map (
            O => \N__32816\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__32813\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__32810\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__7936\ : InMux
    port map (
            O => \N__32799\,
            I => \N__32795\
        );

    \I__7935\ : InMux
    port map (
            O => \N__32798\,
            I => \N__32790\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__32795\,
            I => \N__32787\
        );

    \I__7933\ : InMux
    port map (
            O => \N__32794\,
            I => \N__32784\
        );

    \I__7932\ : InMux
    port map (
            O => \N__32793\,
            I => \N__32781\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__32790\,
            I => \N__32778\
        );

    \I__7930\ : Span4Mux_h
    port map (
            O => \N__32787\,
            I => \N__32775\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__32784\,
            I => \N__32770\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__32781\,
            I => \N__32770\
        );

    \I__7927\ : Span4Mux_h
    port map (
            O => \N__32778\,
            I => \N__32767\
        );

    \I__7926\ : Span4Mux_h
    port map (
            O => \N__32775\,
            I => \N__32764\
        );

    \I__7925\ : Span4Mux_v
    port map (
            O => \N__32770\,
            I => \N__32761\
        );

    \I__7924\ : Odrv4
    port map (
            O => \N__32767\,
            I => \M_this_oam_ram_read_data_8\
        );

    \I__7923\ : Odrv4
    port map (
            O => \N__32764\,
            I => \M_this_oam_ram_read_data_8\
        );

    \I__7922\ : Odrv4
    port map (
            O => \N__32761\,
            I => \M_this_oam_ram_read_data_8\
        );

    \I__7921\ : CascadeMux
    port map (
            O => \N__32754\,
            I => \N__32751\
        );

    \I__7920\ : InMux
    port map (
            O => \N__32751\,
            I => \N__32748\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__32748\,
            I => \N__32744\
        );

    \I__7918\ : CascadeMux
    port map (
            O => \N__32747\,
            I => \N__32740\
        );

    \I__7917\ : Span4Mux_v
    port map (
            O => \N__32744\,
            I => \N__32734\
        );

    \I__7916\ : InMux
    port map (
            O => \N__32743\,
            I => \N__32731\
        );

    \I__7915\ : InMux
    port map (
            O => \N__32740\,
            I => \N__32728\
        );

    \I__7914\ : InMux
    port map (
            O => \N__32739\,
            I => \N__32725\
        );

    \I__7913\ : CascadeMux
    port map (
            O => \N__32738\,
            I => \N__32722\
        );

    \I__7912\ : CascadeMux
    port map (
            O => \N__32737\,
            I => \N__32717\
        );

    \I__7911\ : Span4Mux_h
    port map (
            O => \N__32734\,
            I => \N__32714\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__32731\,
            I => \N__32711\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__32728\,
            I => \N__32706\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__32725\,
            I => \N__32706\
        );

    \I__7907\ : InMux
    port map (
            O => \N__32722\,
            I => \N__32701\
        );

    \I__7906\ : InMux
    port map (
            O => \N__32721\,
            I => \N__32701\
        );

    \I__7905\ : InMux
    port map (
            O => \N__32720\,
            I => \N__32698\
        );

    \I__7904\ : InMux
    port map (
            O => \N__32717\,
            I => \N__32695\
        );

    \I__7903\ : Span4Mux_h
    port map (
            O => \N__32714\,
            I => \N__32692\
        );

    \I__7902\ : Span4Mux_v
    port map (
            O => \N__32711\,
            I => \N__32689\
        );

    \I__7901\ : Span12Mux_v
    port map (
            O => \N__32706\,
            I => \N__32686\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__32701\,
            I => \N__32681\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__32698\,
            I => \N__32681\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__32695\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__7897\ : Odrv4
    port map (
            O => \N__32692\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__7896\ : Odrv4
    port map (
            O => \N__32689\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__7895\ : Odrv12
    port map (
            O => \N__32686\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__7894\ : Odrv12
    port map (
            O => \N__32681\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__7893\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32667\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__32667\,
            I => \N__32664\
        );

    \I__7891\ : Odrv4
    port map (
            O => \N__32664\,
            I => \this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0\
        );

    \I__7890\ : CascadeMux
    port map (
            O => \N__32661\,
            I => \N__32657\
        );

    \I__7889\ : CascadeMux
    port map (
            O => \N__32660\,
            I => \N__32654\
        );

    \I__7888\ : InMux
    port map (
            O => \N__32657\,
            I => \N__32645\
        );

    \I__7887\ : InMux
    port map (
            O => \N__32654\,
            I => \N__32642\
        );

    \I__7886\ : CascadeMux
    port map (
            O => \N__32653\,
            I => \N__32639\
        );

    \I__7885\ : CascadeMux
    port map (
            O => \N__32652\,
            I => \N__32636\
        );

    \I__7884\ : CascadeMux
    port map (
            O => \N__32651\,
            I => \N__32631\
        );

    \I__7883\ : CascadeMux
    port map (
            O => \N__32650\,
            I => \N__32628\
        );

    \I__7882\ : CascadeMux
    port map (
            O => \N__32649\,
            I => \N__32625\
        );

    \I__7881\ : CascadeMux
    port map (
            O => \N__32648\,
            I => \N__32622\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__32645\,
            I => \N__32616\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__32642\,
            I => \N__32616\
        );

    \I__7878\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32613\
        );

    \I__7877\ : InMux
    port map (
            O => \N__32636\,
            I => \N__32610\
        );

    \I__7876\ : CascadeMux
    port map (
            O => \N__32635\,
            I => \N__32607\
        );

    \I__7875\ : CascadeMux
    port map (
            O => \N__32634\,
            I => \N__32604\
        );

    \I__7874\ : InMux
    port map (
            O => \N__32631\,
            I => \N__32599\
        );

    \I__7873\ : InMux
    port map (
            O => \N__32628\,
            I => \N__32596\
        );

    \I__7872\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32593\
        );

    \I__7871\ : InMux
    port map (
            O => \N__32622\,
            I => \N__32590\
        );

    \I__7870\ : CascadeMux
    port map (
            O => \N__32621\,
            I => \N__32587\
        );

    \I__7869\ : Span4Mux_v
    port map (
            O => \N__32616\,
            I => \N__32580\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__32613\,
            I => \N__32580\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__32610\,
            I => \N__32580\
        );

    \I__7866\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32577\
        );

    \I__7865\ : InMux
    port map (
            O => \N__32604\,
            I => \N__32574\
        );

    \I__7864\ : CascadeMux
    port map (
            O => \N__32603\,
            I => \N__32571\
        );

    \I__7863\ : CascadeMux
    port map (
            O => \N__32602\,
            I => \N__32568\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__32599\,
            I => \N__32557\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__32596\,
            I => \N__32557\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__32593\,
            I => \N__32557\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__32590\,
            I => \N__32557\
        );

    \I__7858\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32554\
        );

    \I__7857\ : Span4Mux_v
    port map (
            O => \N__32580\,
            I => \N__32547\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__32577\,
            I => \N__32547\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__32574\,
            I => \N__32547\
        );

    \I__7854\ : InMux
    port map (
            O => \N__32571\,
            I => \N__32544\
        );

    \I__7853\ : InMux
    port map (
            O => \N__32568\,
            I => \N__32541\
        );

    \I__7852\ : CascadeMux
    port map (
            O => \N__32567\,
            I => \N__32538\
        );

    \I__7851\ : CascadeMux
    port map (
            O => \N__32566\,
            I => \N__32535\
        );

    \I__7850\ : Span12Mux_v
    port map (
            O => \N__32557\,
            I => \N__32531\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__32554\,
            I => \N__32528\
        );

    \I__7848\ : Span4Mux_v
    port map (
            O => \N__32547\,
            I => \N__32521\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__32544\,
            I => \N__32521\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__32541\,
            I => \N__32521\
        );

    \I__7845\ : InMux
    port map (
            O => \N__32538\,
            I => \N__32518\
        );

    \I__7844\ : InMux
    port map (
            O => \N__32535\,
            I => \N__32515\
        );

    \I__7843\ : CascadeMux
    port map (
            O => \N__32534\,
            I => \N__32512\
        );

    \I__7842\ : Span12Mux_h
    port map (
            O => \N__32531\,
            I => \N__32509\
        );

    \I__7841\ : Span4Mux_v
    port map (
            O => \N__32528\,
            I => \N__32502\
        );

    \I__7840\ : Span4Mux_v
    port map (
            O => \N__32521\,
            I => \N__32502\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__32518\,
            I => \N__32502\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__32515\,
            I => \N__32499\
        );

    \I__7837\ : InMux
    port map (
            O => \N__32512\,
            I => \N__32496\
        );

    \I__7836\ : Odrv12
    port map (
            O => \N__32509\,
            I => \M_this_ppu_sprites_addr_2\
        );

    \I__7835\ : Odrv4
    port map (
            O => \N__32502\,
            I => \M_this_ppu_sprites_addr_2\
        );

    \I__7834\ : Odrv4
    port map (
            O => \N__32499\,
            I => \M_this_ppu_sprites_addr_2\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__32496\,
            I => \M_this_ppu_sprites_addr_2\
        );

    \I__7832\ : InMux
    port map (
            O => \N__32487\,
            I => \N__32484\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__32484\,
            I => \N__32481\
        );

    \I__7830\ : Span4Mux_v
    port map (
            O => \N__32481\,
            I => \N__32478\
        );

    \I__7829\ : Odrv4
    port map (
            O => \N__32478\,
            I => \M_this_data_tmp_qZ0Z_22\
        );

    \I__7828\ : InMux
    port map (
            O => \N__32475\,
            I => \N__32472\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__32472\,
            I => \N__32469\
        );

    \I__7826\ : Odrv4
    port map (
            O => \N__32469\,
            I => \M_this_oam_ram_write_data_22\
        );

    \I__7825\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32463\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__32463\,
            I => \M_this_oam_ram_write_data_31\
        );

    \I__7823\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32457\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__32457\,
            I => \M_this_data_tmp_qZ0Z_18\
        );

    \I__7821\ : InMux
    port map (
            O => \N__32454\,
            I => \N__32451\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__32451\,
            I => \M_this_data_tmp_qZ0Z_20\
        );

    \I__7819\ : InMux
    port map (
            O => \N__32448\,
            I => \N__32445\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__32445\,
            I => \N__32438\
        );

    \I__7817\ : InMux
    port map (
            O => \N__32444\,
            I => \N__32435\
        );

    \I__7816\ : InMux
    port map (
            O => \N__32443\,
            I => \N__32430\
        );

    \I__7815\ : InMux
    port map (
            O => \N__32442\,
            I => \N__32430\
        );

    \I__7814\ : CascadeMux
    port map (
            O => \N__32441\,
            I => \N__32427\
        );

    \I__7813\ : Span4Mux_v
    port map (
            O => \N__32438\,
            I => \N__32421\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__32435\,
            I => \N__32421\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__32430\,
            I => \N__32418\
        );

    \I__7810\ : InMux
    port map (
            O => \N__32427\,
            I => \N__32414\
        );

    \I__7809\ : CascadeMux
    port map (
            O => \N__32426\,
            I => \N__32410\
        );

    \I__7808\ : Span4Mux_v
    port map (
            O => \N__32421\,
            I => \N__32407\
        );

    \I__7807\ : Span4Mux_v
    port map (
            O => \N__32418\,
            I => \N__32402\
        );

    \I__7806\ : InMux
    port map (
            O => \N__32417\,
            I => \N__32399\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__32414\,
            I => \N__32396\
        );

    \I__7804\ : CascadeMux
    port map (
            O => \N__32413\,
            I => \N__32393\
        );

    \I__7803\ : InMux
    port map (
            O => \N__32410\,
            I => \N__32390\
        );

    \I__7802\ : Span4Mux_v
    port map (
            O => \N__32407\,
            I => \N__32387\
        );

    \I__7801\ : InMux
    port map (
            O => \N__32406\,
            I => \N__32384\
        );

    \I__7800\ : CascadeMux
    port map (
            O => \N__32405\,
            I => \N__32380\
        );

    \I__7799\ : Span4Mux_v
    port map (
            O => \N__32402\,
            I => \N__32377\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__32399\,
            I => \N__32374\
        );

    \I__7797\ : Span4Mux_v
    port map (
            O => \N__32396\,
            I => \N__32371\
        );

    \I__7796\ : InMux
    port map (
            O => \N__32393\,
            I => \N__32368\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__32390\,
            I => \N__32365\
        );

    \I__7794\ : Span4Mux_v
    port map (
            O => \N__32387\,
            I => \N__32360\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__32384\,
            I => \N__32360\
        );

    \I__7792\ : InMux
    port map (
            O => \N__32383\,
            I => \N__32357\
        );

    \I__7791\ : InMux
    port map (
            O => \N__32380\,
            I => \N__32354\
        );

    \I__7790\ : Sp12to4
    port map (
            O => \N__32377\,
            I => \N__32351\
        );

    \I__7789\ : Span4Mux_v
    port map (
            O => \N__32374\,
            I => \N__32348\
        );

    \I__7788\ : Span4Mux_h
    port map (
            O => \N__32371\,
            I => \N__32343\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__32368\,
            I => \N__32343\
        );

    \I__7786\ : Span4Mux_v
    port map (
            O => \N__32365\,
            I => \N__32340\
        );

    \I__7785\ : Span4Mux_v
    port map (
            O => \N__32360\,
            I => \N__32337\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__32357\,
            I => \N__32332\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__32354\,
            I => \N__32332\
        );

    \I__7782\ : Span12Mux_h
    port map (
            O => \N__32351\,
            I => \N__32329\
        );

    \I__7781\ : Sp12to4
    port map (
            O => \N__32348\,
            I => \N__32326\
        );

    \I__7780\ : Sp12to4
    port map (
            O => \N__32343\,
            I => \N__32323\
        );

    \I__7779\ : Span4Mux_h
    port map (
            O => \N__32340\,
            I => \N__32318\
        );

    \I__7778\ : Span4Mux_v
    port map (
            O => \N__32337\,
            I => \N__32318\
        );

    \I__7777\ : Span4Mux_v
    port map (
            O => \N__32332\,
            I => \N__32315\
        );

    \I__7776\ : Span12Mux_v
    port map (
            O => \N__32329\,
            I => \N__32312\
        );

    \I__7775\ : Span12Mux_h
    port map (
            O => \N__32326\,
            I => \N__32303\
        );

    \I__7774\ : Span12Mux_v
    port map (
            O => \N__32323\,
            I => \N__32303\
        );

    \I__7773\ : Sp12to4
    port map (
            O => \N__32318\,
            I => \N__32303\
        );

    \I__7772\ : Sp12to4
    port map (
            O => \N__32315\,
            I => \N__32303\
        );

    \I__7771\ : Odrv12
    port map (
            O => \N__32312\,
            I => port_data_c_4
        );

    \I__7770\ : Odrv12
    port map (
            O => \N__32303\,
            I => port_data_c_4
        );

    \I__7769\ : InMux
    port map (
            O => \N__32298\,
            I => \N__32295\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__32295\,
            I => \N__32292\
        );

    \I__7767\ : Odrv4
    port map (
            O => \N__32292\,
            I => \M_this_oam_ram_write_data_28\
        );

    \I__7766\ : InMux
    port map (
            O => \N__32289\,
            I => \N__32286\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__32286\,
            I => \N__32283\
        );

    \I__7764\ : Odrv4
    port map (
            O => \N__32283\,
            I => \M_this_data_tmp_qZ0Z_21\
        );

    \I__7763\ : InMux
    port map (
            O => \N__32280\,
            I => \N__32277\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__32277\,
            I => \M_this_oam_ram_write_data_21\
        );

    \I__7761\ : CascadeMux
    port map (
            O => \N__32274\,
            I => \N__32271\
        );

    \I__7760\ : CascadeBuf
    port map (
            O => \N__32271\,
            I => \N__32268\
        );

    \I__7759\ : CascadeMux
    port map (
            O => \N__32268\,
            I => \N__32263\
        );

    \I__7758\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32258\
        );

    \I__7757\ : InMux
    port map (
            O => \N__32266\,
            I => \N__32258\
        );

    \I__7756\ : InMux
    port map (
            O => \N__32263\,
            I => \N__32255\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__32258\,
            I => \M_this_oam_address_qZ0Z_6\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__32255\,
            I => \M_this_oam_address_qZ0Z_6\
        );

    \I__7753\ : InMux
    port map (
            O => \N__32250\,
            I => \N__32244\
        );

    \I__7752\ : InMux
    port map (
            O => \N__32249\,
            I => \N__32244\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__32244\,
            I => \un1_M_this_oam_address_q_c6\
        );

    \I__7750\ : CascadeMux
    port map (
            O => \N__32241\,
            I => \N__32238\
        );

    \I__7749\ : CascadeBuf
    port map (
            O => \N__32238\,
            I => \N__32234\
        );

    \I__7748\ : CascadeMux
    port map (
            O => \N__32237\,
            I => \N__32231\
        );

    \I__7747\ : CascadeMux
    port map (
            O => \N__32234\,
            I => \N__32228\
        );

    \I__7746\ : InMux
    port map (
            O => \N__32231\,
            I => \N__32225\
        );

    \I__7745\ : InMux
    port map (
            O => \N__32228\,
            I => \N__32222\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__32225\,
            I => \M_this_oam_address_qZ0Z_7\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__32222\,
            I => \M_this_oam_address_qZ0Z_7\
        );

    \I__7742\ : SRMux
    port map (
            O => \N__32217\,
            I => \N__32172\
        );

    \I__7741\ : SRMux
    port map (
            O => \N__32216\,
            I => \N__32172\
        );

    \I__7740\ : SRMux
    port map (
            O => \N__32215\,
            I => \N__32172\
        );

    \I__7739\ : SRMux
    port map (
            O => \N__32214\,
            I => \N__32172\
        );

    \I__7738\ : SRMux
    port map (
            O => \N__32213\,
            I => \N__32172\
        );

    \I__7737\ : SRMux
    port map (
            O => \N__32212\,
            I => \N__32172\
        );

    \I__7736\ : SRMux
    port map (
            O => \N__32211\,
            I => \N__32172\
        );

    \I__7735\ : SRMux
    port map (
            O => \N__32210\,
            I => \N__32172\
        );

    \I__7734\ : SRMux
    port map (
            O => \N__32209\,
            I => \N__32172\
        );

    \I__7733\ : SRMux
    port map (
            O => \N__32208\,
            I => \N__32172\
        );

    \I__7732\ : SRMux
    port map (
            O => \N__32207\,
            I => \N__32172\
        );

    \I__7731\ : SRMux
    port map (
            O => \N__32206\,
            I => \N__32172\
        );

    \I__7730\ : SRMux
    port map (
            O => \N__32205\,
            I => \N__32172\
        );

    \I__7729\ : SRMux
    port map (
            O => \N__32204\,
            I => \N__32172\
        );

    \I__7728\ : SRMux
    port map (
            O => \N__32203\,
            I => \N__32172\
        );

    \I__7727\ : GlobalMux
    port map (
            O => \N__32172\,
            I => \N__32169\
        );

    \I__7726\ : gio2CtrlBuf
    port map (
            O => \N__32169\,
            I => \N_404_g\
        );

    \I__7725\ : InMux
    port map (
            O => \N__32166\,
            I => \N__32163\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__32163\,
            I => \N__32160\
        );

    \I__7723\ : Odrv12
    port map (
            O => \N__32160\,
            I => \M_this_data_tmp_qZ0Z_9\
        );

    \I__7722\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32154\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__32154\,
            I => \N__32151\
        );

    \I__7720\ : Odrv4
    port map (
            O => \N__32151\,
            I => \M_this_data_tmp_qZ0Z_12\
        );

    \I__7719\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32145\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__32145\,
            I => \M_this_oam_ram_write_data_12\
        );

    \I__7717\ : CascadeMux
    port map (
            O => \N__32142\,
            I => \N__32139\
        );

    \I__7716\ : InMux
    port map (
            O => \N__32139\,
            I => \N__32134\
        );

    \I__7715\ : InMux
    port map (
            O => \N__32138\,
            I => \N__32129\
        );

    \I__7714\ : InMux
    port map (
            O => \N__32137\,
            I => \N__32129\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__32134\,
            I => \N__32125\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__32129\,
            I => \N__32122\
        );

    \I__7711\ : InMux
    port map (
            O => \N__32128\,
            I => \N__32119\
        );

    \I__7710\ : Span12Mux_h
    port map (
            O => \N__32125\,
            I => \N__32116\
        );

    \I__7709\ : Span4Mux_h
    port map (
            O => \N__32122\,
            I => \N__32113\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__32119\,
            I => \N__32110\
        );

    \I__7707\ : Odrv12
    port map (
            O => \N__32116\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__7706\ : Odrv4
    port map (
            O => \N__32113\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__7705\ : Odrv4
    port map (
            O => \N__32110\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__7704\ : InMux
    port map (
            O => \N__32103\,
            I => \N__32100\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__32100\,
            I => \N__32094\
        );

    \I__7702\ : InMux
    port map (
            O => \N__32099\,
            I => \N__32089\
        );

    \I__7701\ : InMux
    port map (
            O => \N__32098\,
            I => \N__32089\
        );

    \I__7700\ : InMux
    port map (
            O => \N__32097\,
            I => \N__32086\
        );

    \I__7699\ : Span4Mux_v
    port map (
            O => \N__32094\,
            I => \N__32081\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__32089\,
            I => \N__32081\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__32086\,
            I => \N__32078\
        );

    \I__7696\ : Span4Mux_h
    port map (
            O => \N__32081\,
            I => \N__32075\
        );

    \I__7695\ : Odrv4
    port map (
            O => \N__32078\,
            I => \M_this_oam_ram_read_data_20\
        );

    \I__7694\ : Odrv4
    port map (
            O => \N__32075\,
            I => \M_this_oam_ram_read_data_20\
        );

    \I__7693\ : InMux
    port map (
            O => \N__32070\,
            I => \N__32067\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__32067\,
            I => \N__32060\
        );

    \I__7691\ : InMux
    port map (
            O => \N__32066\,
            I => \N__32057\
        );

    \I__7690\ : InMux
    port map (
            O => \N__32065\,
            I => \N__32052\
        );

    \I__7689\ : InMux
    port map (
            O => \N__32064\,
            I => \N__32052\
        );

    \I__7688\ : InMux
    port map (
            O => \N__32063\,
            I => \N__32049\
        );

    \I__7687\ : Span4Mux_v
    port map (
            O => \N__32060\,
            I => \N__32042\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__32057\,
            I => \N__32042\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__32052\,
            I => \N__32042\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__32049\,
            I => \N__32039\
        );

    \I__7683\ : Span4Mux_h
    port map (
            O => \N__32042\,
            I => \N__32036\
        );

    \I__7682\ : Odrv4
    port map (
            O => \N__32039\,
            I => \M_this_oam_ram_read_data_19\
        );

    \I__7681\ : Odrv4
    port map (
            O => \N__32036\,
            I => \M_this_oam_ram_read_data_19\
        );

    \I__7680\ : InMux
    port map (
            O => \N__32031\,
            I => \N__32028\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__32028\,
            I => \N__32025\
        );

    \I__7678\ : Odrv4
    port map (
            O => \N__32025\,
            I => \this_ppu.un1_M_vaddress_q_3_5\
        );

    \I__7677\ : InMux
    port map (
            O => \N__32022\,
            I => \N__32019\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__32019\,
            I => \N__32016\
        );

    \I__7675\ : Span4Mux_h
    port map (
            O => \N__32016\,
            I => \N__32013\
        );

    \I__7674\ : Span4Mux_h
    port map (
            O => \N__32013\,
            I => \N__32010\
        );

    \I__7673\ : Odrv4
    port map (
            O => \N__32010\,
            I => \M_this_data_tmp_qZ0Z_5\
        );

    \I__7672\ : InMux
    port map (
            O => \N__32007\,
            I => \N__32004\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__32004\,
            I => \M_this_oam_ram_write_data_5\
        );

    \I__7670\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31997\
        );

    \I__7669\ : CascadeMux
    port map (
            O => \N__32000\,
            I => \N__31994\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__31997\,
            I => \N__31991\
        );

    \I__7667\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31988\
        );

    \I__7666\ : Span4Mux_h
    port map (
            O => \N__31991\,
            I => \N__31985\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__31988\,
            I => \N__31981\
        );

    \I__7664\ : Span4Mux_h
    port map (
            O => \N__31985\,
            I => \N__31978\
        );

    \I__7663\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31975\
        );

    \I__7662\ : Odrv12
    port map (
            O => \N__31981\,
            I => \M_this_oam_ram_read_data_9\
        );

    \I__7661\ : Odrv4
    port map (
            O => \N__31978\,
            I => \M_this_oam_ram_read_data_9\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__31975\,
            I => \M_this_oam_ram_read_data_9\
        );

    \I__7659\ : InMux
    port map (
            O => \N__31968\,
            I => \N__31965\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__31965\,
            I => \M_this_oam_ram_write_data_9\
        );

    \I__7657\ : InMux
    port map (
            O => \N__31962\,
            I => \N__31959\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__31959\,
            I => \M_this_oam_ram_write_data_18\
        );

    \I__7655\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31953\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__31953\,
            I => \M_this_oam_ram_write_data_20\
        );

    \I__7653\ : InMux
    port map (
            O => \N__31950\,
            I => \N__31947\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__31947\,
            I => \M_this_oam_ram_write_data_29\
        );

    \I__7651\ : InMux
    port map (
            O => \N__31944\,
            I => \N__31941\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__31941\,
            I => \M_this_oam_ram_write_data_30\
        );

    \I__7649\ : InMux
    port map (
            O => \N__31938\,
            I => \N__31935\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__31935\,
            I => \N__31932\
        );

    \I__7647\ : Odrv4
    port map (
            O => \N__31932\,
            I => \M_this_external_address_q_3_0_12\
        );

    \I__7646\ : CEMux
    port map (
            O => \N__31929\,
            I => \N__31926\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__31926\,
            I => \N__31922\
        );

    \I__7644\ : CEMux
    port map (
            O => \N__31925\,
            I => \N__31919\
        );

    \I__7643\ : Span4Mux_h
    port map (
            O => \N__31922\,
            I => \N__31916\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__31919\,
            I => \N__31913\
        );

    \I__7641\ : Span4Mux_h
    port map (
            O => \N__31916\,
            I => \N__31910\
        );

    \I__7640\ : Span4Mux_h
    port map (
            O => \N__31913\,
            I => \N__31907\
        );

    \I__7639\ : Odrv4
    port map (
            O => \N__31910\,
            I => \this_sprites_ram.mem_WE_4\
        );

    \I__7638\ : Odrv4
    port map (
            O => \N__31907\,
            I => \this_sprites_ram.mem_WE_4\
        );

    \I__7637\ : InMux
    port map (
            O => \N__31902\,
            I => \N__31899\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__31899\,
            I => \N__31896\
        );

    \I__7635\ : Span4Mux_h
    port map (
            O => \N__31896\,
            I => \N__31893\
        );

    \I__7634\ : Span4Mux_h
    port map (
            O => \N__31893\,
            I => \N__31890\
        );

    \I__7633\ : Odrv4
    port map (
            O => \N__31890\,
            I => \this_ppu.un1_M_haddress_q_2_5\
        );

    \I__7632\ : InMux
    port map (
            O => \N__31887\,
            I => \N__31884\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__31884\,
            I => \M_this_oam_ram_write_data_13\
        );

    \I__7630\ : InMux
    port map (
            O => \N__31881\,
            I => \N__31878\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__31878\,
            I => \M_this_oam_ram_write_data_15\
        );

    \I__7628\ : InMux
    port map (
            O => \N__31875\,
            I => \N__31872\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__31872\,
            I => \N__31868\
        );

    \I__7626\ : CascadeMux
    port map (
            O => \N__31871\,
            I => \N__31865\
        );

    \I__7625\ : Span4Mux_h
    port map (
            O => \N__31868\,
            I => \N__31862\
        );

    \I__7624\ : InMux
    port map (
            O => \N__31865\,
            I => \N__31859\
        );

    \I__7623\ : Odrv4
    port map (
            O => \N__31862\,
            I => \M_this_oam_ram_read_data_15\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__31859\,
            I => \M_this_oam_ram_read_data_15\
        );

    \I__7621\ : InMux
    port map (
            O => \N__31854\,
            I => \N__31851\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__31851\,
            I => \N__31848\
        );

    \I__7619\ : Span4Mux_h
    port map (
            O => \N__31848\,
            I => \N__31845\
        );

    \I__7618\ : Span4Mux_h
    port map (
            O => \N__31845\,
            I => \N__31842\
        );

    \I__7617\ : Odrv4
    port map (
            O => \N__31842\,
            I => \this_ppu.un1_M_haddress_q_2_7\
        );

    \I__7616\ : InMux
    port map (
            O => \N__31839\,
            I => \N__31835\
        );

    \I__7615\ : InMux
    port map (
            O => \N__31838\,
            I => \N__31832\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__31835\,
            I => \N__31825\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__31832\,
            I => \N__31825\
        );

    \I__7612\ : InMux
    port map (
            O => \N__31831\,
            I => \N__31820\
        );

    \I__7611\ : InMux
    port map (
            O => \N__31830\,
            I => \N__31820\
        );

    \I__7610\ : Odrv12
    port map (
            O => \N__31825\,
            I => \M_this_oam_ram_read_data_12\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__31820\,
            I => \M_this_oam_ram_read_data_12\
        );

    \I__7608\ : InMux
    port map (
            O => \N__31815\,
            I => \N__31812\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__31812\,
            I => \N__31807\
        );

    \I__7606\ : InMux
    port map (
            O => \N__31811\,
            I => \N__31804\
        );

    \I__7605\ : InMux
    port map (
            O => \N__31810\,
            I => \N__31801\
        );

    \I__7604\ : Span4Mux_h
    port map (
            O => \N__31807\,
            I => \N__31798\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__31804\,
            I => \N__31791\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__31801\,
            I => \N__31791\
        );

    \I__7601\ : Span4Mux_h
    port map (
            O => \N__31798\,
            I => \N__31788\
        );

    \I__7600\ : InMux
    port map (
            O => \N__31797\,
            I => \N__31783\
        );

    \I__7599\ : InMux
    port map (
            O => \N__31796\,
            I => \N__31783\
        );

    \I__7598\ : Odrv12
    port map (
            O => \N__31791\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__7597\ : Odrv4
    port map (
            O => \N__31788\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__31783\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__7595\ : InMux
    port map (
            O => \N__31776\,
            I => \N__31773\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__31773\,
            I => \this_ppu.un1_oam_data_1_c2\
        );

    \I__7593\ : InMux
    port map (
            O => \N__31770\,
            I => \N__31767\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__31767\,
            I => \N__31764\
        );

    \I__7591\ : Span4Mux_h
    port map (
            O => \N__31764\,
            I => \N__31759\
        );

    \I__7590\ : InMux
    port map (
            O => \N__31763\,
            I => \N__31756\
        );

    \I__7589\ : InMux
    port map (
            O => \N__31762\,
            I => \N__31753\
        );

    \I__7588\ : Odrv4
    port map (
            O => \N__31759\,
            I => \M_this_oam_ram_read_data_14\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__31756\,
            I => \M_this_oam_ram_read_data_14\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__31753\,
            I => \M_this_oam_ram_read_data_14\
        );

    \I__7585\ : CascadeMux
    port map (
            O => \N__31746\,
            I => \this_ppu.un1_oam_data_1_c2_cascade_\
        );

    \I__7584\ : InMux
    port map (
            O => \N__31743\,
            I => \N__31740\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__31740\,
            I => \N__31734\
        );

    \I__7582\ : InMux
    port map (
            O => \N__31739\,
            I => \N__31727\
        );

    \I__7581\ : InMux
    port map (
            O => \N__31738\,
            I => \N__31727\
        );

    \I__7580\ : InMux
    port map (
            O => \N__31737\,
            I => \N__31727\
        );

    \I__7579\ : Odrv12
    port map (
            O => \N__31734\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__31727\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__7577\ : InMux
    port map (
            O => \N__31722\,
            I => \N__31719\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__31719\,
            I => \N__31716\
        );

    \I__7575\ : Span4Mux_h
    port map (
            O => \N__31716\,
            I => \N__31713\
        );

    \I__7574\ : Span4Mux_h
    port map (
            O => \N__31713\,
            I => \N__31710\
        );

    \I__7573\ : Odrv4
    port map (
            O => \N__31710\,
            I => \this_ppu.un1_M_haddress_q_2_6\
        );

    \I__7572\ : InMux
    port map (
            O => \N__31707\,
            I => \N__31703\
        );

    \I__7571\ : InMux
    port map (
            O => \N__31706\,
            I => \N__31699\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__31703\,
            I => \N__31696\
        );

    \I__7569\ : InMux
    port map (
            O => \N__31702\,
            I => \N__31693\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__31699\,
            I => \N__31690\
        );

    \I__7567\ : Span4Mux_v
    port map (
            O => \N__31696\,
            I => \N__31685\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__31693\,
            I => \N__31685\
        );

    \I__7565\ : Span4Mux_v
    port map (
            O => \N__31690\,
            I => \N__31680\
        );

    \I__7564\ : Span4Mux_h
    port map (
            O => \N__31685\,
            I => \N__31680\
        );

    \I__7563\ : Odrv4
    port map (
            O => \N__31680\,
            I => \this_vga_signals.N_746\
        );

    \I__7562\ : InMux
    port map (
            O => \N__31677\,
            I => \N__31674\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__31674\,
            I => \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0Z0Z_12\
        );

    \I__7560\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31667\
        );

    \I__7559\ : InMux
    port map (
            O => \N__31670\,
            I => \N__31664\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__31667\,
            I => \N__31661\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__31664\,
            I => \M_this_oam_address_q_0_i_o3_0_a2_5\
        );

    \I__7556\ : Odrv4
    port map (
            O => \N__31661\,
            I => \M_this_oam_address_q_0_i_o3_0_a2_5\
        );

    \I__7555\ : CascadeMux
    port map (
            O => \N__31656\,
            I => \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0Z0Z_12_cascade_\
        );

    \I__7554\ : IoInMux
    port map (
            O => \N__31653\,
            I => \N__31650\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__31650\,
            I => \N__31647\
        );

    \I__7552\ : IoSpan4Mux
    port map (
            O => \N__31647\,
            I => \N__31643\
        );

    \I__7551\ : InMux
    port map (
            O => \N__31646\,
            I => \N__31640\
        );

    \I__7550\ : Span4Mux_s2_h
    port map (
            O => \N__31643\,
            I => \N__31635\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__31640\,
            I => \N__31632\
        );

    \I__7548\ : InMux
    port map (
            O => \N__31639\,
            I => \N__31629\
        );

    \I__7547\ : InMux
    port map (
            O => \N__31638\,
            I => \N__31626\
        );

    \I__7546\ : Sp12to4
    port map (
            O => \N__31635\,
            I => \N__31621\
        );

    \I__7545\ : Span4Mux_h
    port map (
            O => \N__31632\,
            I => \N__31618\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__31629\,
            I => \N__31615\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__31626\,
            I => \N__31612\
        );

    \I__7542\ : InMux
    port map (
            O => \N__31625\,
            I => \N__31609\
        );

    \I__7541\ : InMux
    port map (
            O => \N__31624\,
            I => \N__31606\
        );

    \I__7540\ : Span12Mux_s11_h
    port map (
            O => \N__31621\,
            I => \N__31603\
        );

    \I__7539\ : Span4Mux_v
    port map (
            O => \N__31618\,
            I => \N__31598\
        );

    \I__7538\ : Span4Mux_h
    port map (
            O => \N__31615\,
            I => \N__31598\
        );

    \I__7537\ : Span4Mux_v
    port map (
            O => \N__31612\,
            I => \N__31595\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__31609\,
            I => \N__31590\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__31606\,
            I => \N__31590\
        );

    \I__7534\ : Span12Mux_v
    port map (
            O => \N__31603\,
            I => \N__31586\
        );

    \I__7533\ : Span4Mux_h
    port map (
            O => \N__31598\,
            I => \N__31583\
        );

    \I__7532\ : Span4Mux_h
    port map (
            O => \N__31595\,
            I => \N__31578\
        );

    \I__7531\ : Span4Mux_v
    port map (
            O => \N__31590\,
            I => \N__31578\
        );

    \I__7530\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31575\
        );

    \I__7529\ : Odrv12
    port map (
            O => \N__31586\,
            I => led_c_1
        );

    \I__7528\ : Odrv4
    port map (
            O => \N__31583\,
            I => led_c_1
        );

    \I__7527\ : Odrv4
    port map (
            O => \N__31578\,
            I => led_c_1
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__31575\,
            I => led_c_1
        );

    \I__7525\ : InMux
    port map (
            O => \N__31566\,
            I => \N__31563\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__31563\,
            I => \N__31559\
        );

    \I__7523\ : InMux
    port map (
            O => \N__31562\,
            I => \N__31556\
        );

    \I__7522\ : Span4Mux_v
    port map (
            O => \N__31559\,
            I => \N__31550\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__31556\,
            I => \N__31550\
        );

    \I__7520\ : InMux
    port map (
            O => \N__31555\,
            I => \N__31547\
        );

    \I__7519\ : Span4Mux_h
    port map (
            O => \N__31550\,
            I => \N__31544\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__31547\,
            I => \M_this_substate_qZ0\
        );

    \I__7517\ : Odrv4
    port map (
            O => \N__31544\,
            I => \M_this_substate_qZ0\
        );

    \I__7516\ : InMux
    port map (
            O => \N__31539\,
            I => \N__31535\
        );

    \I__7515\ : InMux
    port map (
            O => \N__31538\,
            I => \N__31532\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__31535\,
            I => \N__31528\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__31532\,
            I => \N__31525\
        );

    \I__7512\ : InMux
    port map (
            O => \N__31531\,
            I => \N__31522\
        );

    \I__7511\ : Span4Mux_v
    port map (
            O => \N__31528\,
            I => \N__31519\
        );

    \I__7510\ : Span4Mux_v
    port map (
            O => \N__31525\,
            I => \N__31516\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__31522\,
            I => \N__31513\
        );

    \I__7508\ : Odrv4
    port map (
            O => \N__31519\,
            I => \this_vga_signals.N_419_0\
        );

    \I__7507\ : Odrv4
    port map (
            O => \N__31516\,
            I => \this_vga_signals.N_419_0\
        );

    \I__7506\ : Odrv12
    port map (
            O => \N__31513\,
            I => \this_vga_signals.N_419_0\
        );

    \I__7505\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31503\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__31503\,
            I => \N__31500\
        );

    \I__7503\ : Span4Mux_h
    port map (
            O => \N__31500\,
            I => \N__31497\
        );

    \I__7502\ : Odrv4
    port map (
            O => \N__31497\,
            I => \M_this_data_count_q_cry_6_THRU_CO\
        );

    \I__7501\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31476\
        );

    \I__7500\ : InMux
    port map (
            O => \N__31493\,
            I => \N__31465\
        );

    \I__7499\ : InMux
    port map (
            O => \N__31492\,
            I => \N__31465\
        );

    \I__7498\ : InMux
    port map (
            O => \N__31491\,
            I => \N__31465\
        );

    \I__7497\ : InMux
    port map (
            O => \N__31490\,
            I => \N__31465\
        );

    \I__7496\ : InMux
    port map (
            O => \N__31489\,
            I => \N__31465\
        );

    \I__7495\ : InMux
    port map (
            O => \N__31488\,
            I => \N__31458\
        );

    \I__7494\ : InMux
    port map (
            O => \N__31487\,
            I => \N__31458\
        );

    \I__7493\ : InMux
    port map (
            O => \N__31486\,
            I => \N__31458\
        );

    \I__7492\ : InMux
    port map (
            O => \N__31485\,
            I => \N__31451\
        );

    \I__7491\ : InMux
    port map (
            O => \N__31484\,
            I => \N__31451\
        );

    \I__7490\ : InMux
    port map (
            O => \N__31483\,
            I => \N__31451\
        );

    \I__7489\ : InMux
    port map (
            O => \N__31482\,
            I => \N__31442\
        );

    \I__7488\ : InMux
    port map (
            O => \N__31481\,
            I => \N__31442\
        );

    \I__7487\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31442\
        );

    \I__7486\ : InMux
    port map (
            O => \N__31479\,
            I => \N__31442\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__31476\,
            I => \N_716_i\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__31465\,
            I => \N_716_i\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__31458\,
            I => \N_716_i\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__31451\,
            I => \N_716_i\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__31442\,
            I => \N_716_i\
        );

    \I__7480\ : CascadeMux
    port map (
            O => \N__31431\,
            I => \N__31428\
        );

    \I__7479\ : InMux
    port map (
            O => \N__31428\,
            I => \N__31424\
        );

    \I__7478\ : CascadeMux
    port map (
            O => \N__31427\,
            I => \N__31421\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__31424\,
            I => \N__31417\
        );

    \I__7476\ : InMux
    port map (
            O => \N__31421\,
            I => \N__31414\
        );

    \I__7475\ : InMux
    port map (
            O => \N__31420\,
            I => \N__31411\
        );

    \I__7474\ : Span4Mux_v
    port map (
            O => \N__31417\,
            I => \N__31406\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__31414\,
            I => \N__31406\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__31411\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__7471\ : Odrv4
    port map (
            O => \N__31406\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__7470\ : CEMux
    port map (
            O => \N__31401\,
            I => \N__31397\
        );

    \I__7469\ : CEMux
    port map (
            O => \N__31400\,
            I => \N__31394\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__31397\,
            I => \N__31389\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__31394\,
            I => \N__31386\
        );

    \I__7466\ : CEMux
    port map (
            O => \N__31393\,
            I => \N__31383\
        );

    \I__7465\ : CEMux
    port map (
            O => \N__31392\,
            I => \N__31380\
        );

    \I__7464\ : Span4Mux_v
    port map (
            O => \N__31389\,
            I => \N__31377\
        );

    \I__7463\ : Span4Mux_v
    port map (
            O => \N__31386\,
            I => \N__31374\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__31383\,
            I => \N__31369\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__31380\,
            I => \N__31369\
        );

    \I__7460\ : Odrv4
    port map (
            O => \N__31377\,
            I => \N_364\
        );

    \I__7459\ : Odrv4
    port map (
            O => \N__31374\,
            I => \N_364\
        );

    \I__7458\ : Odrv4
    port map (
            O => \N__31369\,
            I => \N_364\
        );

    \I__7457\ : CascadeMux
    port map (
            O => \N__31362\,
            I => \N__31357\
        );

    \I__7456\ : InMux
    port map (
            O => \N__31361\,
            I => \N__31352\
        );

    \I__7455\ : CascadeMux
    port map (
            O => \N__31360\,
            I => \N__31347\
        );

    \I__7454\ : InMux
    port map (
            O => \N__31357\,
            I => \N__31344\
        );

    \I__7453\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31341\
        );

    \I__7452\ : CascadeMux
    port map (
            O => \N__31355\,
            I => \N__31338\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__31352\,
            I => \N__31334\
        );

    \I__7450\ : InMux
    port map (
            O => \N__31351\,
            I => \N__31331\
        );

    \I__7449\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31328\
        );

    \I__7448\ : InMux
    port map (
            O => \N__31347\,
            I => \N__31325\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__31344\,
            I => \N__31321\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__31341\,
            I => \N__31318\
        );

    \I__7445\ : InMux
    port map (
            O => \N__31338\,
            I => \N__31315\
        );

    \I__7444\ : CascadeMux
    port map (
            O => \N__31337\,
            I => \N__31312\
        );

    \I__7443\ : Span4Mux_v
    port map (
            O => \N__31334\,
            I => \N__31307\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__31331\,
            I => \N__31307\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__31328\,
            I => \N__31304\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__31325\,
            I => \N__31300\
        );

    \I__7439\ : InMux
    port map (
            O => \N__31324\,
            I => \N__31297\
        );

    \I__7438\ : Span4Mux_v
    port map (
            O => \N__31321\,
            I => \N__31292\
        );

    \I__7437\ : Span4Mux_v
    port map (
            O => \N__31318\,
            I => \N__31292\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__31315\,
            I => \N__31289\
        );

    \I__7435\ : InMux
    port map (
            O => \N__31312\,
            I => \N__31286\
        );

    \I__7434\ : Span4Mux_v
    port map (
            O => \N__31307\,
            I => \N__31283\
        );

    \I__7433\ : Span4Mux_v
    port map (
            O => \N__31304\,
            I => \N__31280\
        );

    \I__7432\ : InMux
    port map (
            O => \N__31303\,
            I => \N__31277\
        );

    \I__7431\ : Span4Mux_v
    port map (
            O => \N__31300\,
            I => \N__31274\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__31297\,
            I => \N__31271\
        );

    \I__7429\ : Span4Mux_h
    port map (
            O => \N__31292\,
            I => \N__31264\
        );

    \I__7428\ : Span4Mux_v
    port map (
            O => \N__31289\,
            I => \N__31264\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__31286\,
            I => \N__31264\
        );

    \I__7426\ : Sp12to4
    port map (
            O => \N__31283\,
            I => \N__31256\
        );

    \I__7425\ : Sp12to4
    port map (
            O => \N__31280\,
            I => \N__31256\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__31277\,
            I => \N__31256\
        );

    \I__7423\ : Span4Mux_v
    port map (
            O => \N__31274\,
            I => \N__31253\
        );

    \I__7422\ : Span4Mux_v
    port map (
            O => \N__31271\,
            I => \N__31250\
        );

    \I__7421\ : Span4Mux_h
    port map (
            O => \N__31264\,
            I => \N__31247\
        );

    \I__7420\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31244\
        );

    \I__7419\ : Span12Mux_h
    port map (
            O => \N__31256\,
            I => \N__31241\
        );

    \I__7418\ : Sp12to4
    port map (
            O => \N__31253\,
            I => \N__31236\
        );

    \I__7417\ : Sp12to4
    port map (
            O => \N__31250\,
            I => \N__31236\
        );

    \I__7416\ : Span4Mux_v
    port map (
            O => \N__31247\,
            I => \N__31231\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__31244\,
            I => \N__31231\
        );

    \I__7414\ : Span12Mux_v
    port map (
            O => \N__31241\,
            I => \N__31228\
        );

    \I__7413\ : Span12Mux_h
    port map (
            O => \N__31236\,
            I => \N__31225\
        );

    \I__7412\ : Span4Mux_v
    port map (
            O => \N__31231\,
            I => \N__31222\
        );

    \I__7411\ : Odrv12
    port map (
            O => \N__31228\,
            I => port_data_c_0
        );

    \I__7410\ : Odrv12
    port map (
            O => \N__31225\,
            I => port_data_c_0
        );

    \I__7409\ : Odrv4
    port map (
            O => \N__31222\,
            I => port_data_c_0
        );

    \I__7408\ : CascadeMux
    port map (
            O => \N__31215\,
            I => \N__31210\
        );

    \I__7407\ : InMux
    port map (
            O => \N__31214\,
            I => \N__31206\
        );

    \I__7406\ : InMux
    port map (
            O => \N__31213\,
            I => \N__31202\
        );

    \I__7405\ : InMux
    port map (
            O => \N__31210\,
            I => \N__31197\
        );

    \I__7404\ : InMux
    port map (
            O => \N__31209\,
            I => \N__31197\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__31206\,
            I => \N__31194\
        );

    \I__7402\ : InMux
    port map (
            O => \N__31205\,
            I => \N__31191\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__31202\,
            I => \N__31188\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__31197\,
            I => \N__31185\
        );

    \I__7399\ : Span4Mux_v
    port map (
            O => \N__31194\,
            I => \N__31179\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__31191\,
            I => \N__31179\
        );

    \I__7397\ : Span4Mux_v
    port map (
            O => \N__31188\,
            I => \N__31173\
        );

    \I__7396\ : Span4Mux_v
    port map (
            O => \N__31185\,
            I => \N__31173\
        );

    \I__7395\ : InMux
    port map (
            O => \N__31184\,
            I => \N__31170\
        );

    \I__7394\ : Span4Mux_h
    port map (
            O => \N__31179\,
            I => \N__31167\
        );

    \I__7393\ : InMux
    port map (
            O => \N__31178\,
            I => \N__31164\
        );

    \I__7392\ : Sp12to4
    port map (
            O => \N__31173\,
            I => \N__31159\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__31170\,
            I => \N__31159\
        );

    \I__7390\ : Span4Mux_v
    port map (
            O => \N__31167\,
            I => \N__31156\
        );

    \I__7389\ : LocalMux
    port map (
            O => \N__31164\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__7388\ : Odrv12
    port map (
            O => \N__31159\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__7387\ : Odrv4
    port map (
            O => \N__31156\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__7386\ : InMux
    port map (
            O => \N__31149\,
            I => \N__31137\
        );

    \I__7385\ : InMux
    port map (
            O => \N__31148\,
            I => \N__31137\
        );

    \I__7384\ : InMux
    port map (
            O => \N__31147\,
            I => \N__31134\
        );

    \I__7383\ : InMux
    port map (
            O => \N__31146\,
            I => \N__31131\
        );

    \I__7382\ : CascadeMux
    port map (
            O => \N__31145\,
            I => \N__31128\
        );

    \I__7381\ : InMux
    port map (
            O => \N__31144\,
            I => \N__31112\
        );

    \I__7380\ : CascadeMux
    port map (
            O => \N__31143\,
            I => \N__31108\
        );

    \I__7379\ : CascadeMux
    port map (
            O => \N__31142\,
            I => \N__31098\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__31137\,
            I => \N__31090\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__31134\,
            I => \N__31090\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__31131\,
            I => \N__31090\
        );

    \I__7375\ : InMux
    port map (
            O => \N__31128\,
            I => \N__31085\
        );

    \I__7374\ : InMux
    port map (
            O => \N__31127\,
            I => \N__31085\
        );

    \I__7373\ : InMux
    port map (
            O => \N__31126\,
            I => \N__31077\
        );

    \I__7372\ : InMux
    port map (
            O => \N__31125\,
            I => \N__31077\
        );

    \I__7371\ : InMux
    port map (
            O => \N__31124\,
            I => \N__31073\
        );

    \I__7370\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31068\
        );

    \I__7369\ : InMux
    port map (
            O => \N__31122\,
            I => \N__31068\
        );

    \I__7368\ : InMux
    port map (
            O => \N__31121\,
            I => \N__31063\
        );

    \I__7367\ : InMux
    port map (
            O => \N__31120\,
            I => \N__31063\
        );

    \I__7366\ : InMux
    port map (
            O => \N__31119\,
            I => \N__31060\
        );

    \I__7365\ : InMux
    port map (
            O => \N__31118\,
            I => \N__31057\
        );

    \I__7364\ : InMux
    port map (
            O => \N__31117\,
            I => \N__31054\
        );

    \I__7363\ : InMux
    port map (
            O => \N__31116\,
            I => \N__31049\
        );

    \I__7362\ : InMux
    port map (
            O => \N__31115\,
            I => \N__31049\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__31112\,
            I => \N__31046\
        );

    \I__7360\ : InMux
    port map (
            O => \N__31111\,
            I => \N__31041\
        );

    \I__7359\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31041\
        );

    \I__7358\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31038\
        );

    \I__7357\ : InMux
    port map (
            O => \N__31106\,
            I => \N__31035\
        );

    \I__7356\ : InMux
    port map (
            O => \N__31105\,
            I => \N__31030\
        );

    \I__7355\ : InMux
    port map (
            O => \N__31104\,
            I => \N__31030\
        );

    \I__7354\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31027\
        );

    \I__7353\ : InMux
    port map (
            O => \N__31102\,
            I => \N__31024\
        );

    \I__7352\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31017\
        );

    \I__7351\ : InMux
    port map (
            O => \N__31098\,
            I => \N__31017\
        );

    \I__7350\ : InMux
    port map (
            O => \N__31097\,
            I => \N__31017\
        );

    \I__7349\ : Span4Mux_v
    port map (
            O => \N__31090\,
            I => \N__31014\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__31085\,
            I => \N__31011\
        );

    \I__7347\ : InMux
    port map (
            O => \N__31084\,
            I => \N__31004\
        );

    \I__7346\ : InMux
    port map (
            O => \N__31083\,
            I => \N__31004\
        );

    \I__7345\ : InMux
    port map (
            O => \N__31082\,
            I => \N__31004\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__31077\,
            I => \N__30997\
        );

    \I__7343\ : InMux
    port map (
            O => \N__31076\,
            I => \N__30994\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__31073\,
            I => \N__30987\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__31068\,
            I => \N__30987\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__31063\,
            I => \N__30987\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__31060\,
            I => \N__30982\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__31057\,
            I => \N__30982\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__31054\,
            I => \N__30973\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__31049\,
            I => \N__30973\
        );

    \I__7335\ : Span4Mux_v
    port map (
            O => \N__31046\,
            I => \N__30973\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__31041\,
            I => \N__30973\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__31038\,
            I => \N__30970\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__31035\,
            I => \N__30967\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__31030\,
            I => \N__30963\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__31027\,
            I => \N__30960\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__31024\,
            I => \N__30949\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__31017\,
            I => \N__30949\
        );

    \I__7327\ : Span4Mux_h
    port map (
            O => \N__31014\,
            I => \N__30949\
        );

    \I__7326\ : Span4Mux_h
    port map (
            O => \N__31011\,
            I => \N__30949\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__31004\,
            I => \N__30949\
        );

    \I__7324\ : InMux
    port map (
            O => \N__31003\,
            I => \N__30940\
        );

    \I__7323\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30935\
        );

    \I__7322\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30935\
        );

    \I__7321\ : InMux
    port map (
            O => \N__31000\,
            I => \N__30932\
        );

    \I__7320\ : Span4Mux_h
    port map (
            O => \N__30997\,
            I => \N__30923\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__30994\,
            I => \N__30923\
        );

    \I__7318\ : Span4Mux_v
    port map (
            O => \N__30987\,
            I => \N__30923\
        );

    \I__7317\ : Span4Mux_v
    port map (
            O => \N__30982\,
            I => \N__30923\
        );

    \I__7316\ : Span4Mux_h
    port map (
            O => \N__30973\,
            I => \N__30918\
        );

    \I__7315\ : Span4Mux_h
    port map (
            O => \N__30970\,
            I => \N__30918\
        );

    \I__7314\ : Span4Mux_h
    port map (
            O => \N__30967\,
            I => \N__30915\
        );

    \I__7313\ : InMux
    port map (
            O => \N__30966\,
            I => \N__30912\
        );

    \I__7312\ : Span4Mux_v
    port map (
            O => \N__30963\,
            I => \N__30905\
        );

    \I__7311\ : Span4Mux_h
    port map (
            O => \N__30960\,
            I => \N__30905\
        );

    \I__7310\ : Span4Mux_v
    port map (
            O => \N__30949\,
            I => \N__30905\
        );

    \I__7309\ : InMux
    port map (
            O => \N__30948\,
            I => \N__30898\
        );

    \I__7308\ : InMux
    port map (
            O => \N__30947\,
            I => \N__30898\
        );

    \I__7307\ : InMux
    port map (
            O => \N__30946\,
            I => \N__30898\
        );

    \I__7306\ : InMux
    port map (
            O => \N__30945\,
            I => \N__30891\
        );

    \I__7305\ : InMux
    port map (
            O => \N__30944\,
            I => \N__30891\
        );

    \I__7304\ : InMux
    port map (
            O => \N__30943\,
            I => \N__30891\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__30940\,
            I => \N_888_0\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__30935\,
            I => \N_888_0\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__30932\,
            I => \N_888_0\
        );

    \I__7300\ : Odrv4
    port map (
            O => \N__30923\,
            I => \N_888_0\
        );

    \I__7299\ : Odrv4
    port map (
            O => \N__30918\,
            I => \N_888_0\
        );

    \I__7298\ : Odrv4
    port map (
            O => \N__30915\,
            I => \N_888_0\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__30912\,
            I => \N_888_0\
        );

    \I__7296\ : Odrv4
    port map (
            O => \N__30905\,
            I => \N_888_0\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__30898\,
            I => \N_888_0\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__30891\,
            I => \N_888_0\
        );

    \I__7293\ : CascadeMux
    port map (
            O => \N__30870\,
            I => \N_760_cascade_\
        );

    \I__7292\ : InMux
    port map (
            O => \N__30867\,
            I => \N__30864\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__30864\,
            I => \N__30861\
        );

    \I__7290\ : Span4Mux_v
    port map (
            O => \N__30861\,
            I => \N__30858\
        );

    \I__7289\ : Odrv4
    port map (
            O => \N__30858\,
            I => \M_this_data_tmp_qZ0Z_8\
        );

    \I__7288\ : CascadeMux
    port map (
            O => \N__30855\,
            I => \N__30849\
        );

    \I__7287\ : CascadeMux
    port map (
            O => \N__30854\,
            I => \N__30846\
        );

    \I__7286\ : CascadeMux
    port map (
            O => \N__30853\,
            I => \N__30841\
        );

    \I__7285\ : CascadeMux
    port map (
            O => \N__30852\,
            I => \N__30838\
        );

    \I__7284\ : InMux
    port map (
            O => \N__30849\,
            I => \N__30835\
        );

    \I__7283\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30832\
        );

    \I__7282\ : CascadeMux
    port map (
            O => \N__30845\,
            I => \N__30829\
        );

    \I__7281\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30826\
        );

    \I__7280\ : InMux
    port map (
            O => \N__30841\,
            I => \N__30823\
        );

    \I__7279\ : InMux
    port map (
            O => \N__30838\,
            I => \N__30820\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__30835\,
            I => \N__30815\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__30832\,
            I => \N__30815\
        );

    \I__7276\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30812\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__30826\,
            I => \N__30808\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__30823\,
            I => \N__30805\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__30820\,
            I => \N__30802\
        );

    \I__7272\ : Span4Mux_v
    port map (
            O => \N__30815\,
            I => \N__30797\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__30812\,
            I => \N__30797\
        );

    \I__7270\ : InMux
    port map (
            O => \N__30811\,
            I => \N__30794\
        );

    \I__7269\ : Span4Mux_v
    port map (
            O => \N__30808\,
            I => \N__30787\
        );

    \I__7268\ : Span4Mux_v
    port map (
            O => \N__30805\,
            I => \N__30787\
        );

    \I__7267\ : Span4Mux_h
    port map (
            O => \N__30802\,
            I => \N__30787\
        );

    \I__7266\ : Sp12to4
    port map (
            O => \N__30797\,
            I => \N__30782\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__30794\,
            I => \N__30782\
        );

    \I__7264\ : Span4Mux_v
    port map (
            O => \N__30787\,
            I => \N__30779\
        );

    \I__7263\ : Span12Mux_v
    port map (
            O => \N__30782\,
            I => \N__30776\
        );

    \I__7262\ : Odrv4
    port map (
            O => \N__30779\,
            I => \N_413_0\
        );

    \I__7261\ : Odrv12
    port map (
            O => \N__30776\,
            I => \N_413_0\
        );

    \I__7260\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30765\
        );

    \I__7259\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30765\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__30765\,
            I => \N__30761\
        );

    \I__7257\ : InMux
    port map (
            O => \N__30764\,
            I => \N__30758\
        );

    \I__7256\ : Span4Mux_v
    port map (
            O => \N__30761\,
            I => \N__30755\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__30758\,
            I => \N__30752\
        );

    \I__7254\ : Odrv4
    port map (
            O => \N__30755\,
            I => \un1_M_this_oam_address_q_c4\
        );

    \I__7253\ : Odrv12
    port map (
            O => \N__30752\,
            I => \un1_M_this_oam_address_q_c4\
        );

    \I__7252\ : CascadeMux
    port map (
            O => \N__30747\,
            I => \N__30744\
        );

    \I__7251\ : CascadeBuf
    port map (
            O => \N__30744\,
            I => \N__30741\
        );

    \I__7250\ : CascadeMux
    port map (
            O => \N__30741\,
            I => \N__30738\
        );

    \I__7249\ : InMux
    port map (
            O => \N__30738\,
            I => \N__30735\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__30735\,
            I => \N__30732\
        );

    \I__7247\ : Span4Mux_h
    port map (
            O => \N__30732\,
            I => \N__30729\
        );

    \I__7246\ : Span4Mux_v
    port map (
            O => \N__30729\,
            I => \N__30724\
        );

    \I__7245\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30721\
        );

    \I__7244\ : InMux
    port map (
            O => \N__30727\,
            I => \N__30718\
        );

    \I__7243\ : Span4Mux_h
    port map (
            O => \N__30724\,
            I => \N__30715\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__30721\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__30718\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__7240\ : Odrv4
    port map (
            O => \N__30715\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__7239\ : CascadeMux
    port map (
            O => \N__30708\,
            I => \N__30705\
        );

    \I__7238\ : CascadeBuf
    port map (
            O => \N__30705\,
            I => \N__30702\
        );

    \I__7237\ : CascadeMux
    port map (
            O => \N__30702\,
            I => \N__30699\
        );

    \I__7236\ : InMux
    port map (
            O => \N__30699\,
            I => \N__30696\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__30696\,
            I => \N__30693\
        );

    \I__7234\ : Span4Mux_h
    port map (
            O => \N__30693\,
            I => \N__30687\
        );

    \I__7233\ : InMux
    port map (
            O => \N__30692\,
            I => \N__30682\
        );

    \I__7232\ : InMux
    port map (
            O => \N__30691\,
            I => \N__30682\
        );

    \I__7231\ : InMux
    port map (
            O => \N__30690\,
            I => \N__30679\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__30687\,
            I => \N__30676\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__30682\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__30679\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__7227\ : Odrv4
    port map (
            O => \N__30676\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__7226\ : InMux
    port map (
            O => \N__30669\,
            I => \N__30662\
        );

    \I__7225\ : InMux
    port map (
            O => \N__30668\,
            I => \N__30659\
        );

    \I__7224\ : InMux
    port map (
            O => \N__30667\,
            I => \N__30655\
        );

    \I__7223\ : InMux
    port map (
            O => \N__30666\,
            I => \N__30652\
        );

    \I__7222\ : InMux
    port map (
            O => \N__30665\,
            I => \N__30649\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__30662\,
            I => \N__30645\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__30659\,
            I => \N__30642\
        );

    \I__7219\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30639\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__30655\,
            I => \N__30636\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__30652\,
            I => \N__30631\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__30649\,
            I => \N__30631\
        );

    \I__7215\ : InMux
    port map (
            O => \N__30648\,
            I => \N__30628\
        );

    \I__7214\ : Span4Mux_h
    port map (
            O => \N__30645\,
            I => \N__30625\
        );

    \I__7213\ : Span4Mux_h
    port map (
            O => \N__30642\,
            I => \N__30620\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__30639\,
            I => \N__30620\
        );

    \I__7211\ : Span4Mux_h
    port map (
            O => \N__30636\,
            I => \N__30615\
        );

    \I__7210\ : Span4Mux_h
    port map (
            O => \N__30631\,
            I => \N__30615\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__30628\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__7208\ : Odrv4
    port map (
            O => \N__30625\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__30620\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__7206\ : Odrv4
    port map (
            O => \N__30615\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__7205\ : InMux
    port map (
            O => \N__30606\,
            I => \N__30601\
        );

    \I__7204\ : CascadeMux
    port map (
            O => \N__30605\,
            I => \N__30598\
        );

    \I__7203\ : InMux
    port map (
            O => \N__30604\,
            I => \N__30594\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__30601\,
            I => \N__30590\
        );

    \I__7201\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30587\
        );

    \I__7200\ : InMux
    port map (
            O => \N__30597\,
            I => \N__30583\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__30594\,
            I => \N__30580\
        );

    \I__7198\ : InMux
    port map (
            O => \N__30593\,
            I => \N__30577\
        );

    \I__7197\ : Span4Mux_h
    port map (
            O => \N__30590\,
            I => \N__30572\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__30587\,
            I => \N__30572\
        );

    \I__7195\ : InMux
    port map (
            O => \N__30586\,
            I => \N__30569\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__30583\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__7193\ : Odrv4
    port map (
            O => \N__30580\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__30577\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__7191\ : Odrv4
    port map (
            O => \N__30572\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__30569\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__7189\ : InMux
    port map (
            O => \N__30558\,
            I => \N__30553\
        );

    \I__7188\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30549\
        );

    \I__7187\ : InMux
    port map (
            O => \N__30556\,
            I => \N__30544\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__30553\,
            I => \N__30541\
        );

    \I__7185\ : InMux
    port map (
            O => \N__30552\,
            I => \N__30538\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__30549\,
            I => \N__30535\
        );

    \I__7183\ : CascadeMux
    port map (
            O => \N__30548\,
            I => \N__30532\
        );

    \I__7182\ : InMux
    port map (
            O => \N__30547\,
            I => \N__30529\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__30544\,
            I => \N__30526\
        );

    \I__7180\ : Span4Mux_v
    port map (
            O => \N__30541\,
            I => \N__30519\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__30538\,
            I => \N__30519\
        );

    \I__7178\ : Span4Mux_h
    port map (
            O => \N__30535\,
            I => \N__30519\
        );

    \I__7177\ : InMux
    port map (
            O => \N__30532\,
            I => \N__30516\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__30529\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__7175\ : Odrv12
    port map (
            O => \N__30526\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__7174\ : Odrv4
    port map (
            O => \N__30519\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__30516\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__7172\ : InMux
    port map (
            O => \N__30507\,
            I => \N__30500\
        );

    \I__7171\ : InMux
    port map (
            O => \N__30506\,
            I => \N__30500\
        );

    \I__7170\ : InMux
    port map (
            O => \N__30505\,
            I => \N__30497\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__30500\,
            I => \N__30492\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__30497\,
            I => \N__30492\
        );

    \I__7167\ : Odrv4
    port map (
            O => \N__30492\,
            I => \un1_M_this_oam_address_q_c2\
        );

    \I__7166\ : InMux
    port map (
            O => \N__30489\,
            I => \N__30485\
        );

    \I__7165\ : InMux
    port map (
            O => \N__30488\,
            I => \N__30482\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__30485\,
            I => \N__30477\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__30482\,
            I => \N__30474\
        );

    \I__7162\ : InMux
    port map (
            O => \N__30481\,
            I => \N__30471\
        );

    \I__7161\ : InMux
    port map (
            O => \N__30480\,
            I => \N__30468\
        );

    \I__7160\ : Odrv4
    port map (
            O => \N__30477\,
            I => \this_vga_signals.N_461_0\
        );

    \I__7159\ : Odrv4
    port map (
            O => \N__30474\,
            I => \this_vga_signals.N_461_0\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__30471\,
            I => \this_vga_signals.N_461_0\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__30468\,
            I => \this_vga_signals.N_461_0\
        );

    \I__7156\ : CascadeMux
    port map (
            O => \N__30459\,
            I => \N__30456\
        );

    \I__7155\ : InMux
    port map (
            O => \N__30456\,
            I => \N__30453\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__30453\,
            I => \N__30450\
        );

    \I__7153\ : Span4Mux_h
    port map (
            O => \N__30450\,
            I => \N__30447\
        );

    \I__7152\ : Odrv4
    port map (
            O => \N__30447\,
            I => \this_vga_signals.N_747\
        );

    \I__7151\ : InMux
    port map (
            O => \N__30444\,
            I => \N__30439\
        );

    \I__7150\ : InMux
    port map (
            O => \N__30443\,
            I => \N__30435\
        );

    \I__7149\ : CascadeMux
    port map (
            O => \N__30442\,
            I => \N__30432\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__30439\,
            I => \N__30428\
        );

    \I__7147\ : InMux
    port map (
            O => \N__30438\,
            I => \N__30425\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__30435\,
            I => \N__30422\
        );

    \I__7145\ : InMux
    port map (
            O => \N__30432\,
            I => \N__30417\
        );

    \I__7144\ : InMux
    port map (
            O => \N__30431\,
            I => \N__30417\
        );

    \I__7143\ : Span4Mux_v
    port map (
            O => \N__30428\,
            I => \N__30411\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__30425\,
            I => \N__30411\
        );

    \I__7141\ : Span4Mux_v
    port map (
            O => \N__30422\,
            I => \N__30408\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__30417\,
            I => \N__30405\
        );

    \I__7139\ : CascadeMux
    port map (
            O => \N__30416\,
            I => \N__30401\
        );

    \I__7138\ : Span4Mux_h
    port map (
            O => \N__30411\,
            I => \N__30398\
        );

    \I__7137\ : Span4Mux_h
    port map (
            O => \N__30408\,
            I => \N__30393\
        );

    \I__7136\ : Span4Mux_v
    port map (
            O => \N__30405\,
            I => \N__30393\
        );

    \I__7135\ : InMux
    port map (
            O => \N__30404\,
            I => \N__30390\
        );

    \I__7134\ : InMux
    port map (
            O => \N__30401\,
            I => \N__30387\
        );

    \I__7133\ : Odrv4
    port map (
            O => \N__30398\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__7132\ : Odrv4
    port map (
            O => \N__30393\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__30390\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__30387\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__7129\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30371\
        );

    \I__7128\ : InMux
    port map (
            O => \N__30377\,
            I => \N__30368\
        );

    \I__7127\ : InMux
    port map (
            O => \N__30376\,
            I => \N__30365\
        );

    \I__7126\ : InMux
    port map (
            O => \N__30375\,
            I => \N__30362\
        );

    \I__7125\ : InMux
    port map (
            O => \N__30374\,
            I => \N__30358\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__30371\,
            I => \N__30355\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__30368\,
            I => \N__30352\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__30365\,
            I => \N__30347\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__30362\,
            I => \N__30347\
        );

    \I__7120\ : InMux
    port map (
            O => \N__30361\,
            I => \N__30344\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__30358\,
            I => \N__30339\
        );

    \I__7118\ : Span4Mux_v
    port map (
            O => \N__30355\,
            I => \N__30339\
        );

    \I__7117\ : Span4Mux_v
    port map (
            O => \N__30352\,
            I => \N__30332\
        );

    \I__7116\ : Span4Mux_v
    port map (
            O => \N__30347\,
            I => \N__30332\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__30344\,
            I => \N__30332\
        );

    \I__7114\ : Odrv4
    port map (
            O => \N__30339\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__7113\ : Odrv4
    port map (
            O => \N__30332\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__7112\ : InMux
    port map (
            O => \N__30327\,
            I => \N__30324\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__30324\,
            I => \N__30320\
        );

    \I__7110\ : InMux
    port map (
            O => \N__30323\,
            I => \N__30317\
        );

    \I__7109\ : Odrv4
    port map (
            O => \N__30320\,
            I => \this_vga_signals.N_433_0\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__30317\,
            I => \this_vga_signals.N_433_0\
        );

    \I__7107\ : InMux
    port map (
            O => \N__30312\,
            I => \N__30309\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__30309\,
            I => \N__30306\
        );

    \I__7105\ : Span4Mux_v
    port map (
            O => \N__30306\,
            I => \N__30303\
        );

    \I__7104\ : Odrv4
    port map (
            O => \N__30303\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_i_1Z0Z_0\
        );

    \I__7103\ : CascadeMux
    port map (
            O => \N__30300\,
            I => \N__30297\
        );

    \I__7102\ : InMux
    port map (
            O => \N__30297\,
            I => \N__30294\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__30294\,
            I => \N__30291\
        );

    \I__7100\ : Span4Mux_v
    port map (
            O => \N__30291\,
            I => \N__30288\
        );

    \I__7099\ : Odrv4
    port map (
            O => \N__30288\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_i_a4_4Z0Z_0\
        );

    \I__7098\ : InMux
    port map (
            O => \N__30285\,
            I => \N__30281\
        );

    \I__7097\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30276\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__30281\,
            I => \N__30273\
        );

    \I__7095\ : InMux
    port map (
            O => \N__30280\,
            I => \N__30270\
        );

    \I__7094\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30267\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__30276\,
            I => \N__30264\
        );

    \I__7092\ : Span4Mux_h
    port map (
            O => \N__30273\,
            I => \N__30261\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__30270\,
            I => \N__30256\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__30267\,
            I => \N__30256\
        );

    \I__7089\ : Odrv4
    port map (
            O => \N__30264\,
            I => \M_this_state_d62\
        );

    \I__7088\ : Odrv4
    port map (
            O => \N__30261\,
            I => \M_this_state_d62\
        );

    \I__7087\ : Odrv4
    port map (
            O => \N__30256\,
            I => \M_this_state_d62\
        );

    \I__7086\ : InMux
    port map (
            O => \N__30249\,
            I => \N__30246\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__30246\,
            I => \M_this_data_tmp_qZ0Z_4\
        );

    \I__7084\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30240\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__30240\,
            I => \M_this_data_tmp_qZ0Z_0\
        );

    \I__7082\ : CEMux
    port map (
            O => \N__30237\,
            I => \N__30234\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__30234\,
            I => \N__30231\
        );

    \I__7080\ : Span4Mux_v
    port map (
            O => \N__30231\,
            I => \N__30225\
        );

    \I__7079\ : CEMux
    port map (
            O => \N__30230\,
            I => \N__30222\
        );

    \I__7078\ : CEMux
    port map (
            O => \N__30229\,
            I => \N__30219\
        );

    \I__7077\ : CEMux
    port map (
            O => \N__30228\,
            I => \N__30216\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__30225\,
            I => \N__30212\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__30222\,
            I => \N__30209\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__30219\,
            I => \N__30206\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__30216\,
            I => \N__30203\
        );

    \I__7072\ : CEMux
    port map (
            O => \N__30215\,
            I => \N__30200\
        );

    \I__7071\ : Span4Mux_h
    port map (
            O => \N__30212\,
            I => \N__30197\
        );

    \I__7070\ : Span4Mux_v
    port map (
            O => \N__30209\,
            I => \N__30194\
        );

    \I__7069\ : Span4Mux_h
    port map (
            O => \N__30206\,
            I => \N__30191\
        );

    \I__7068\ : Span4Mux_h
    port map (
            O => \N__30203\,
            I => \N__30188\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__30200\,
            I => \N__30185\
        );

    \I__7066\ : Odrv4
    port map (
            O => \N__30197\,
            I => \N_1412_0\
        );

    \I__7065\ : Odrv4
    port map (
            O => \N__30194\,
            I => \N_1412_0\
        );

    \I__7064\ : Odrv4
    port map (
            O => \N__30191\,
            I => \N_1412_0\
        );

    \I__7063\ : Odrv4
    port map (
            O => \N__30188\,
            I => \N_1412_0\
        );

    \I__7062\ : Odrv12
    port map (
            O => \N__30185\,
            I => \N_1412_0\
        );

    \I__7061\ : InMux
    port map (
            O => \N__30174\,
            I => \N__30171\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__30171\,
            I => \N__30168\
        );

    \I__7059\ : Span4Mux_h
    port map (
            O => \N__30168\,
            I => \N__30165\
        );

    \I__7058\ : Odrv4
    port map (
            O => \N__30165\,
            I => \M_this_data_tmp_qZ0Z_3\
        );

    \I__7057\ : InMux
    port map (
            O => \N__30162\,
            I => \N__30159\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__30159\,
            I => \N__30156\
        );

    \I__7055\ : Span4Mux_h
    port map (
            O => \N__30156\,
            I => \N__30153\
        );

    \I__7054\ : Odrv4
    port map (
            O => \N__30153\,
            I => \M_this_oam_ram_write_data_3\
        );

    \I__7053\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30147\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__30147\,
            I => \N__30144\
        );

    \I__7051\ : Span4Mux_h
    port map (
            O => \N__30144\,
            I => \N__30141\
        );

    \I__7050\ : Odrv4
    port map (
            O => \N__30141\,
            I => \M_this_oam_ram_write_data_10\
        );

    \I__7049\ : InMux
    port map (
            O => \N__30138\,
            I => \N__30135\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__30135\,
            I => \M_this_data_tmp_qZ0Z_10\
        );

    \I__7047\ : InMux
    port map (
            O => \N__30132\,
            I => \N__30129\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__30129\,
            I => \N__30126\
        );

    \I__7045\ : Span4Mux_h
    port map (
            O => \N__30126\,
            I => \N__30123\
        );

    \I__7044\ : Odrv4
    port map (
            O => \N__30123\,
            I => \M_this_oam_ram_write_data_11\
        );

    \I__7043\ : CascadeMux
    port map (
            O => \N__30120\,
            I => \N__30117\
        );

    \I__7042\ : CascadeBuf
    port map (
            O => \N__30117\,
            I => \N__30114\
        );

    \I__7041\ : CascadeMux
    port map (
            O => \N__30114\,
            I => \N__30111\
        );

    \I__7040\ : InMux
    port map (
            O => \N__30111\,
            I => \N__30107\
        );

    \I__7039\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30103\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__30107\,
            I => \N__30100\
        );

    \I__7037\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30097\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__30103\,
            I => \N__30094\
        );

    \I__7035\ : Span4Mux_v
    port map (
            O => \N__30100\,
            I => \N__30091\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__30097\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__7033\ : Odrv4
    port map (
            O => \N__30094\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__7032\ : Odrv4
    port map (
            O => \N__30091\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__7031\ : CascadeMux
    port map (
            O => \N__30084\,
            I => \N__30081\
        );

    \I__7030\ : CascadeBuf
    port map (
            O => \N__30081\,
            I => \N__30078\
        );

    \I__7029\ : CascadeMux
    port map (
            O => \N__30078\,
            I => \N__30074\
        );

    \I__7028\ : InMux
    port map (
            O => \N__30077\,
            I => \N__30071\
        );

    \I__7027\ : InMux
    port map (
            O => \N__30074\,
            I => \N__30068\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__30071\,
            I => \N__30063\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__30068\,
            I => \N__30060\
        );

    \I__7024\ : InMux
    port map (
            O => \N__30067\,
            I => \N__30055\
        );

    \I__7023\ : InMux
    port map (
            O => \N__30066\,
            I => \N__30055\
        );

    \I__7022\ : Span4Mux_h
    port map (
            O => \N__30063\,
            I => \N__30052\
        );

    \I__7021\ : Span4Mux_v
    port map (
            O => \N__30060\,
            I => \N__30049\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__30055\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__7019\ : Odrv4
    port map (
            O => \N__30052\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__7018\ : Odrv4
    port map (
            O => \N__30049\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__7017\ : InMux
    port map (
            O => \N__30042\,
            I => \N__30039\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__30039\,
            I => \M_this_data_tmp_qZ0Z_11\
        );

    \I__7015\ : InMux
    port map (
            O => \N__30036\,
            I => \N__30033\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__30033\,
            I => \M_this_data_count_q_cry_0_THRU_CO\
        );

    \I__7013\ : CascadeMux
    port map (
            O => \N__30030\,
            I => \N__30026\
        );

    \I__7012\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30022\
        );

    \I__7011\ : InMux
    port map (
            O => \N__30026\,
            I => \N__30019\
        );

    \I__7010\ : InMux
    port map (
            O => \N__30025\,
            I => \N__30016\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__30022\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__30019\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__30016\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__7006\ : CascadeMux
    port map (
            O => \N__30009\,
            I => \N__30006\
        );

    \I__7005\ : InMux
    port map (
            O => \N__30006\,
            I => \N__30003\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__30003\,
            I => \M_this_data_count_q_cry_2_THRU_CO\
        );

    \I__7003\ : CascadeMux
    port map (
            O => \N__30000\,
            I => \N__29995\
        );

    \I__7002\ : CascadeMux
    port map (
            O => \N__29999\,
            I => \N__29992\
        );

    \I__7001\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29989\
        );

    \I__7000\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29986\
        );

    \I__6999\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29983\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__29989\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__29986\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__29983\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__6995\ : InMux
    port map (
            O => \N__29976\,
            I => \N__29973\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__29973\,
            I => \M_this_data_count_q_cry_3_THRU_CO\
        );

    \I__6993\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29965\
        );

    \I__6992\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29962\
        );

    \I__6991\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29959\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__29965\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__29962\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__29959\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__6987\ : InMux
    port map (
            O => \N__29952\,
            I => \N__29949\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__29949\,
            I => \M_this_data_count_q_cry_4_THRU_CO\
        );

    \I__6985\ : CascadeMux
    port map (
            O => \N__29946\,
            I => \N__29942\
        );

    \I__6984\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29938\
        );

    \I__6983\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29935\
        );

    \I__6982\ : InMux
    port map (
            O => \N__29941\,
            I => \N__29932\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__29938\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__29935\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__29932\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__6978\ : InMux
    port map (
            O => \N__29925\,
            I => \N__29922\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__29922\,
            I => \M_this_data_count_q_cry_5_THRU_CO\
        );

    \I__6976\ : InMux
    port map (
            O => \N__29919\,
            I => \N__29914\
        );

    \I__6975\ : InMux
    port map (
            O => \N__29918\,
            I => \N__29911\
        );

    \I__6974\ : InMux
    port map (
            O => \N__29917\,
            I => \N__29908\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__29914\,
            I => \N__29905\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__29911\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__29908\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__6970\ : Odrv4
    port map (
            O => \N__29905\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__6969\ : InMux
    port map (
            O => \N__29898\,
            I => \N__29895\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__29895\,
            I => \N__29892\
        );

    \I__6967\ : Span4Mux_h
    port map (
            O => \N__29892\,
            I => \N__29889\
        );

    \I__6966\ : Odrv4
    port map (
            O => \N__29889\,
            I => \M_this_oam_ram_write_data_4\
        );

    \I__6965\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29883\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__29883\,
            I => \N__29880\
        );

    \I__6963\ : Span4Mux_h
    port map (
            O => \N__29880\,
            I => \N__29877\
        );

    \I__6962\ : Span4Mux_v
    port map (
            O => \N__29877\,
            I => \N__29874\
        );

    \I__6961\ : Odrv4
    port map (
            O => \N__29874\,
            I => \M_this_data_tmp_qZ0Z_7\
        );

    \I__6960\ : InMux
    port map (
            O => \N__29871\,
            I => \N__29868\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__29868\,
            I => \N__29865\
        );

    \I__6958\ : Span4Mux_h
    port map (
            O => \N__29865\,
            I => \N__29862\
        );

    \I__6957\ : Odrv4
    port map (
            O => \N__29862\,
            I => \M_this_oam_ram_write_data_7\
        );

    \I__6956\ : InMux
    port map (
            O => \N__29859\,
            I => \N__29856\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__29856\,
            I => \N__29853\
        );

    \I__6954\ : Odrv12
    port map (
            O => \N__29853\,
            I => \M_this_oam_ram_write_data_8\
        );

    \I__6953\ : InMux
    port map (
            O => \N__29850\,
            I => \N__29847\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__29847\,
            I => \N__29844\
        );

    \I__6951\ : Span4Mux_h
    port map (
            O => \N__29844\,
            I => \N__29841\
        );

    \I__6950\ : Odrv4
    port map (
            O => \N__29841\,
            I => \M_this_oam_ram_write_data_0\
        );

    \I__6949\ : CascadeMux
    port map (
            O => \N__29838\,
            I => \N__29835\
        );

    \I__6948\ : InMux
    port map (
            O => \N__29835\,
            I => \N__29832\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__29832\,
            I => \N__29828\
        );

    \I__6946\ : InMux
    port map (
            O => \N__29831\,
            I => \N__29825\
        );

    \I__6945\ : Odrv4
    port map (
            O => \N__29828\,
            I => \M_this_data_count_qZ0Z_14\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__29825\,
            I => \M_this_data_count_qZ0Z_14\
        );

    \I__6943\ : InMux
    port map (
            O => \N__29820\,
            I => \N__29816\
        );

    \I__6942\ : InMux
    port map (
            O => \N__29819\,
            I => \N__29812\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__29816\,
            I => \N__29809\
        );

    \I__6940\ : InMux
    port map (
            O => \N__29815\,
            I => \N__29806\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__29812\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__6938\ : Odrv4
    port map (
            O => \N__29809\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__29806\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__6936\ : InMux
    port map (
            O => \N__29799\,
            I => \N__29795\
        );

    \I__6935\ : CascadeMux
    port map (
            O => \N__29798\,
            I => \N__29792\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__29795\,
            I => \N__29789\
        );

    \I__6933\ : InMux
    port map (
            O => \N__29792\,
            I => \N__29786\
        );

    \I__6932\ : Odrv4
    port map (
            O => \N__29789\,
            I => \M_this_data_count_qZ0Z_15\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__29786\,
            I => \M_this_data_count_qZ0Z_15\
        );

    \I__6930\ : CascadeMux
    port map (
            O => \N__29781\,
            I => \N__29778\
        );

    \I__6929\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29775\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__29775\,
            I => \N__29771\
        );

    \I__6927\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29768\
        );

    \I__6926\ : Odrv12
    port map (
            O => \N__29771\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__29768\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__6924\ : InMux
    port map (
            O => \N__29763\,
            I => \N__29758\
        );

    \I__6923\ : InMux
    port map (
            O => \N__29762\,
            I => \N__29755\
        );

    \I__6922\ : InMux
    port map (
            O => \N__29761\,
            I => \N__29752\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__29758\,
            I => \N__29747\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__29755\,
            I => \N__29744\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__29752\,
            I => \N__29741\
        );

    \I__6918\ : InMux
    port map (
            O => \N__29751\,
            I => \N__29736\
        );

    \I__6917\ : InMux
    port map (
            O => \N__29750\,
            I => \N__29736\
        );

    \I__6916\ : Odrv4
    port map (
            O => \N__29747\,
            I => \this_vga_signals.N_745\
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__29744\,
            I => \this_vga_signals.N_745\
        );

    \I__6914\ : Odrv4
    port map (
            O => \N__29741\,
            I => \this_vga_signals.N_745\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__29736\,
            I => \this_vga_signals.N_745\
        );

    \I__6912\ : InMux
    port map (
            O => \N__29727\,
            I => \N__29724\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__29724\,
            I => \this_vga_signals.M_this_external_address_qlde_i_0_aZ0Z2\
        );

    \I__6910\ : InMux
    port map (
            O => \N__29721\,
            I => \N__29718\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__29718\,
            I => \this_vga_signals.N_442_0\
        );

    \I__6908\ : InMux
    port map (
            O => \N__29715\,
            I => \N__29712\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__29712\,
            I => \N__29707\
        );

    \I__6906\ : InMux
    port map (
            O => \N__29711\,
            I => \N__29704\
        );

    \I__6905\ : InMux
    port map (
            O => \N__29710\,
            I => \N__29701\
        );

    \I__6904\ : Span4Mux_v
    port map (
            O => \N__29707\,
            I => \N__29692\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__29704\,
            I => \N__29692\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__29701\,
            I => \N__29689\
        );

    \I__6901\ : InMux
    port map (
            O => \N__29700\,
            I => \N__29686\
        );

    \I__6900\ : CascadeMux
    port map (
            O => \N__29699\,
            I => \N__29681\
        );

    \I__6899\ : IoInMux
    port map (
            O => \N__29698\,
            I => \N__29675\
        );

    \I__6898\ : InMux
    port map (
            O => \N__29697\,
            I => \N__29672\
        );

    \I__6897\ : Span4Mux_h
    port map (
            O => \N__29692\,
            I => \N__29669\
        );

    \I__6896\ : Span4Mux_h
    port map (
            O => \N__29689\,
            I => \N__29666\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__29686\,
            I => \N__29663\
        );

    \I__6894\ : InMux
    port map (
            O => \N__29685\,
            I => \N__29657\
        );

    \I__6893\ : InMux
    port map (
            O => \N__29684\,
            I => \N__29657\
        );

    \I__6892\ : InMux
    port map (
            O => \N__29681\,
            I => \N__29652\
        );

    \I__6891\ : InMux
    port map (
            O => \N__29680\,
            I => \N__29652\
        );

    \I__6890\ : InMux
    port map (
            O => \N__29679\,
            I => \N__29649\
        );

    \I__6889\ : InMux
    port map (
            O => \N__29678\,
            I => \N__29646\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__29675\,
            I => \N__29643\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__29672\,
            I => \N__29640\
        );

    \I__6886\ : Span4Mux_h
    port map (
            O => \N__29669\,
            I => \N__29633\
        );

    \I__6885\ : Span4Mux_h
    port map (
            O => \N__29666\,
            I => \N__29633\
        );

    \I__6884\ : Span4Mux_h
    port map (
            O => \N__29663\,
            I => \N__29633\
        );

    \I__6883\ : InMux
    port map (
            O => \N__29662\,
            I => \N__29630\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__29657\,
            I => \N__29619\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__29652\,
            I => \N__29619\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__29649\,
            I => \N__29619\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__29646\,
            I => \N__29619\
        );

    \I__6878\ : Span12Mux_s9_h
    port map (
            O => \N__29643\,
            I => \N__29619\
        );

    \I__6877\ : Odrv4
    port map (
            O => \N__29640\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6876\ : Odrv4
    port map (
            O => \N__29633\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__29630\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6874\ : Odrv12
    port map (
            O => \N__29619\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6873\ : CascadeMux
    port map (
            O => \N__29610\,
            I => \this_vga_signals.M_this_external_address_qlde_i_0_aZ0Z2_cascade_\
        );

    \I__6872\ : InMux
    port map (
            O => \N__29607\,
            I => \N__29604\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__29604\,
            I => \this_vga_signals.M_this_data_count_qlde_iZ0Z_1\
        );

    \I__6870\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29598\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__29598\,
            I => \N__29594\
        );

    \I__6868\ : InMux
    port map (
            O => \N__29597\,
            I => \N__29591\
        );

    \I__6867\ : Odrv4
    port map (
            O => \N__29594\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__29591\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__6865\ : InMux
    port map (
            O => \N__29586\,
            I => \N__29581\
        );

    \I__6864\ : InMux
    port map (
            O => \N__29585\,
            I => \N__29578\
        );

    \I__6863\ : InMux
    port map (
            O => \N__29584\,
            I => \N__29575\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__29581\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__29578\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__29575\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__6859\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29565\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__29565\,
            I => \N__29562\
        );

    \I__6857\ : Odrv4
    port map (
            O => \N__29562\,
            I => \M_this_state_d62_11\
        );

    \I__6856\ : CascadeMux
    port map (
            O => \N__29559\,
            I => \M_this_state_d62_8_cascade_\
        );

    \I__6855\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29553\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__29553\,
            I => \N__29549\
        );

    \I__6853\ : InMux
    port map (
            O => \N__29552\,
            I => \N__29545\
        );

    \I__6852\ : Span4Mux_h
    port map (
            O => \N__29549\,
            I => \N__29542\
        );

    \I__6851\ : InMux
    port map (
            O => \N__29548\,
            I => \N__29539\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__29545\,
            I => \N__29536\
        );

    \I__6849\ : Odrv4
    port map (
            O => \N__29542\,
            I => \un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__29539\,
            I => \un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2\
        );

    \I__6847\ : Odrv12
    port map (
            O => \N__29536\,
            I => \un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2\
        );

    \I__6846\ : CascadeMux
    port map (
            O => \N__29529\,
            I => \M_this_state_d62_cascade_\
        );

    \I__6845\ : CascadeMux
    port map (
            O => \N__29526\,
            I => \N__29523\
        );

    \I__6844\ : InMux
    port map (
            O => \N__29523\,
            I => \N__29520\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__29520\,
            I => \N__29515\
        );

    \I__6842\ : InMux
    port map (
            O => \N__29519\,
            I => \N__29512\
        );

    \I__6841\ : InMux
    port map (
            O => \N__29518\,
            I => \N__29509\
        );

    \I__6840\ : Span4Mux_v
    port map (
            O => \N__29515\,
            I => \N__29506\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__29512\,
            I => \N__29503\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__29509\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__6837\ : Odrv4
    port map (
            O => \N__29506\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__6836\ : Odrv4
    port map (
            O => \N__29503\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__6835\ : InMux
    port map (
            O => \N__29496\,
            I => \N__29493\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__29493\,
            I => \N__29489\
        );

    \I__6833\ : InMux
    port map (
            O => \N__29492\,
            I => \N__29486\
        );

    \I__6832\ : Odrv4
    port map (
            O => \N__29489\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__29486\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__6830\ : CascadeMux
    port map (
            O => \N__29481\,
            I => \N__29477\
        );

    \I__6829\ : InMux
    port map (
            O => \N__29480\,
            I => \N__29474\
        );

    \I__6828\ : InMux
    port map (
            O => \N__29477\,
            I => \N__29471\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__29474\,
            I => \N__29468\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__29471\,
            I => \N__29465\
        );

    \I__6825\ : Odrv4
    port map (
            O => \N__29468\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__6824\ : Odrv4
    port map (
            O => \N__29465\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__6823\ : CascadeMux
    port map (
            O => \N__29460\,
            I => \N__29457\
        );

    \I__6822\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29454\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__29454\,
            I => \N__29450\
        );

    \I__6820\ : InMux
    port map (
            O => \N__29453\,
            I => \N__29447\
        );

    \I__6819\ : Odrv4
    port map (
            O => \N__29450\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__29447\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__6817\ : InMux
    port map (
            O => \N__29442\,
            I => \N__29439\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__29439\,
            I => \M_this_state_d62_10\
        );

    \I__6815\ : InMux
    port map (
            O => \N__29436\,
            I => \N__29433\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__29433\,
            I => \M_this_state_d62_9\
        );

    \I__6813\ : InMux
    port map (
            O => \N__29430\,
            I => \N__29427\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__29427\,
            I => \N__29424\
        );

    \I__6811\ : Span4Mux_h
    port map (
            O => \N__29424\,
            I => \N__29421\
        );

    \I__6810\ : Odrv4
    port map (
            O => \N__29421\,
            I => \M_this_oam_ram_write_data_24\
        );

    \I__6809\ : InMux
    port map (
            O => \N__29418\,
            I => \N__29413\
        );

    \I__6808\ : InMux
    port map (
            O => \N__29417\,
            I => \N__29410\
        );

    \I__6807\ : InMux
    port map (
            O => \N__29416\,
            I => \N__29407\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__29413\,
            I => \N__29403\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__29410\,
            I => \N__29397\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__29407\,
            I => \N__29397\
        );

    \I__6803\ : InMux
    port map (
            O => \N__29406\,
            I => \N__29394\
        );

    \I__6802\ : Span4Mux_h
    port map (
            O => \N__29403\,
            I => \N__29391\
        );

    \I__6801\ : InMux
    port map (
            O => \N__29402\,
            I => \N__29388\
        );

    \I__6800\ : Span4Mux_h
    port map (
            O => \N__29397\,
            I => \N__29385\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__29394\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6798\ : Odrv4
    port map (
            O => \N__29391\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__29388\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__29385\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6795\ : CascadeMux
    port map (
            O => \N__29376\,
            I => \N__29370\
        );

    \I__6794\ : InMux
    port map (
            O => \N__29375\,
            I => \N__29367\
        );

    \I__6793\ : CascadeMux
    port map (
            O => \N__29374\,
            I => \N__29364\
        );

    \I__6792\ : InMux
    port map (
            O => \N__29373\,
            I => \N__29360\
        );

    \I__6791\ : InMux
    port map (
            O => \N__29370\,
            I => \N__29357\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__29367\,
            I => \N__29354\
        );

    \I__6789\ : InMux
    port map (
            O => \N__29364\,
            I => \N__29349\
        );

    \I__6788\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29349\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__29360\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__29357\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__6785\ : Odrv4
    port map (
            O => \N__29354\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__29349\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__6783\ : CascadeMux
    port map (
            O => \N__29340\,
            I => \this_vga_signals.N_469_0_cascade_\
        );

    \I__6782\ : CascadeMux
    port map (
            O => \N__29337\,
            I => \this_vga_signals.N_506_cascade_\
        );

    \I__6781\ : InMux
    port map (
            O => \N__29334\,
            I => \N__29331\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__29331\,
            I => \N__29326\
        );

    \I__6779\ : InMux
    port map (
            O => \N__29330\,
            I => \N__29323\
        );

    \I__6778\ : InMux
    port map (
            O => \N__29329\,
            I => \N__29320\
        );

    \I__6777\ : Span4Mux_h
    port map (
            O => \N__29326\,
            I => \N__29312\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__29323\,
            I => \N__29307\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__29320\,
            I => \N__29307\
        );

    \I__6774\ : InMux
    port map (
            O => \N__29319\,
            I => \N__29300\
        );

    \I__6773\ : InMux
    port map (
            O => \N__29318\,
            I => \N__29300\
        );

    \I__6772\ : InMux
    port map (
            O => \N__29317\,
            I => \N__29300\
        );

    \I__6771\ : InMux
    port map (
            O => \N__29316\,
            I => \N__29292\
        );

    \I__6770\ : InMux
    port map (
            O => \N__29315\,
            I => \N__29292\
        );

    \I__6769\ : Span4Mux_v
    port map (
            O => \N__29312\,
            I => \N__29289\
        );

    \I__6768\ : Span4Mux_v
    port map (
            O => \N__29307\,
            I => \N__29284\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__29300\,
            I => \N__29284\
        );

    \I__6766\ : InMux
    port map (
            O => \N__29299\,
            I => \N__29277\
        );

    \I__6765\ : InMux
    port map (
            O => \N__29298\,
            I => \N__29277\
        );

    \I__6764\ : InMux
    port map (
            O => \N__29297\,
            I => \N__29277\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__29292\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__6762\ : Odrv4
    port map (
            O => \N__29289\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__6761\ : Odrv4
    port map (
            O => \N__29284\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__29277\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__6759\ : CascadeMux
    port map (
            O => \N__29268\,
            I => \this_ppu.un1_oam_data_c2_cascade_\
        );

    \I__6758\ : InMux
    port map (
            O => \N__29265\,
            I => \N__29262\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__29262\,
            I => \this_ppu.un1_M_vaddress_q_3_6\
        );

    \I__6756\ : InMux
    port map (
            O => \N__29259\,
            I => \N__29256\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__29256\,
            I => \M_this_data_tmp_qZ0Z_23\
        );

    \I__6754\ : InMux
    port map (
            O => \N__29253\,
            I => \N__29250\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__29250\,
            I => \N__29247\
        );

    \I__6752\ : Span4Mux_h
    port map (
            O => \N__29247\,
            I => \N__29244\
        );

    \I__6751\ : Odrv4
    port map (
            O => \N__29244\,
            I => \M_this_oam_ram_write_data_23\
        );

    \I__6750\ : InMux
    port map (
            O => \N__29241\,
            I => \N__29236\
        );

    \I__6749\ : InMux
    port map (
            O => \N__29240\,
            I => \N__29231\
        );

    \I__6748\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29231\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__29236\,
            I => \N__29228\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__29231\,
            I => \N__29225\
        );

    \I__6745\ : Span12Mux_s7_v
    port map (
            O => \N__29228\,
            I => \N__29222\
        );

    \I__6744\ : Span4Mux_v
    port map (
            O => \N__29225\,
            I => \N__29219\
        );

    \I__6743\ : Odrv12
    port map (
            O => \N__29222\,
            I => \M_this_oam_ram_read_data_22\
        );

    \I__6742\ : Odrv4
    port map (
            O => \N__29219\,
            I => \M_this_oam_ram_read_data_22\
        );

    \I__6741\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29210\
        );

    \I__6740\ : CascadeMux
    port map (
            O => \N__29213\,
            I => \N__29207\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__29210\,
            I => \N__29204\
        );

    \I__6738\ : InMux
    port map (
            O => \N__29207\,
            I => \N__29201\
        );

    \I__6737\ : Span4Mux_h
    port map (
            O => \N__29204\,
            I => \N__29198\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__29201\,
            I => \N__29195\
        );

    \I__6735\ : Span4Mux_h
    port map (
            O => \N__29198\,
            I => \N__29192\
        );

    \I__6734\ : Span4Mux_v
    port map (
            O => \N__29195\,
            I => \N__29189\
        );

    \I__6733\ : Odrv4
    port map (
            O => \N__29192\,
            I => \M_this_oam_ram_read_data_23\
        );

    \I__6732\ : Odrv4
    port map (
            O => \N__29189\,
            I => \M_this_oam_ram_read_data_23\
        );

    \I__6731\ : InMux
    port map (
            O => \N__29184\,
            I => \N__29181\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__29181\,
            I => \this_ppu.un1_oam_data_c2\
        );

    \I__6729\ : InMux
    port map (
            O => \N__29178\,
            I => \N__29175\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__29175\,
            I => \this_ppu.un1_M_vaddress_q_3_7\
        );

    \I__6727\ : InMux
    port map (
            O => \N__29172\,
            I => \N__29169\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__29169\,
            I => \N__29166\
        );

    \I__6725\ : Odrv4
    port map (
            O => \N__29166\,
            I => \M_this_oam_ram_write_data_25\
        );

    \I__6724\ : CascadeMux
    port map (
            O => \N__29163\,
            I => \N__29160\
        );

    \I__6723\ : InMux
    port map (
            O => \N__29160\,
            I => \N__29157\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__29157\,
            I => \M_this_data_tmp_qZ0Z_17\
        );

    \I__6721\ : InMux
    port map (
            O => \N__29154\,
            I => \N__29151\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__29151\,
            I => \N__29148\
        );

    \I__6719\ : Span4Mux_h
    port map (
            O => \N__29148\,
            I => \N__29145\
        );

    \I__6718\ : Odrv4
    port map (
            O => \N__29145\,
            I => \M_this_oam_ram_write_data_17\
        );

    \I__6717\ : InMux
    port map (
            O => \N__29142\,
            I => \N__29139\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__29139\,
            I => \this_ppu.un1_M_vaddress_q_3_4\
        );

    \I__6715\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29133\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__29133\,
            I => \N__29130\
        );

    \I__6713\ : Odrv4
    port map (
            O => \N__29130\,
            I => \M_this_data_count_q_cry_12_THRU_CO\
        );

    \I__6712\ : InMux
    port map (
            O => \N__29127\,
            I => \M_this_data_count_q_cry_12\
        );

    \I__6711\ : IoInMux
    port map (
            O => \N__29124\,
            I => \N__29118\
        );

    \I__6710\ : SRMux
    port map (
            O => \N__29123\,
            I => \N__29114\
        );

    \I__6709\ : SRMux
    port map (
            O => \N__29122\,
            I => \N__29111\
        );

    \I__6708\ : SRMux
    port map (
            O => \N__29121\,
            I => \N__29108\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__29118\,
            I => \N__29103\
        );

    \I__6706\ : SRMux
    port map (
            O => \N__29117\,
            I => \N__29099\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__29114\,
            I => \N__29093\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__29111\,
            I => \N__29093\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__29108\,
            I => \N__29090\
        );

    \I__6702\ : SRMux
    port map (
            O => \N__29107\,
            I => \N__29087\
        );

    \I__6701\ : SRMux
    port map (
            O => \N__29106\,
            I => \N__29084\
        );

    \I__6700\ : IoSpan4Mux
    port map (
            O => \N__29103\,
            I => \N__29078\
        );

    \I__6699\ : SRMux
    port map (
            O => \N__29102\,
            I => \N__29075\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__29099\,
            I => \N__29072\
        );

    \I__6697\ : SRMux
    port map (
            O => \N__29098\,
            I => \N__29069\
        );

    \I__6696\ : Span4Mux_s3_v
    port map (
            O => \N__29093\,
            I => \N__29052\
        );

    \I__6695\ : Span4Mux_h
    port map (
            O => \N__29090\,
            I => \N__29052\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__29087\,
            I => \N__29052\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__29084\,
            I => \N__29052\
        );

    \I__6692\ : SRMux
    port map (
            O => \N__29083\,
            I => \N__29049\
        );

    \I__6691\ : SRMux
    port map (
            O => \N__29082\,
            I => \N__29043\
        );

    \I__6690\ : SRMux
    port map (
            O => \N__29081\,
            I => \N__29039\
        );

    \I__6689\ : Span4Mux_s2_h
    port map (
            O => \N__29078\,
            I => \N__29036\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__29075\,
            I => \N__29029\
        );

    \I__6687\ : Span4Mux_h
    port map (
            O => \N__29072\,
            I => \N__29029\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__29069\,
            I => \N__29029\
        );

    \I__6685\ : SRMux
    port map (
            O => \N__29068\,
            I => \N__29026\
        );

    \I__6684\ : SRMux
    port map (
            O => \N__29067\,
            I => \N__29020\
        );

    \I__6683\ : SRMux
    port map (
            O => \N__29066\,
            I => \N__29017\
        );

    \I__6682\ : SRMux
    port map (
            O => \N__29065\,
            I => \N__29012\
        );

    \I__6681\ : CascadeMux
    port map (
            O => \N__29064\,
            I => \N__29007\
        );

    \I__6680\ : CascadeMux
    port map (
            O => \N__29063\,
            I => \N__29004\
        );

    \I__6679\ : CascadeMux
    port map (
            O => \N__29062\,
            I => \N__28998\
        );

    \I__6678\ : SRMux
    port map (
            O => \N__29061\,
            I => \N__28995\
        );

    \I__6677\ : Span4Mux_v
    port map (
            O => \N__29052\,
            I => \N__28990\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__29049\,
            I => \N__28990\
        );

    \I__6675\ : CascadeMux
    port map (
            O => \N__29048\,
            I => \N__28986\
        );

    \I__6674\ : CascadeMux
    port map (
            O => \N__29047\,
            I => \N__28982\
        );

    \I__6673\ : CascadeMux
    port map (
            O => \N__29046\,
            I => \N__28977\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__29043\,
            I => \N__28974\
        );

    \I__6671\ : SRMux
    port map (
            O => \N__29042\,
            I => \N__28971\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__29039\,
            I => \N__28968\
        );

    \I__6669\ : Span4Mux_h
    port map (
            O => \N__29036\,
            I => \N__28961\
        );

    \I__6668\ : Span4Mux_v
    port map (
            O => \N__29029\,
            I => \N__28961\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__29026\,
            I => \N__28961\
        );

    \I__6666\ : SRMux
    port map (
            O => \N__29025\,
            I => \N__28958\
        );

    \I__6665\ : SRMux
    port map (
            O => \N__29024\,
            I => \N__28955\
        );

    \I__6664\ : SRMux
    port map (
            O => \N__29023\,
            I => \N__28952\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__29020\,
            I => \N__28949\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__29017\,
            I => \N__28946\
        );

    \I__6661\ : SRMux
    port map (
            O => \N__29016\,
            I => \N__28943\
        );

    \I__6660\ : SRMux
    port map (
            O => \N__29015\,
            I => \N__28940\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__29012\,
            I => \N__28931\
        );

    \I__6658\ : SRMux
    port map (
            O => \N__29011\,
            I => \N__28928\
        );

    \I__6657\ : InMux
    port map (
            O => \N__29010\,
            I => \N__28913\
        );

    \I__6656\ : InMux
    port map (
            O => \N__29007\,
            I => \N__28913\
        );

    \I__6655\ : InMux
    port map (
            O => \N__29004\,
            I => \N__28913\
        );

    \I__6654\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28913\
        );

    \I__6653\ : InMux
    port map (
            O => \N__29002\,
            I => \N__28913\
        );

    \I__6652\ : InMux
    port map (
            O => \N__29001\,
            I => \N__28913\
        );

    \I__6651\ : InMux
    port map (
            O => \N__28998\,
            I => \N__28913\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__28995\,
            I => \N__28910\
        );

    \I__6649\ : Span4Mux_v
    port map (
            O => \N__28990\,
            I => \N__28907\
        );

    \I__6648\ : InMux
    port map (
            O => \N__28989\,
            I => \N__28892\
        );

    \I__6647\ : InMux
    port map (
            O => \N__28986\,
            I => \N__28892\
        );

    \I__6646\ : InMux
    port map (
            O => \N__28985\,
            I => \N__28892\
        );

    \I__6645\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28892\
        );

    \I__6644\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28892\
        );

    \I__6643\ : InMux
    port map (
            O => \N__28980\,
            I => \N__28892\
        );

    \I__6642\ : InMux
    port map (
            O => \N__28977\,
            I => \N__28892\
        );

    \I__6641\ : Span4Mux_v
    port map (
            O => \N__28974\,
            I => \N__28887\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__28971\,
            I => \N__28887\
        );

    \I__6639\ : Span4Mux_v
    port map (
            O => \N__28968\,
            I => \N__28878\
        );

    \I__6638\ : Span4Mux_h
    port map (
            O => \N__28961\,
            I => \N__28878\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__28958\,
            I => \N__28878\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__28955\,
            I => \N__28878\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__28952\,
            I => \N__28875\
        );

    \I__6634\ : Span4Mux_v
    port map (
            O => \N__28949\,
            I => \N__28866\
        );

    \I__6633\ : Span4Mux_h
    port map (
            O => \N__28946\,
            I => \N__28866\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__28943\,
            I => \N__28866\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__28940\,
            I => \N__28866\
        );

    \I__6630\ : SRMux
    port map (
            O => \N__28939\,
            I => \N__28863\
        );

    \I__6629\ : SRMux
    port map (
            O => \N__28938\,
            I => \N__28860\
        );

    \I__6628\ : SRMux
    port map (
            O => \N__28937\,
            I => \N__28857\
        );

    \I__6627\ : SRMux
    port map (
            O => \N__28936\,
            I => \N__28854\
        );

    \I__6626\ : SRMux
    port map (
            O => \N__28935\,
            I => \N__28847\
        );

    \I__6625\ : SRMux
    port map (
            O => \N__28934\,
            I => \N__28844\
        );

    \I__6624\ : Span4Mux_v
    port map (
            O => \N__28931\,
            I => \N__28839\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__28928\,
            I => \N__28836\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__28913\,
            I => \N__28833\
        );

    \I__6621\ : Span4Mux_h
    port map (
            O => \N__28910\,
            I => \N__28826\
        );

    \I__6620\ : Span4Mux_h
    port map (
            O => \N__28907\,
            I => \N__28826\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__28892\,
            I => \N__28826\
        );

    \I__6618\ : Span4Mux_v
    port map (
            O => \N__28887\,
            I => \N__28813\
        );

    \I__6617\ : Span4Mux_v
    port map (
            O => \N__28878\,
            I => \N__28813\
        );

    \I__6616\ : Span4Mux_v
    port map (
            O => \N__28875\,
            I => \N__28813\
        );

    \I__6615\ : Span4Mux_v
    port map (
            O => \N__28866\,
            I => \N__28813\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__28863\,
            I => \N__28813\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__28860\,
            I => \N__28813\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__28857\,
            I => \N__28810\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__28854\,
            I => \N__28804\
        );

    \I__6610\ : SRMux
    port map (
            O => \N__28853\,
            I => \N__28801\
        );

    \I__6609\ : SRMux
    port map (
            O => \N__28852\,
            I => \N__28798\
        );

    \I__6608\ : SRMux
    port map (
            O => \N__28851\,
            I => \N__28795\
        );

    \I__6607\ : SRMux
    port map (
            O => \N__28850\,
            I => \N__28792\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__28847\,
            I => \N__28789\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__28844\,
            I => \N__28786\
        );

    \I__6604\ : SRMux
    port map (
            O => \N__28843\,
            I => \N__28783\
        );

    \I__6603\ : SRMux
    port map (
            O => \N__28842\,
            I => \N__28780\
        );

    \I__6602\ : Span4Mux_h
    port map (
            O => \N__28839\,
            I => \N__28772\
        );

    \I__6601\ : Span4Mux_h
    port map (
            O => \N__28836\,
            I => \N__28772\
        );

    \I__6600\ : Span4Mux_v
    port map (
            O => \N__28833\,
            I => \N__28767\
        );

    \I__6599\ : Span4Mux_v
    port map (
            O => \N__28826\,
            I => \N__28767\
        );

    \I__6598\ : Span4Mux_v
    port map (
            O => \N__28813\,
            I => \N__28764\
        );

    \I__6597\ : Span4Mux_v
    port map (
            O => \N__28810\,
            I => \N__28761\
        );

    \I__6596\ : CascadeMux
    port map (
            O => \N__28809\,
            I => \N__28758\
        );

    \I__6595\ : CascadeMux
    port map (
            O => \N__28808\,
            I => \N__28754\
        );

    \I__6594\ : CascadeMux
    port map (
            O => \N__28807\,
            I => \N__28750\
        );

    \I__6593\ : Span4Mux_h
    port map (
            O => \N__28804\,
            I => \N__28746\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__28801\,
            I => \N__28743\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__28798\,
            I => \N__28738\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__28795\,
            I => \N__28738\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__28792\,
            I => \N__28733\
        );

    \I__6588\ : Span4Mux_v
    port map (
            O => \N__28789\,
            I => \N__28724\
        );

    \I__6587\ : Span4Mux_h
    port map (
            O => \N__28786\,
            I => \N__28724\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__28783\,
            I => \N__28724\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__28780\,
            I => \N__28724\
        );

    \I__6584\ : SRMux
    port map (
            O => \N__28779\,
            I => \N__28721\
        );

    \I__6583\ : SRMux
    port map (
            O => \N__28778\,
            I => \N__28718\
        );

    \I__6582\ : IoInMux
    port map (
            O => \N__28777\,
            I => \N__28714\
        );

    \I__6581\ : Span4Mux_h
    port map (
            O => \N__28772\,
            I => \N__28711\
        );

    \I__6580\ : Span4Mux_v
    port map (
            O => \N__28767\,
            I => \N__28704\
        );

    \I__6579\ : Span4Mux_h
    port map (
            O => \N__28764\,
            I => \N__28704\
        );

    \I__6578\ : Span4Mux_h
    port map (
            O => \N__28761\,
            I => \N__28704\
        );

    \I__6577\ : InMux
    port map (
            O => \N__28758\,
            I => \N__28691\
        );

    \I__6576\ : InMux
    port map (
            O => \N__28757\,
            I => \N__28691\
        );

    \I__6575\ : InMux
    port map (
            O => \N__28754\,
            I => \N__28691\
        );

    \I__6574\ : InMux
    port map (
            O => \N__28753\,
            I => \N__28691\
        );

    \I__6573\ : InMux
    port map (
            O => \N__28750\,
            I => \N__28691\
        );

    \I__6572\ : InMux
    port map (
            O => \N__28749\,
            I => \N__28691\
        );

    \I__6571\ : Span4Mux_v
    port map (
            O => \N__28746\,
            I => \N__28686\
        );

    \I__6570\ : Span4Mux_h
    port map (
            O => \N__28743\,
            I => \N__28686\
        );

    \I__6569\ : Span4Mux_v
    port map (
            O => \N__28738\,
            I => \N__28683\
        );

    \I__6568\ : SRMux
    port map (
            O => \N__28737\,
            I => \N__28680\
        );

    \I__6567\ : SRMux
    port map (
            O => \N__28736\,
            I => \N__28677\
        );

    \I__6566\ : Span4Mux_v
    port map (
            O => \N__28733\,
            I => \N__28670\
        );

    \I__6565\ : Span4Mux_v
    port map (
            O => \N__28724\,
            I => \N__28670\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__28721\,
            I => \N__28670\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__28718\,
            I => \N__28667\
        );

    \I__6562\ : SRMux
    port map (
            O => \N__28717\,
            I => \N__28664\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__28714\,
            I => \N__28661\
        );

    \I__6560\ : Span4Mux_v
    port map (
            O => \N__28711\,
            I => \N__28653\
        );

    \I__6559\ : Span4Mux_h
    port map (
            O => \N__28704\,
            I => \N__28653\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__28691\,
            I => \N__28653\
        );

    \I__6557\ : Sp12to4
    port map (
            O => \N__28686\,
            I => \N__28649\
        );

    \I__6556\ : Span4Mux_v
    port map (
            O => \N__28683\,
            I => \N__28642\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__28680\,
            I => \N__28642\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__28677\,
            I => \N__28642\
        );

    \I__6553\ : Span4Mux_v
    port map (
            O => \N__28670\,
            I => \N__28635\
        );

    \I__6552\ : Span4Mux_v
    port map (
            O => \N__28667\,
            I => \N__28635\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__28664\,
            I => \N__28635\
        );

    \I__6550\ : IoSpan4Mux
    port map (
            O => \N__28661\,
            I => \N__28632\
        );

    \I__6549\ : SRMux
    port map (
            O => \N__28660\,
            I => \N__28629\
        );

    \I__6548\ : Span4Mux_h
    port map (
            O => \N__28653\,
            I => \N__28626\
        );

    \I__6547\ : SRMux
    port map (
            O => \N__28652\,
            I => \N__28623\
        );

    \I__6546\ : Span12Mux_h
    port map (
            O => \N__28649\,
            I => \N__28620\
        );

    \I__6545\ : Span4Mux_v
    port map (
            O => \N__28642\,
            I => \N__28617\
        );

    \I__6544\ : Span4Mux_h
    port map (
            O => \N__28635\,
            I => \N__28614\
        );

    \I__6543\ : Span4Mux_s3_h
    port map (
            O => \N__28632\,
            I => \N__28611\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__28629\,
            I => \N__28608\
        );

    \I__6541\ : Span4Mux_h
    port map (
            O => \N__28626\,
            I => \N__28603\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__28623\,
            I => \N__28603\
        );

    \I__6539\ : Span12Mux_v
    port map (
            O => \N__28620\,
            I => \N__28600\
        );

    \I__6538\ : Span4Mux_v
    port map (
            O => \N__28617\,
            I => \N__28595\
        );

    \I__6537\ : Span4Mux_v
    port map (
            O => \N__28614\,
            I => \N__28595\
        );

    \I__6536\ : Span4Mux_v
    port map (
            O => \N__28611\,
            I => \N__28590\
        );

    \I__6535\ : Span4Mux_v
    port map (
            O => \N__28608\,
            I => \N__28590\
        );

    \I__6534\ : Span4Mux_h
    port map (
            O => \N__28603\,
            I => \N__28587\
        );

    \I__6533\ : Odrv12
    port map (
            O => \N__28600\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6532\ : Odrv4
    port map (
            O => \N__28595\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6531\ : Odrv4
    port map (
            O => \N__28590\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6530\ : Odrv4
    port map (
            O => \N__28587\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6529\ : InMux
    port map (
            O => \N__28578\,
            I => \N__28575\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__28575\,
            I => \N__28572\
        );

    \I__6527\ : Odrv12
    port map (
            O => \N__28572\,
            I => \M_this_data_count_q_s_14\
        );

    \I__6526\ : InMux
    port map (
            O => \N__28569\,
            I => \M_this_data_count_q_cry_13\
        );

    \I__6525\ : InMux
    port map (
            O => \N__28566\,
            I => \M_this_data_count_q_cry_14\
        );

    \I__6524\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28560\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__28560\,
            I => \N__28557\
        );

    \I__6522\ : Span4Mux_h
    port map (
            O => \N__28557\,
            I => \N__28554\
        );

    \I__6521\ : Odrv4
    port map (
            O => \N__28554\,
            I => \M_this_data_count_q_s_15\
        );

    \I__6520\ : InMux
    port map (
            O => \N__28551\,
            I => \N__28548\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__28548\,
            I => \N__28542\
        );

    \I__6518\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28537\
        );

    \I__6517\ : InMux
    port map (
            O => \N__28546\,
            I => \N__28537\
        );

    \I__6516\ : InMux
    port map (
            O => \N__28545\,
            I => \N__28534\
        );

    \I__6515\ : Odrv4
    port map (
            O => \N__28542\,
            I => \this_vga_signals.N_431_0\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__28537\,
            I => \this_vga_signals.N_431_0\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__28534\,
            I => \this_vga_signals.N_431_0\
        );

    \I__6512\ : InMux
    port map (
            O => \N__28527\,
            I => \N__28524\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28518\
        );

    \I__6510\ : InMux
    port map (
            O => \N__28523\,
            I => \N__28511\
        );

    \I__6509\ : InMux
    port map (
            O => \N__28522\,
            I => \N__28511\
        );

    \I__6508\ : InMux
    port map (
            O => \N__28521\,
            I => \N__28511\
        );

    \I__6507\ : Span4Mux_v
    port map (
            O => \N__28518\,
            I => \N__28507\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__28511\,
            I => \N__28504\
        );

    \I__6505\ : InMux
    port map (
            O => \N__28510\,
            I => \N__28501\
        );

    \I__6504\ : Odrv4
    port map (
            O => \N__28507\,
            I => \this_vga_signals.N_428_0\
        );

    \I__6503\ : Odrv12
    port map (
            O => \N__28504\,
            I => \this_vga_signals.N_428_0\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__28501\,
            I => \this_vga_signals.N_428_0\
        );

    \I__6501\ : InMux
    port map (
            O => \N__28494\,
            I => \N__28490\
        );

    \I__6500\ : InMux
    port map (
            O => \N__28493\,
            I => \N__28486\
        );

    \I__6499\ : LocalMux
    port map (
            O => \N__28490\,
            I => \N__28482\
        );

    \I__6498\ : InMux
    port map (
            O => \N__28489\,
            I => \N__28479\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__28486\,
            I => \N__28476\
        );

    \I__6496\ : InMux
    port map (
            O => \N__28485\,
            I => \N__28473\
        );

    \I__6495\ : Span4Mux_h
    port map (
            O => \N__28482\,
            I => \N__28470\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__28479\,
            I => \N__28467\
        );

    \I__6493\ : Span4Mux_v
    port map (
            O => \N__28476\,
            I => \N__28462\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__28473\,
            I => \N__28462\
        );

    \I__6491\ : Span4Mux_v
    port map (
            O => \N__28470\,
            I => \N__28455\
        );

    \I__6490\ : Span4Mux_h
    port map (
            O => \N__28467\,
            I => \N__28455\
        );

    \I__6489\ : Span4Mux_v
    port map (
            O => \N__28462\,
            I => \N__28452\
        );

    \I__6488\ : InMux
    port map (
            O => \N__28461\,
            I => \N__28449\
        );

    \I__6487\ : InMux
    port map (
            O => \N__28460\,
            I => \N__28446\
        );

    \I__6486\ : Span4Mux_h
    port map (
            O => \N__28455\,
            I => \N__28441\
        );

    \I__6485\ : Span4Mux_v
    port map (
            O => \N__28452\,
            I => \N__28436\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__28449\,
            I => \N__28436\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__28446\,
            I => \N__28433\
        );

    \I__6482\ : InMux
    port map (
            O => \N__28445\,
            I => \N__28430\
        );

    \I__6481\ : InMux
    port map (
            O => \N__28444\,
            I => \N__28427\
        );

    \I__6480\ : Span4Mux_h
    port map (
            O => \N__28441\,
            I => \N__28424\
        );

    \I__6479\ : Span4Mux_h
    port map (
            O => \N__28436\,
            I => \N__28421\
        );

    \I__6478\ : Span4Mux_v
    port map (
            O => \N__28433\,
            I => \N__28416\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__28430\,
            I => \N__28416\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__28427\,
            I => \N__28413\
        );

    \I__6475\ : Span4Mux_h
    port map (
            O => \N__28424\,
            I => \N__28404\
        );

    \I__6474\ : Span4Mux_v
    port map (
            O => \N__28421\,
            I => \N__28404\
        );

    \I__6473\ : Span4Mux_h
    port map (
            O => \N__28416\,
            I => \N__28404\
        );

    \I__6472\ : Span4Mux_h
    port map (
            O => \N__28413\,
            I => \N__28404\
        );

    \I__6471\ : Odrv4
    port map (
            O => \N__28404\,
            I => \N_226\
        );

    \I__6470\ : InMux
    port map (
            O => \N__28401\,
            I => \N__28398\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__28398\,
            I => \M_this_data_tmp_qZ0Z_6\
        );

    \I__6468\ : InMux
    port map (
            O => \N__28395\,
            I => \N__28392\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__28392\,
            I => \N__28389\
        );

    \I__6466\ : Span4Mux_h
    port map (
            O => \N__28389\,
            I => \N__28386\
        );

    \I__6465\ : Odrv4
    port map (
            O => \N__28386\,
            I => \M_this_oam_ram_write_data_6\
        );

    \I__6464\ : InMux
    port map (
            O => \N__28383\,
            I => \N__28380\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__28380\,
            I => \N__28377\
        );

    \I__6462\ : Span12Mux_s8_v
    port map (
            O => \N__28377\,
            I => \N__28374\
        );

    \I__6461\ : Odrv12
    port map (
            O => \N__28374\,
            I => \M_this_data_tmp_qZ0Z_2\
        );

    \I__6460\ : InMux
    port map (
            O => \N__28371\,
            I => \N__28368\
        );

    \I__6459\ : LocalMux
    port map (
            O => \N__28368\,
            I => \N__28365\
        );

    \I__6458\ : Span4Mux_v
    port map (
            O => \N__28365\,
            I => \N__28362\
        );

    \I__6457\ : Odrv4
    port map (
            O => \N__28362\,
            I => \M_this_oam_ram_write_data_2\
        );

    \I__6456\ : InMux
    port map (
            O => \N__28359\,
            I => \N__28356\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__28356\,
            I => \M_this_data_tmp_qZ0Z_1\
        );

    \I__6454\ : InMux
    port map (
            O => \N__28353\,
            I => \N__28350\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__28350\,
            I => \N__28347\
        );

    \I__6452\ : Span4Mux_h
    port map (
            O => \N__28347\,
            I => \N__28344\
        );

    \I__6451\ : Odrv4
    port map (
            O => \N__28344\,
            I => \M_this_oam_ram_write_data_1\
        );

    \I__6450\ : InMux
    port map (
            O => \N__28341\,
            I => \M_this_data_count_q_cry_3\
        );

    \I__6449\ : InMux
    port map (
            O => \N__28338\,
            I => \M_this_data_count_q_cry_4\
        );

    \I__6448\ : InMux
    port map (
            O => \N__28335\,
            I => \M_this_data_count_q_cry_5\
        );

    \I__6447\ : InMux
    port map (
            O => \N__28332\,
            I => \M_this_data_count_q_cry_6\
        );

    \I__6446\ : InMux
    port map (
            O => \N__28329\,
            I => \N__28326\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__28326\,
            I => \N__28323\
        );

    \I__6444\ : Odrv4
    port map (
            O => \N__28323\,
            I => \M_this_data_count_q_s_8\
        );

    \I__6443\ : InMux
    port map (
            O => \N__28320\,
            I => \bfn_21_23_0_\
        );

    \I__6442\ : InMux
    port map (
            O => \N__28317\,
            I => \N__28314\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__28314\,
            I => \N__28311\
        );

    \I__6440\ : Span4Mux_v
    port map (
            O => \N__28311\,
            I => \N__28308\
        );

    \I__6439\ : Odrv4
    port map (
            O => \N__28308\,
            I => \M_this_data_count_q_s_9\
        );

    \I__6438\ : InMux
    port map (
            O => \N__28305\,
            I => \M_this_data_count_q_cry_8\
        );

    \I__6437\ : InMux
    port map (
            O => \N__28302\,
            I => \N__28299\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__28299\,
            I => \N__28296\
        );

    \I__6435\ : Odrv12
    port map (
            O => \N__28296\,
            I => \M_this_data_count_q_cry_9_THRU_CO\
        );

    \I__6434\ : InMux
    port map (
            O => \N__28293\,
            I => \M_this_data_count_q_cry_9\
        );

    \I__6433\ : InMux
    port map (
            O => \N__28290\,
            I => \N__28287\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__28287\,
            I => \N__28284\
        );

    \I__6431\ : Odrv4
    port map (
            O => \N__28284\,
            I => \M_this_data_count_q_s_11\
        );

    \I__6430\ : InMux
    port map (
            O => \N__28281\,
            I => \M_this_data_count_q_cry_10\
        );

    \I__6429\ : InMux
    port map (
            O => \N__28278\,
            I => \N__28275\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__28275\,
            I => \N__28272\
        );

    \I__6427\ : Odrv4
    port map (
            O => \N__28272\,
            I => \M_this_data_count_q_s_12\
        );

    \I__6426\ : InMux
    port map (
            O => \N__28269\,
            I => \M_this_data_count_q_cry_11\
        );

    \I__6425\ : InMux
    port map (
            O => \N__28266\,
            I => \N__28246\
        );

    \I__6424\ : InMux
    port map (
            O => \N__28265\,
            I => \N__28246\
        );

    \I__6423\ : InMux
    port map (
            O => \N__28264\,
            I => \N__28246\
        );

    \I__6422\ : InMux
    port map (
            O => \N__28263\,
            I => \N__28246\
        );

    \I__6421\ : InMux
    port map (
            O => \N__28262\,
            I => \N__28246\
        );

    \I__6420\ : InMux
    port map (
            O => \N__28261\,
            I => \N__28246\
        );

    \I__6419\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28241\
        );

    \I__6418\ : InMux
    port map (
            O => \N__28259\,
            I => \N__28241\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__28246\,
            I => \N_755\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__28241\,
            I => \N_755\
        );

    \I__6415\ : InMux
    port map (
            O => \N__28236\,
            I => \M_this_data_count_q_cry_0\
        );

    \I__6414\ : CascadeMux
    port map (
            O => \N__28233\,
            I => \N__28230\
        );

    \I__6413\ : InMux
    port map (
            O => \N__28230\,
            I => \N__28227\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__28227\,
            I => \N__28224\
        );

    \I__6411\ : Odrv4
    port map (
            O => \N__28224\,
            I => \M_this_data_count_q_s_2\
        );

    \I__6410\ : InMux
    port map (
            O => \N__28221\,
            I => \M_this_data_count_q_cry_1\
        );

    \I__6409\ : InMux
    port map (
            O => \N__28218\,
            I => \M_this_data_count_q_cry_2\
        );

    \I__6408\ : InMux
    port map (
            O => \N__28215\,
            I => \N__28212\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__28212\,
            I => \this_vga_signals_M_this_data_count_q_3_0_a3_0_a4_0_2\
        );

    \I__6406\ : CascadeMux
    port map (
            O => \N__28209\,
            I => \this_vga_signals_M_this_data_count_q_3_0_a3_0_a4_0_2_cascade_\
        );

    \I__6405\ : CascadeMux
    port map (
            O => \N__28206\,
            I => \N_307_0_cascade_\
        );

    \I__6404\ : InMux
    port map (
            O => \N__28203\,
            I => \N__28199\
        );

    \I__6403\ : InMux
    port map (
            O => \N__28202\,
            I => \N__28196\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__28199\,
            I => \N__28188\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__28196\,
            I => \N__28185\
        );

    \I__6400\ : InMux
    port map (
            O => \N__28195\,
            I => \N__28180\
        );

    \I__6399\ : InMux
    port map (
            O => \N__28194\,
            I => \N__28180\
        );

    \I__6398\ : InMux
    port map (
            O => \N__28193\,
            I => \N__28177\
        );

    \I__6397\ : InMux
    port map (
            O => \N__28192\,
            I => \N__28174\
        );

    \I__6396\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28171\
        );

    \I__6395\ : Span4Mux_h
    port map (
            O => \N__28188\,
            I => \N__28168\
        );

    \I__6394\ : Span4Mux_v
    port map (
            O => \N__28185\,
            I => \N__28165\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__28180\,
            I => \N__28160\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__28177\,
            I => \N__28160\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__28174\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__28171\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__28168\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__6388\ : Odrv4
    port map (
            O => \N__28165\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__6387\ : Odrv4
    port map (
            O => \N__28160\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__6386\ : CascadeMux
    port map (
            O => \N__28149\,
            I => \this_vga_signals.N_665_1_cascade_\
        );

    \I__6385\ : CascadeMux
    port map (
            O => \N__28146\,
            I => \M_this_data_count_q_3_0_13_cascade_\
        );

    \I__6384\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28140\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__28140\,
            I => this_vga_signals_un20_i_a2_0_a3_0_a4_2_2
        );

    \I__6382\ : InMux
    port map (
            O => \N__28137\,
            I => \N__28134\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__28134\,
            I => \N__28131\
        );

    \I__6380\ : Span4Mux_h
    port map (
            O => \N__28131\,
            I => \N__28128\
        );

    \I__6379\ : Sp12to4
    port map (
            O => \N__28128\,
            I => \N__28125\
        );

    \I__6378\ : Odrv12
    port map (
            O => \N__28125\,
            I => \this_sprites_ram.mem_out_bus5_0\
        );

    \I__6377\ : InMux
    port map (
            O => \N__28122\,
            I => \N__28119\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__28119\,
            I => \N__28116\
        );

    \I__6375\ : Span4Mux_v
    port map (
            O => \N__28116\,
            I => \N__28113\
        );

    \I__6374\ : Odrv4
    port map (
            O => \N__28113\,
            I => \this_sprites_ram.mem_out_bus1_0\
        );

    \I__6373\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28105\
        );

    \I__6372\ : InMux
    port map (
            O => \N__28109\,
            I => \N__28102\
        );

    \I__6371\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28099\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__28105\,
            I => \N__28091\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__28102\,
            I => \N__28083\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__28099\,
            I => \N__28080\
        );

    \I__6367\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28071\
        );

    \I__6366\ : InMux
    port map (
            O => \N__28097\,
            I => \N__28071\
        );

    \I__6365\ : InMux
    port map (
            O => \N__28096\,
            I => \N__28071\
        );

    \I__6364\ : InMux
    port map (
            O => \N__28095\,
            I => \N__28071\
        );

    \I__6363\ : InMux
    port map (
            O => \N__28094\,
            I => \N__28065\
        );

    \I__6362\ : Span4Mux_h
    port map (
            O => \N__28091\,
            I => \N__28062\
        );

    \I__6361\ : InMux
    port map (
            O => \N__28090\,
            I => \N__28053\
        );

    \I__6360\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28053\
        );

    \I__6359\ : InMux
    port map (
            O => \N__28088\,
            I => \N__28053\
        );

    \I__6358\ : InMux
    port map (
            O => \N__28087\,
            I => \N__28053\
        );

    \I__6357\ : InMux
    port map (
            O => \N__28086\,
            I => \N__28050\
        );

    \I__6356\ : Span4Mux_h
    port map (
            O => \N__28083\,
            I => \N__28043\
        );

    \I__6355\ : Span4Mux_v
    port map (
            O => \N__28080\,
            I => \N__28043\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__28071\,
            I => \N__28043\
        );

    \I__6353\ : InMux
    port map (
            O => \N__28070\,
            I => \N__28036\
        );

    \I__6352\ : InMux
    port map (
            O => \N__28069\,
            I => \N__28036\
        );

    \I__6351\ : InMux
    port map (
            O => \N__28068\,
            I => \N__28036\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__28065\,
            I => \N__28033\
        );

    \I__6349\ : Odrv4
    port map (
            O => \N__28062\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__28053\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__28050\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__6346\ : Odrv4
    port map (
            O => \N__28043\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__28036\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__6344\ : Odrv4
    port map (
            O => \N__28033\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__6343\ : InMux
    port map (
            O => \N__28020\,
            I => \N__28017\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__28017\,
            I => \N__28014\
        );

    \I__6341\ : Odrv4
    port map (
            O => \N__28014\,
            I => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\
        );

    \I__6340\ : InMux
    port map (
            O => \N__28011\,
            I => \N__28002\
        );

    \I__6339\ : InMux
    port map (
            O => \N__28010\,
            I => \N__28002\
        );

    \I__6338\ : InMux
    port map (
            O => \N__28009\,
            I => \N__27997\
        );

    \I__6337\ : InMux
    port map (
            O => \N__28008\,
            I => \N__27997\
        );

    \I__6336\ : InMux
    port map (
            O => \N__28007\,
            I => \N__27994\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__28002\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6334\ : LocalMux
    port map (
            O => \N__27997\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__27994\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6332\ : CascadeMux
    port map (
            O => \N__27987\,
            I => \this_vga_signals.N_433_0_cascade_\
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__27984\,
            I => \this_vga_signals.N_442_0_cascade_\
        );

    \I__6330\ : CascadeMux
    port map (
            O => \N__27981\,
            I => \this_vga_signals.N_719_cascade_\
        );

    \I__6329\ : CascadeMux
    port map (
            O => \N__27978\,
            I => \N__27975\
        );

    \I__6328\ : CascadeBuf
    port map (
            O => \N__27975\,
            I => \N__27972\
        );

    \I__6327\ : CascadeMux
    port map (
            O => \N__27972\,
            I => \N__27969\
        );

    \I__6326\ : InMux
    port map (
            O => \N__27969\,
            I => \N__27965\
        );

    \I__6325\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27962\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__27965\,
            I => \N__27959\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__27962\,
            I => \N__27955\
        );

    \I__6322\ : Span4Mux_v
    port map (
            O => \N__27959\,
            I => \N__27952\
        );

    \I__6321\ : CascadeMux
    port map (
            O => \N__27958\,
            I => \N__27949\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__27955\,
            I => \N__27946\
        );

    \I__6319\ : Sp12to4
    port map (
            O => \N__27952\,
            I => \N__27943\
        );

    \I__6318\ : InMux
    port map (
            O => \N__27949\,
            I => \N__27940\
        );

    \I__6317\ : Sp12to4
    port map (
            O => \N__27946\,
            I => \N__27937\
        );

    \I__6316\ : Span12Mux_h
    port map (
            O => \N__27943\,
            I => \N__27934\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__27940\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__6314\ : Odrv12
    port map (
            O => \N__27937\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__6313\ : Odrv12
    port map (
            O => \N__27934\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__6312\ : CascadeMux
    port map (
            O => \N__27927\,
            I => \N__27924\
        );

    \I__6311\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27920\
        );

    \I__6310\ : CascadeMux
    port map (
            O => \N__27923\,
            I => \N__27917\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__27920\,
            I => \N__27914\
        );

    \I__6308\ : InMux
    port map (
            O => \N__27917\,
            I => \N__27911\
        );

    \I__6307\ : Odrv4
    port map (
            O => \N__27914\,
            I => \this_ppu.M_this_ppu_map_addr_i_9\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__27911\,
            I => \this_ppu.M_this_ppu_map_addr_i_9\
        );

    \I__6305\ : InMux
    port map (
            O => \N__27906\,
            I => \bfn_21_7_0_\
        );

    \I__6304\ : InMux
    port map (
            O => \N__27903\,
            I => \N__27900\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__27900\,
            I => \N__27897\
        );

    \I__6302\ : Odrv4
    port map (
            O => \N__27897\,
            I => \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO\
        );

    \I__6301\ : InMux
    port map (
            O => \N__27894\,
            I => \N__27891\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__27891\,
            I => \N__27888\
        );

    \I__6299\ : Span4Mux_h
    port map (
            O => \N__27888\,
            I => \N__27885\
        );

    \I__6298\ : Odrv4
    port map (
            O => \N__27885\,
            I => \M_this_oam_ram_write_data_16\
        );

    \I__6297\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27879\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__27879\,
            I => \M_this_oam_ram_read_data_i_19\
        );

    \I__6295\ : InMux
    port map (
            O => \N__27876\,
            I => \N__27873\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__27873\,
            I => \M_this_data_tmp_qZ0Z_16\
        );

    \I__6293\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27865\
        );

    \I__6292\ : InMux
    port map (
            O => \N__27869\,
            I => \N__27861\
        );

    \I__6291\ : InMux
    port map (
            O => \N__27868\,
            I => \N__27858\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__27865\,
            I => \N__27855\
        );

    \I__6289\ : InMux
    port map (
            O => \N__27864\,
            I => \N__27852\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__27861\,
            I => \N__27849\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__27858\,
            I => \N__27846\
        );

    \I__6286\ : Span4Mux_h
    port map (
            O => \N__27855\,
            I => \N__27841\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__27852\,
            I => \N__27841\
        );

    \I__6284\ : Span4Mux_v
    port map (
            O => \N__27849\,
            I => \N__27836\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__27846\,
            I => \N__27836\
        );

    \I__6282\ : Span4Mux_h
    port map (
            O => \N__27841\,
            I => \N__27833\
        );

    \I__6281\ : Span4Mux_h
    port map (
            O => \N__27836\,
            I => \N__27830\
        );

    \I__6280\ : Odrv4
    port map (
            O => \N__27833\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__27830\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__6278\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27820\
        );

    \I__6277\ : CascadeMux
    port map (
            O => \N__27824\,
            I => \N__27817\
        );

    \I__6276\ : CascadeMux
    port map (
            O => \N__27823\,
            I => \N__27812\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__27820\,
            I => \N__27809\
        );

    \I__6274\ : InMux
    port map (
            O => \N__27817\,
            I => \N__27806\
        );

    \I__6273\ : InMux
    port map (
            O => \N__27816\,
            I => \N__27803\
        );

    \I__6272\ : InMux
    port map (
            O => \N__27815\,
            I => \N__27799\
        );

    \I__6271\ : InMux
    port map (
            O => \N__27812\,
            I => \N__27796\
        );

    \I__6270\ : Span4Mux_h
    port map (
            O => \N__27809\,
            I => \N__27793\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__27806\,
            I => \N__27790\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__27803\,
            I => \N__27784\
        );

    \I__6267\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27781\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__27799\,
            I => \N__27778\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__27796\,
            I => \N__27773\
        );

    \I__6264\ : Span4Mux_v
    port map (
            O => \N__27793\,
            I => \N__27773\
        );

    \I__6263\ : Span12Mux_v
    port map (
            O => \N__27790\,
            I => \N__27770\
        );

    \I__6262\ : InMux
    port map (
            O => \N__27789\,
            I => \N__27767\
        );

    \I__6261\ : InMux
    port map (
            O => \N__27788\,
            I => \N__27762\
        );

    \I__6260\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27762\
        );

    \I__6259\ : Span4Mux_h
    port map (
            O => \N__27784\,
            I => \N__27759\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__27781\,
            I => \N__27756\
        );

    \I__6257\ : Span4Mux_h
    port map (
            O => \N__27778\,
            I => \N__27751\
        );

    \I__6256\ : Span4Mux_v
    port map (
            O => \N__27773\,
            I => \N__27751\
        );

    \I__6255\ : Odrv12
    port map (
            O => \N__27770\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__27767\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__27762\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__6252\ : Odrv4
    port map (
            O => \N__27759\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__6251\ : Odrv4
    port map (
            O => \N__27756\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__6250\ : Odrv4
    port map (
            O => \N__27751\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__6249\ : CascadeMux
    port map (
            O => \N__27738\,
            I => \N__27734\
        );

    \I__6248\ : CascadeMux
    port map (
            O => \N__27737\,
            I => \N__27731\
        );

    \I__6247\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27728\
        );

    \I__6246\ : InMux
    port map (
            O => \N__27731\,
            I => \N__27725\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__27728\,
            I => \this_ppu.M_this_ppu_vram_addr_i_7\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__27725\,
            I => \this_ppu.M_this_ppu_vram_addr_i_7\
        );

    \I__6243\ : CascadeMux
    port map (
            O => \N__27720\,
            I => \N__27717\
        );

    \I__6242\ : InMux
    port map (
            O => \N__27717\,
            I => \N__27710\
        );

    \I__6241\ : InMux
    port map (
            O => \N__27716\,
            I => \N__27707\
        );

    \I__6240\ : CascadeMux
    port map (
            O => \N__27715\,
            I => \N__27704\
        );

    \I__6239\ : InMux
    port map (
            O => \N__27714\,
            I => \N__27700\
        );

    \I__6238\ : InMux
    port map (
            O => \N__27713\,
            I => \N__27697\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__27710\,
            I => \N__27694\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__27707\,
            I => \N__27691\
        );

    \I__6235\ : InMux
    port map (
            O => \N__27704\,
            I => \N__27688\
        );

    \I__6234\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27685\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__27700\,
            I => \N__27682\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__27697\,
            I => \N__27679\
        );

    \I__6231\ : Span4Mux_v
    port map (
            O => \N__27694\,
            I => \N__27676\
        );

    \I__6230\ : Span12Mux_h
    port map (
            O => \N__27691\,
            I => \N__27673\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__27688\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__27685\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__6227\ : Odrv4
    port map (
            O => \N__27682\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__6226\ : Odrv4
    port map (
            O => \N__27679\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__6225\ : Odrv4
    port map (
            O => \N__27676\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__6224\ : Odrv12
    port map (
            O => \N__27673\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__6223\ : InMux
    port map (
            O => \N__27660\,
            I => \N__27656\
        );

    \I__6222\ : InMux
    port map (
            O => \N__27659\,
            I => \N__27652\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__27656\,
            I => \N__27649\
        );

    \I__6220\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27646\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__27652\,
            I => \N__27643\
        );

    \I__6218\ : Span4Mux_h
    port map (
            O => \N__27649\,
            I => \N__27638\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__27646\,
            I => \N__27638\
        );

    \I__6216\ : Span4Mux_h
    port map (
            O => \N__27643\,
            I => \N__27635\
        );

    \I__6215\ : Span4Mux_h
    port map (
            O => \N__27638\,
            I => \N__27632\
        );

    \I__6214\ : Span4Mux_h
    port map (
            O => \N__27635\,
            I => \N__27629\
        );

    \I__6213\ : Odrv4
    port map (
            O => \N__27632\,
            I => \M_this_oam_ram_read_data_17\
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__27629\,
            I => \M_this_oam_ram_read_data_17\
        );

    \I__6211\ : CascadeMux
    port map (
            O => \N__27624\,
            I => \N__27620\
        );

    \I__6210\ : CascadeMux
    port map (
            O => \N__27623\,
            I => \N__27617\
        );

    \I__6209\ : InMux
    port map (
            O => \N__27620\,
            I => \N__27614\
        );

    \I__6208\ : InMux
    port map (
            O => \N__27617\,
            I => \N__27611\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__27614\,
            I => \this_ppu.M_vaddress_q_i_1\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__27611\,
            I => \this_ppu.M_vaddress_q_i_1\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__27606\,
            I => \N__27598\
        );

    \I__6204\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27595\
        );

    \I__6203\ : InMux
    port map (
            O => \N__27604\,
            I => \N__27592\
        );

    \I__6202\ : InMux
    port map (
            O => \N__27603\,
            I => \N__27589\
        );

    \I__6201\ : CascadeMux
    port map (
            O => \N__27602\,
            I => \N__27586\
        );

    \I__6200\ : InMux
    port map (
            O => \N__27601\,
            I => \N__27580\
        );

    \I__6199\ : InMux
    port map (
            O => \N__27598\,
            I => \N__27580\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__27595\,
            I => \N__27577\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__27592\,
            I => \N__27574\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__27589\,
            I => \N__27571\
        );

    \I__6195\ : InMux
    port map (
            O => \N__27586\,
            I => \N__27568\
        );

    \I__6194\ : InMux
    port map (
            O => \N__27585\,
            I => \N__27565\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__27580\,
            I => \N__27562\
        );

    \I__6192\ : Span4Mux_h
    port map (
            O => \N__27577\,
            I => \N__27557\
        );

    \I__6191\ : Span4Mux_h
    port map (
            O => \N__27574\,
            I => \N__27557\
        );

    \I__6190\ : Span12Mux_v
    port map (
            O => \N__27571\,
            I => \N__27554\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__27568\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__27565\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__6187\ : Odrv4
    port map (
            O => \N__27562\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__6186\ : Odrv4
    port map (
            O => \N__27557\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__6185\ : Odrv12
    port map (
            O => \N__27554\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__6184\ : CascadeMux
    port map (
            O => \N__27543\,
            I => \N__27540\
        );

    \I__6183\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27535\
        );

    \I__6182\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27532\
        );

    \I__6181\ : CascadeMux
    port map (
            O => \N__27538\,
            I => \N__27529\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__27535\,
            I => \N__27526\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__27532\,
            I => \N__27523\
        );

    \I__6178\ : InMux
    port map (
            O => \N__27529\,
            I => \N__27520\
        );

    \I__6177\ : Span4Mux_v
    port map (
            O => \N__27526\,
            I => \N__27517\
        );

    \I__6176\ : Span4Mux_v
    port map (
            O => \N__27523\,
            I => \N__27514\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__27520\,
            I => \N__27511\
        );

    \I__6174\ : Span4Mux_h
    port map (
            O => \N__27517\,
            I => \N__27508\
        );

    \I__6173\ : Span4Mux_h
    port map (
            O => \N__27514\,
            I => \N__27503\
        );

    \I__6172\ : Span4Mux_v
    port map (
            O => \N__27511\,
            I => \N__27503\
        );

    \I__6171\ : Odrv4
    port map (
            O => \N__27508\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__6170\ : Odrv4
    port map (
            O => \N__27503\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__6169\ : InMux
    port map (
            O => \N__27498\,
            I => \N__27494\
        );

    \I__6168\ : InMux
    port map (
            O => \N__27497\,
            I => \N__27491\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__27494\,
            I => \this_ppu.M_vaddress_q_i_2\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__27491\,
            I => \this_ppu.M_vaddress_q_i_2\
        );

    \I__6165\ : CascadeMux
    port map (
            O => \N__27486\,
            I => \N__27483\
        );

    \I__6164\ : CascadeBuf
    port map (
            O => \N__27483\,
            I => \N__27480\
        );

    \I__6163\ : CascadeMux
    port map (
            O => \N__27480\,
            I => \N__27477\
        );

    \I__6162\ : InMux
    port map (
            O => \N__27477\,
            I => \N__27473\
        );

    \I__6161\ : InMux
    port map (
            O => \N__27476\,
            I => \N__27469\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__27473\,
            I => \N__27466\
        );

    \I__6159\ : InMux
    port map (
            O => \N__27472\,
            I => \N__27463\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__27469\,
            I => \N__27458\
        );

    \I__6157\ : Sp12to4
    port map (
            O => \N__27466\,
            I => \N__27455\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__27463\,
            I => \N__27452\
        );

    \I__6155\ : InMux
    port map (
            O => \N__27462\,
            I => \N__27447\
        );

    \I__6154\ : InMux
    port map (
            O => \N__27461\,
            I => \N__27447\
        );

    \I__6153\ : Span12Mux_v
    port map (
            O => \N__27458\,
            I => \N__27442\
        );

    \I__6152\ : Span12Mux_v
    port map (
            O => \N__27455\,
            I => \N__27442\
        );

    \I__6151\ : Odrv4
    port map (
            O => \N__27452\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__27447\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__6149\ : Odrv12
    port map (
            O => \N__27442\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__6148\ : CascadeMux
    port map (
            O => \N__27435\,
            I => \N__27431\
        );

    \I__6147\ : CascadeMux
    port map (
            O => \N__27434\,
            I => \N__27428\
        );

    \I__6146\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27425\
        );

    \I__6145\ : InMux
    port map (
            O => \N__27428\,
            I => \N__27422\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__27425\,
            I => \this_ppu.M_this_ppu_map_addr_i_5\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__27422\,
            I => \this_ppu.M_this_ppu_map_addr_i_5\
        );

    \I__6142\ : CascadeMux
    port map (
            O => \N__27417\,
            I => \N__27414\
        );

    \I__6141\ : CascadeBuf
    port map (
            O => \N__27414\,
            I => \N__27411\
        );

    \I__6140\ : CascadeMux
    port map (
            O => \N__27411\,
            I => \N__27408\
        );

    \I__6139\ : InMux
    port map (
            O => \N__27408\,
            I => \N__27405\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__27405\,
            I => \N__27401\
        );

    \I__6137\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27396\
        );

    \I__6136\ : Span4Mux_v
    port map (
            O => \N__27401\,
            I => \N__27393\
        );

    \I__6135\ : CascadeMux
    port map (
            O => \N__27400\,
            I => \N__27390\
        );

    \I__6134\ : InMux
    port map (
            O => \N__27399\,
            I => \N__27387\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__27396\,
            I => \N__27384\
        );

    \I__6132\ : Sp12to4
    port map (
            O => \N__27393\,
            I => \N__27381\
        );

    \I__6131\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27378\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__27387\,
            I => \N__27375\
        );

    \I__6129\ : Span12Mux_v
    port map (
            O => \N__27384\,
            I => \N__27370\
        );

    \I__6128\ : Span12Mux_v
    port map (
            O => \N__27381\,
            I => \N__27370\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__27378\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__6126\ : Odrv4
    port map (
            O => \N__27375\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__6125\ : Odrv12
    port map (
            O => \N__27370\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__6124\ : CascadeMux
    port map (
            O => \N__27363\,
            I => \N__27359\
        );

    \I__6123\ : CascadeMux
    port map (
            O => \N__27362\,
            I => \N__27356\
        );

    \I__6122\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27353\
        );

    \I__6121\ : InMux
    port map (
            O => \N__27356\,
            I => \N__27350\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__27353\,
            I => \N__27347\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__27350\,
            I => \this_ppu.M_this_ppu_map_addr_i_6\
        );

    \I__6118\ : Odrv4
    port map (
            O => \N__27347\,
            I => \this_ppu.M_this_ppu_map_addr_i_6\
        );

    \I__6117\ : CascadeMux
    port map (
            O => \N__27342\,
            I => \N__27339\
        );

    \I__6116\ : CascadeBuf
    port map (
            O => \N__27339\,
            I => \N__27336\
        );

    \I__6115\ : CascadeMux
    port map (
            O => \N__27336\,
            I => \N__27332\
        );

    \I__6114\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27329\
        );

    \I__6113\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27326\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__27329\,
            I => \N__27323\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__27326\,
            I => \N__27320\
        );

    \I__6110\ : Span4Mux_h
    port map (
            O => \N__27323\,
            I => \N__27314\
        );

    \I__6109\ : Span12Mux_h
    port map (
            O => \N__27320\,
            I => \N__27311\
        );

    \I__6108\ : InMux
    port map (
            O => \N__27319\,
            I => \N__27308\
        );

    \I__6107\ : InMux
    port map (
            O => \N__27318\,
            I => \N__27303\
        );

    \I__6106\ : InMux
    port map (
            O => \N__27317\,
            I => \N__27303\
        );

    \I__6105\ : Sp12to4
    port map (
            O => \N__27314\,
            I => \N__27298\
        );

    \I__6104\ : Span12Mux_v
    port map (
            O => \N__27311\,
            I => \N__27298\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__27308\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__27303\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__6101\ : Odrv12
    port map (
            O => \N__27298\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__27291\,
            I => \N__27287\
        );

    \I__6099\ : InMux
    port map (
            O => \N__27290\,
            I => \N__27284\
        );

    \I__6098\ : InMux
    port map (
            O => \N__27287\,
            I => \N__27281\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__27284\,
            I => \this_ppu.M_this_ppu_map_addr_i_7\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__27281\,
            I => \this_ppu.M_this_ppu_map_addr_i_7\
        );

    \I__6095\ : CascadeMux
    port map (
            O => \N__27276\,
            I => \N__27273\
        );

    \I__6094\ : CascadeBuf
    port map (
            O => \N__27273\,
            I => \N__27269\
        );

    \I__6093\ : InMux
    port map (
            O => \N__27272\,
            I => \N__27266\
        );

    \I__6092\ : CascadeMux
    port map (
            O => \N__27269\,
            I => \N__27263\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__27266\,
            I => \N__27260\
        );

    \I__6090\ : InMux
    port map (
            O => \N__27263\,
            I => \N__27257\
        );

    \I__6089\ : Span4Mux_h
    port map (
            O => \N__27260\,
            I => \N__27254\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__27257\,
            I => \N__27251\
        );

    \I__6087\ : Span4Mux_v
    port map (
            O => \N__27254\,
            I => \N__27246\
        );

    \I__6086\ : Span12Mux_s5_v
    port map (
            O => \N__27251\,
            I => \N__27243\
        );

    \I__6085\ : InMux
    port map (
            O => \N__27250\,
            I => \N__27240\
        );

    \I__6084\ : InMux
    port map (
            O => \N__27249\,
            I => \N__27237\
        );

    \I__6083\ : Span4Mux_v
    port map (
            O => \N__27246\,
            I => \N__27234\
        );

    \I__6082\ : Span12Mux_v
    port map (
            O => \N__27243\,
            I => \N__27231\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__27240\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__27237\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__6079\ : Odrv4
    port map (
            O => \N__27234\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__6078\ : Odrv12
    port map (
            O => \N__27231\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__6077\ : CascadeMux
    port map (
            O => \N__27222\,
            I => \N__27218\
        );

    \I__6076\ : CascadeMux
    port map (
            O => \N__27221\,
            I => \N__27215\
        );

    \I__6075\ : InMux
    port map (
            O => \N__27218\,
            I => \N__27212\
        );

    \I__6074\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27209\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__27212\,
            I => \this_ppu.M_this_ppu_map_addr_i_8\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__27209\,
            I => \this_ppu.M_this_ppu_map_addr_i_8\
        );

    \I__6071\ : CascadeMux
    port map (
            O => \N__27204\,
            I => \N__27201\
        );

    \I__6070\ : InMux
    port map (
            O => \N__27201\,
            I => \N__27198\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__27198\,
            I => \N__27194\
        );

    \I__6068\ : CascadeMux
    port map (
            O => \N__27197\,
            I => \N__27191\
        );

    \I__6067\ : Span4Mux_v
    port map (
            O => \N__27194\,
            I => \N__27188\
        );

    \I__6066\ : InMux
    port map (
            O => \N__27191\,
            I => \N__27185\
        );

    \I__6065\ : Odrv4
    port map (
            O => \N__27188\,
            I => \N_460_0\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__27185\,
            I => \N_460_0\
        );

    \I__6063\ : CascadeMux
    port map (
            O => \N__27180\,
            I => \N__27176\
        );

    \I__6062\ : InMux
    port map (
            O => \N__27179\,
            I => \N__27173\
        );

    \I__6061\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27170\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__27173\,
            I => \N__27165\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__27170\,
            I => \N__27162\
        );

    \I__6058\ : InMux
    port map (
            O => \N__27169\,
            I => \N__27155\
        );

    \I__6057\ : InMux
    port map (
            O => \N__27168\,
            I => \N__27155\
        );

    \I__6056\ : Span4Mux_v
    port map (
            O => \N__27165\,
            I => \N__27151\
        );

    \I__6055\ : Span4Mux_v
    port map (
            O => \N__27162\,
            I => \N__27148\
        );

    \I__6054\ : InMux
    port map (
            O => \N__27161\,
            I => \N__27143\
        );

    \I__6053\ : InMux
    port map (
            O => \N__27160\,
            I => \N__27143\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__27155\,
            I => \N__27140\
        );

    \I__6051\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27137\
        );

    \I__6050\ : Odrv4
    port map (
            O => \N__27151\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6049\ : Odrv4
    port map (
            O => \N__27148\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__27143\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6047\ : Odrv12
    port map (
            O => \N__27140\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__27137\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6045\ : InMux
    port map (
            O => \N__27126\,
            I => \N__27118\
        );

    \I__6044\ : InMux
    port map (
            O => \N__27125\,
            I => \N__27118\
        );

    \I__6043\ : InMux
    port map (
            O => \N__27124\,
            I => \N__27115\
        );

    \I__6042\ : InMux
    port map (
            O => \N__27123\,
            I => \N__27112\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__27118\,
            I => \N__27107\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__27115\,
            I => \N__27102\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__27112\,
            I => \N__27102\
        );

    \I__6038\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27097\
        );

    \I__6037\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27097\
        );

    \I__6036\ : Odrv4
    port map (
            O => \N__27107\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__6035\ : Odrv12
    port map (
            O => \N__27102\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__27097\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__6033\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27087\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__27087\,
            I => \N__27084\
        );

    \I__6031\ : Odrv4
    port map (
            O => \N__27084\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0Z0Z_2\
        );

    \I__6030\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27077\
        );

    \I__6029\ : InMux
    port map (
            O => \N__27080\,
            I => \N__27074\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__27077\,
            I => \N__27068\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__27074\,
            I => \N__27068\
        );

    \I__6026\ : InMux
    port map (
            O => \N__27073\,
            I => \N__27065\
        );

    \I__6025\ : Span4Mux_h
    port map (
            O => \N__27068\,
            I => \N__27062\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__27065\,
            I => \N__27059\
        );

    \I__6023\ : Odrv4
    port map (
            O => \N__27062\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a2Z0Z_1\
        );

    \I__6022\ : Odrv4
    port map (
            O => \N__27059\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a2Z0Z_1\
        );

    \I__6021\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27039\
        );

    \I__6020\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27033\
        );

    \I__6019\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27026\
        );

    \I__6018\ : InMux
    port map (
            O => \N__27051\,
            I => \N__27026\
        );

    \I__6017\ : InMux
    port map (
            O => \N__27050\,
            I => \N__27026\
        );

    \I__6016\ : InMux
    port map (
            O => \N__27049\,
            I => \N__27023\
        );

    \I__6015\ : InMux
    port map (
            O => \N__27048\,
            I => \N__27018\
        );

    \I__6014\ : InMux
    port map (
            O => \N__27047\,
            I => \N__27018\
        );

    \I__6013\ : InMux
    port map (
            O => \N__27046\,
            I => \N__27011\
        );

    \I__6012\ : InMux
    port map (
            O => \N__27045\,
            I => \N__27011\
        );

    \I__6011\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27008\
        );

    \I__6010\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27002\
        );

    \I__6009\ : InMux
    port map (
            O => \N__27042\,
            I => \N__26999\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__27039\,
            I => \N__26996\
        );

    \I__6007\ : InMux
    port map (
            O => \N__27038\,
            I => \N__26993\
        );

    \I__6006\ : InMux
    port map (
            O => \N__27037\,
            I => \N__26990\
        );

    \I__6005\ : CascadeMux
    port map (
            O => \N__27036\,
            I => \N__26986\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__27033\,
            I => \N__26980\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__27026\,
            I => \N__26980\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__27023\,
            I => \N__26975\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__27018\,
            I => \N__26975\
        );

    \I__6000\ : InMux
    port map (
            O => \N__27017\,
            I => \N__26970\
        );

    \I__5999\ : InMux
    port map (
            O => \N__27016\,
            I => \N__26970\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__27011\,
            I => \N__26965\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__27008\,
            I => \N__26965\
        );

    \I__5996\ : InMux
    port map (
            O => \N__27007\,
            I => \N__26960\
        );

    \I__5995\ : InMux
    port map (
            O => \N__27006\,
            I => \N__26960\
        );

    \I__5994\ : InMux
    port map (
            O => \N__27005\,
            I => \N__26957\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__27002\,
            I => \N__26954\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__26999\,
            I => \N__26951\
        );

    \I__5991\ : Span4Mux_v
    port map (
            O => \N__26996\,
            I => \N__26946\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__26993\,
            I => \N__26946\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__26990\,
            I => \N__26943\
        );

    \I__5988\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26936\
        );

    \I__5987\ : InMux
    port map (
            O => \N__26986\,
            I => \N__26931\
        );

    \I__5986\ : InMux
    port map (
            O => \N__26985\,
            I => \N__26931\
        );

    \I__5985\ : Span4Mux_h
    port map (
            O => \N__26980\,
            I => \N__26920\
        );

    \I__5984\ : Span4Mux_v
    port map (
            O => \N__26975\,
            I => \N__26920\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__26970\,
            I => \N__26920\
        );

    \I__5982\ : Span4Mux_v
    port map (
            O => \N__26965\,
            I => \N__26920\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__26960\,
            I => \N__26920\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__26957\,
            I => \N__26915\
        );

    \I__5979\ : Span4Mux_h
    port map (
            O => \N__26954\,
            I => \N__26915\
        );

    \I__5978\ : Span4Mux_v
    port map (
            O => \N__26951\,
            I => \N__26910\
        );

    \I__5977\ : Span4Mux_h
    port map (
            O => \N__26946\,
            I => \N__26910\
        );

    \I__5976\ : Span12Mux_v
    port map (
            O => \N__26943\,
            I => \N__26907\
        );

    \I__5975\ : InMux
    port map (
            O => \N__26942\,
            I => \N__26898\
        );

    \I__5974\ : InMux
    port map (
            O => \N__26941\,
            I => \N__26898\
        );

    \I__5973\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26898\
        );

    \I__5972\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26898\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__26936\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__26931\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5969\ : Odrv4
    port map (
            O => \N__26920\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5968\ : Odrv4
    port map (
            O => \N__26915\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5967\ : Odrv4
    port map (
            O => \N__26910\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5966\ : Odrv12
    port map (
            O => \N__26907\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__26898\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__5964\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26880\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__26880\,
            I => \N__26874\
        );

    \I__5962\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26871\
        );

    \I__5961\ : InMux
    port map (
            O => \N__26878\,
            I => \N__26868\
        );

    \I__5960\ : InMux
    port map (
            O => \N__26877\,
            I => \N__26865\
        );

    \I__5959\ : Span4Mux_v
    port map (
            O => \N__26874\,
            I => \N__26860\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__26871\,
            I => \N__26860\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__26868\,
            I => \N__26857\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__26865\,
            I => \N__26850\
        );

    \I__5955\ : Span4Mux_v
    port map (
            O => \N__26860\,
            I => \N__26845\
        );

    \I__5954\ : Span4Mux_h
    port map (
            O => \N__26857\,
            I => \N__26845\
        );

    \I__5953\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26842\
        );

    \I__5952\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26839\
        );

    \I__5951\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26836\
        );

    \I__5950\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26833\
        );

    \I__5949\ : Span4Mux_s3_v
    port map (
            O => \N__26850\,
            I => \N__26830\
        );

    \I__5948\ : Span4Mux_v
    port map (
            O => \N__26845\,
            I => \N__26827\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__26842\,
            I => \N__26824\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__26839\,
            I => \N__26821\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__26836\,
            I => \N__26818\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__26833\,
            I => \N__26815\
        );

    \I__5943\ : Span4Mux_v
    port map (
            O => \N__26830\,
            I => \N__26808\
        );

    \I__5942\ : Span4Mux_v
    port map (
            O => \N__26827\,
            I => \N__26808\
        );

    \I__5941\ : Span4Mux_h
    port map (
            O => \N__26824\,
            I => \N__26808\
        );

    \I__5940\ : Span12Mux_h
    port map (
            O => \N__26821\,
            I => \N__26805\
        );

    \I__5939\ : Span12Mux_h
    port map (
            O => \N__26818\,
            I => \N__26800\
        );

    \I__5938\ : Span12Mux_h
    port map (
            O => \N__26815\,
            I => \N__26800\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__26808\,
            I => \N__26797\
        );

    \I__5936\ : Odrv12
    port map (
            O => \N__26805\,
            I => \N_250\
        );

    \I__5935\ : Odrv12
    port map (
            O => \N__26800\,
            I => \N_250\
        );

    \I__5934\ : Odrv4
    port map (
            O => \N__26797\,
            I => \N_250\
        );

    \I__5933\ : CascadeMux
    port map (
            O => \N__26790\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_3Z0Z_0_cascade_\
        );

    \I__5932\ : CascadeMux
    port map (
            O => \N__26787\,
            I => \N__26784\
        );

    \I__5931\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26780\
        );

    \I__5930\ : CascadeMux
    port map (
            O => \N__26783\,
            I => \N__26777\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__26780\,
            I => \N__26772\
        );

    \I__5928\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26765\
        );

    \I__5927\ : InMux
    port map (
            O => \N__26776\,
            I => \N__26765\
        );

    \I__5926\ : InMux
    port map (
            O => \N__26775\,
            I => \N__26765\
        );

    \I__5925\ : Span4Mux_h
    port map (
            O => \N__26772\,
            I => \N__26762\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__26765\,
            I => \N__26759\
        );

    \I__5923\ : Odrv4
    port map (
            O => \N__26762\,
            I => \this_vga_signals.N_743\
        );

    \I__5922\ : Odrv12
    port map (
            O => \N__26759\,
            I => \this_vga_signals.N_743\
        );

    \I__5921\ : InMux
    port map (
            O => \N__26754\,
            I => \N__26750\
        );

    \I__5920\ : InMux
    port map (
            O => \N__26753\,
            I => \N__26741\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__26750\,
            I => \N__26738\
        );

    \I__5918\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26735\
        );

    \I__5917\ : InMux
    port map (
            O => \N__26748\,
            I => \N__26732\
        );

    \I__5916\ : InMux
    port map (
            O => \N__26747\,
            I => \N__26729\
        );

    \I__5915\ : InMux
    port map (
            O => \N__26746\,
            I => \N__26726\
        );

    \I__5914\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26723\
        );

    \I__5913\ : InMux
    port map (
            O => \N__26744\,
            I => \N__26720\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__26741\,
            I => \N__26717\
        );

    \I__5911\ : Span4Mux_v
    port map (
            O => \N__26738\,
            I => \N__26714\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__26735\,
            I => \N__26709\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__26732\,
            I => \N__26709\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__26729\,
            I => \N__26706\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__26726\,
            I => \N__26703\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__26723\,
            I => \N__26698\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__26720\,
            I => \N__26698\
        );

    \I__5904\ : Span4Mux_v
    port map (
            O => \N__26717\,
            I => \N__26693\
        );

    \I__5903\ : Span4Mux_v
    port map (
            O => \N__26714\,
            I => \N__26693\
        );

    \I__5902\ : Span4Mux_v
    port map (
            O => \N__26709\,
            I => \N__26690\
        );

    \I__5901\ : Span4Mux_v
    port map (
            O => \N__26706\,
            I => \N__26685\
        );

    \I__5900\ : Span4Mux_v
    port map (
            O => \N__26703\,
            I => \N__26685\
        );

    \I__5899\ : Span12Mux_v
    port map (
            O => \N__26698\,
            I => \N__26682\
        );

    \I__5898\ : Sp12to4
    port map (
            O => \N__26693\,
            I => \N__26679\
        );

    \I__5897\ : Span4Mux_h
    port map (
            O => \N__26690\,
            I => \N__26674\
        );

    \I__5896\ : Span4Mux_h
    port map (
            O => \N__26685\,
            I => \N__26674\
        );

    \I__5895\ : Span12Mux_h
    port map (
            O => \N__26682\,
            I => \N__26669\
        );

    \I__5894\ : Span12Mux_h
    port map (
            O => \N__26679\,
            I => \N__26669\
        );

    \I__5893\ : Odrv4
    port map (
            O => \N__26674\,
            I => \N_228\
        );

    \I__5892\ : Odrv12
    port map (
            O => \N__26669\,
            I => \N_228\
        );

    \I__5891\ : InMux
    port map (
            O => \N__26664\,
            I => \N__26657\
        );

    \I__5890\ : InMux
    port map (
            O => \N__26663\,
            I => \N__26654\
        );

    \I__5889\ : InMux
    port map (
            O => \N__26662\,
            I => \N__26648\
        );

    \I__5888\ : InMux
    port map (
            O => \N__26661\,
            I => \N__26645\
        );

    \I__5887\ : InMux
    port map (
            O => \N__26660\,
            I => \N__26642\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__26657\,
            I => \N__26639\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__26654\,
            I => \N__26636\
        );

    \I__5884\ : InMux
    port map (
            O => \N__26653\,
            I => \N__26633\
        );

    \I__5883\ : InMux
    port map (
            O => \N__26652\,
            I => \N__26630\
        );

    \I__5882\ : InMux
    port map (
            O => \N__26651\,
            I => \N__26627\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__26648\,
            I => \N__26624\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__26645\,
            I => \N__26621\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__26642\,
            I => \N__26618\
        );

    \I__5878\ : Span4Mux_v
    port map (
            O => \N__26639\,
            I => \N__26613\
        );

    \I__5877\ : Span4Mux_v
    port map (
            O => \N__26636\,
            I => \N__26613\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__26633\,
            I => \N__26610\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__26630\,
            I => \N__26607\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__26627\,
            I => \N__26604\
        );

    \I__5873\ : Span4Mux_v
    port map (
            O => \N__26624\,
            I => \N__26599\
        );

    \I__5872\ : Span4Mux_h
    port map (
            O => \N__26621\,
            I => \N__26599\
        );

    \I__5871\ : Span4Mux_s2_v
    port map (
            O => \N__26618\,
            I => \N__26596\
        );

    \I__5870\ : Span4Mux_h
    port map (
            O => \N__26613\,
            I => \N__26593\
        );

    \I__5869\ : Span12Mux_s9_h
    port map (
            O => \N__26610\,
            I => \N__26590\
        );

    \I__5868\ : Span4Mux_h
    port map (
            O => \N__26607\,
            I => \N__26583\
        );

    \I__5867\ : Span4Mux_v
    port map (
            O => \N__26604\,
            I => \N__26583\
        );

    \I__5866\ : Span4Mux_v
    port map (
            O => \N__26599\,
            I => \N__26583\
        );

    \I__5865\ : Span4Mux_h
    port map (
            O => \N__26596\,
            I => \N__26580\
        );

    \I__5864\ : Span4Mux_h
    port map (
            O => \N__26593\,
            I => \N__26577\
        );

    \I__5863\ : Span12Mux_v
    port map (
            O => \N__26590\,
            I => \N__26574\
        );

    \I__5862\ : Span4Mux_h
    port map (
            O => \N__26583\,
            I => \N__26569\
        );

    \I__5861\ : Span4Mux_v
    port map (
            O => \N__26580\,
            I => \N__26569\
        );

    \I__5860\ : Odrv4
    port map (
            O => \N__26577\,
            I => \N_248\
        );

    \I__5859\ : Odrv12
    port map (
            O => \N__26574\,
            I => \N_248\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__26569\,
            I => \N_248\
        );

    \I__5857\ : InMux
    port map (
            O => \N__26562\,
            I => \N__26559\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__26559\,
            I => \M_this_sprites_address_qc_12_0\
        );

    \I__5855\ : InMux
    port map (
            O => \N__26556\,
            I => \N__26545\
        );

    \I__5854\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26542\
        );

    \I__5853\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26539\
        );

    \I__5852\ : InMux
    port map (
            O => \N__26553\,
            I => \N__26533\
        );

    \I__5851\ : CascadeMux
    port map (
            O => \N__26552\,
            I => \N__26530\
        );

    \I__5850\ : InMux
    port map (
            O => \N__26551\,
            I => \N__26523\
        );

    \I__5849\ : InMux
    port map (
            O => \N__26550\,
            I => \N__26523\
        );

    \I__5848\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26523\
        );

    \I__5847\ : InMux
    port map (
            O => \N__26548\,
            I => \N__26520\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__26545\,
            I => \N__26515\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__26542\,
            I => \N__26510\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__26539\,
            I => \N__26510\
        );

    \I__5843\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26506\
        );

    \I__5842\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26501\
        );

    \I__5841\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26501\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__26533\,
            I => \N__26498\
        );

    \I__5839\ : InMux
    port map (
            O => \N__26530\,
            I => \N__26495\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__26523\,
            I => \N__26492\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__26520\,
            I => \N__26489\
        );

    \I__5836\ : InMux
    port map (
            O => \N__26519\,
            I => \N__26486\
        );

    \I__5835\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26483\
        );

    \I__5834\ : Span4Mux_h
    port map (
            O => \N__26515\,
            I => \N__26478\
        );

    \I__5833\ : Span4Mux_h
    port map (
            O => \N__26510\,
            I => \N__26478\
        );

    \I__5832\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26475\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__26506\,
            I => \N__26468\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__26501\,
            I => \N__26468\
        );

    \I__5829\ : Span4Mux_v
    port map (
            O => \N__26498\,
            I => \N__26468\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__26495\,
            I => \N__26463\
        );

    \I__5827\ : Span12Mux_s10_v
    port map (
            O => \N__26492\,
            I => \N__26463\
        );

    \I__5826\ : Span4Mux_h
    port map (
            O => \N__26489\,
            I => \N__26460\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__26486\,
            I => \N__26457\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__26483\,
            I => \N__26454\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__26478\,
            I => \this_vga_signals.N_427_0\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__26475\,
            I => \this_vga_signals.N_427_0\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__26468\,
            I => \this_vga_signals.N_427_0\
        );

    \I__5820\ : Odrv12
    port map (
            O => \N__26463\,
            I => \this_vga_signals.N_427_0\
        );

    \I__5819\ : Odrv4
    port map (
            O => \N__26460\,
            I => \this_vga_signals.N_427_0\
        );

    \I__5818\ : Odrv12
    port map (
            O => \N__26457\,
            I => \this_vga_signals.N_427_0\
        );

    \I__5817\ : Odrv4
    port map (
            O => \N__26454\,
            I => \this_vga_signals.N_427_0\
        );

    \I__5816\ : CascadeMux
    port map (
            O => \N__26439\,
            I => \N__26426\
        );

    \I__5815\ : InMux
    port map (
            O => \N__26438\,
            I => \N__26405\
        );

    \I__5814\ : InMux
    port map (
            O => \N__26437\,
            I => \N__26405\
        );

    \I__5813\ : InMux
    port map (
            O => \N__26436\,
            I => \N__26405\
        );

    \I__5812\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26398\
        );

    \I__5811\ : InMux
    port map (
            O => \N__26434\,
            I => \N__26398\
        );

    \I__5810\ : InMux
    port map (
            O => \N__26433\,
            I => \N__26391\
        );

    \I__5809\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26391\
        );

    \I__5808\ : InMux
    port map (
            O => \N__26431\,
            I => \N__26391\
        );

    \I__5807\ : InMux
    port map (
            O => \N__26430\,
            I => \N__26388\
        );

    \I__5806\ : InMux
    port map (
            O => \N__26429\,
            I => \N__26385\
        );

    \I__5805\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26382\
        );

    \I__5804\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26377\
        );

    \I__5803\ : InMux
    port map (
            O => \N__26424\,
            I => \N__26377\
        );

    \I__5802\ : InMux
    port map (
            O => \N__26423\,
            I => \N__26370\
        );

    \I__5801\ : InMux
    port map (
            O => \N__26422\,
            I => \N__26370\
        );

    \I__5800\ : InMux
    port map (
            O => \N__26421\,
            I => \N__26370\
        );

    \I__5799\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26365\
        );

    \I__5798\ : InMux
    port map (
            O => \N__26419\,
            I => \N__26365\
        );

    \I__5797\ : InMux
    port map (
            O => \N__26418\,
            I => \N__26358\
        );

    \I__5796\ : InMux
    port map (
            O => \N__26417\,
            I => \N__26358\
        );

    \I__5795\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26358\
        );

    \I__5794\ : InMux
    port map (
            O => \N__26415\,
            I => \N__26353\
        );

    \I__5793\ : InMux
    port map (
            O => \N__26414\,
            I => \N__26353\
        );

    \I__5792\ : InMux
    port map (
            O => \N__26413\,
            I => \N__26348\
        );

    \I__5791\ : InMux
    port map (
            O => \N__26412\,
            I => \N__26348\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__26405\,
            I => \N__26345\
        );

    \I__5789\ : InMux
    port map (
            O => \N__26404\,
            I => \N__26340\
        );

    \I__5788\ : InMux
    port map (
            O => \N__26403\,
            I => \N__26340\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__26398\,
            I => \N__26335\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__26391\,
            I => \N__26335\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__26388\,
            I => \N__26332\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__26385\,
            I => \N__26317\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__26382\,
            I => \N__26317\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__26377\,
            I => \N__26317\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__26370\,
            I => \N__26317\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__26365\,
            I => \N__26317\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__26358\,
            I => \N__26317\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__26353\,
            I => \N__26317\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__26348\,
            I => \N__26302\
        );

    \I__5776\ : Span4Mux_v
    port map (
            O => \N__26345\,
            I => \N__26302\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__26340\,
            I => \N__26302\
        );

    \I__5774\ : Span4Mux_v
    port map (
            O => \N__26335\,
            I => \N__26302\
        );

    \I__5773\ : Span4Mux_h
    port map (
            O => \N__26332\,
            I => \N__26299\
        );

    \I__5772\ : Span4Mux_v
    port map (
            O => \N__26317\,
            I => \N__26296\
        );

    \I__5771\ : InMux
    port map (
            O => \N__26316\,
            I => \N__26291\
        );

    \I__5770\ : InMux
    port map (
            O => \N__26315\,
            I => \N__26291\
        );

    \I__5769\ : InMux
    port map (
            O => \N__26314\,
            I => \N__26282\
        );

    \I__5768\ : InMux
    port map (
            O => \N__26313\,
            I => \N__26282\
        );

    \I__5767\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26282\
        );

    \I__5766\ : InMux
    port map (
            O => \N__26311\,
            I => \N__26282\
        );

    \I__5765\ : Odrv4
    port map (
            O => \N__26302\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5764\ : Odrv4
    port map (
            O => \N__26299\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5763\ : Odrv4
    port map (
            O => \N__26296\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__26291\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__26282\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__5760\ : CascadeMux
    port map (
            O => \N__26271\,
            I => \this_vga_signals.N_427_0_cascade_\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__26268\,
            I => \N__26265\
        );

    \I__5758\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26262\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__26262\,
            I => \N__26259\
        );

    \I__5756\ : Span12Mux_s10_v
    port map (
            O => \N__26259\,
            I => \N__26256\
        );

    \I__5755\ : Odrv12
    port map (
            O => \N__26256\,
            I => \N_1274_tz_0\
        );

    \I__5754\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26250\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__26250\,
            I => \N__26247\
        );

    \I__5752\ : Span4Mux_h
    port map (
            O => \N__26247\,
            I => \N__26244\
        );

    \I__5751\ : Odrv4
    port map (
            O => \N__26244\,
            I => \M_this_sprites_address_qc_0_2\
        );

    \I__5750\ : InMux
    port map (
            O => \N__26241\,
            I => \N__26237\
        );

    \I__5749\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26234\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__26237\,
            I => \N__26229\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__26234\,
            I => \N__26229\
        );

    \I__5746\ : Span4Mux_h
    port map (
            O => \N__26229\,
            I => \N__26226\
        );

    \I__5745\ : Odrv4
    port map (
            O => \N__26226\,
            I => \this_vga_signals.N_889_0\
        );

    \I__5744\ : CascadeMux
    port map (
            O => \N__26223\,
            I => \this_vga_signals.N_889_0_cascade_\
        );

    \I__5743\ : CascadeMux
    port map (
            O => \N__26220\,
            I => \N__26211\
        );

    \I__5742\ : InMux
    port map (
            O => \N__26219\,
            I => \N__26208\
        );

    \I__5741\ : InMux
    port map (
            O => \N__26218\,
            I => \N__26199\
        );

    \I__5740\ : InMux
    port map (
            O => \N__26217\,
            I => \N__26199\
        );

    \I__5739\ : InMux
    port map (
            O => \N__26216\,
            I => \N__26196\
        );

    \I__5738\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26191\
        );

    \I__5737\ : InMux
    port map (
            O => \N__26214\,
            I => \N__26191\
        );

    \I__5736\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26188\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__26208\,
            I => \N__26185\
        );

    \I__5734\ : InMux
    port map (
            O => \N__26207\,
            I => \N__26179\
        );

    \I__5733\ : InMux
    port map (
            O => \N__26206\,
            I => \N__26179\
        );

    \I__5732\ : InMux
    port map (
            O => \N__26205\,
            I => \N__26174\
        );

    \I__5731\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26174\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__26199\,
            I => \N__26170\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__26196\,
            I => \N__26165\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__26191\,
            I => \N__26165\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__26188\,
            I => \N__26162\
        );

    \I__5726\ : Span4Mux_v
    port map (
            O => \N__26185\,
            I => \N__26159\
        );

    \I__5725\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26156\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__26179\,
            I => \N__26151\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__26174\,
            I => \N__26151\
        );

    \I__5722\ : InMux
    port map (
            O => \N__26173\,
            I => \N__26148\
        );

    \I__5721\ : Span4Mux_h
    port map (
            O => \N__26170\,
            I => \N__26143\
        );

    \I__5720\ : Span4Mux_h
    port map (
            O => \N__26165\,
            I => \N__26143\
        );

    \I__5719\ : Odrv4
    port map (
            O => \N__26162\,
            I => \N_750\
        );

    \I__5718\ : Odrv4
    port map (
            O => \N__26159\,
            I => \N_750\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__26156\,
            I => \N_750\
        );

    \I__5716\ : Odrv12
    port map (
            O => \N__26151\,
            I => \N_750\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__26148\,
            I => \N_750\
        );

    \I__5714\ : Odrv4
    port map (
            O => \N__26143\,
            I => \N_750\
        );

    \I__5713\ : CascadeMux
    port map (
            O => \N__26130\,
            I => \N__26126\
        );

    \I__5712\ : CascadeMux
    port map (
            O => \N__26129\,
            I => \N__26120\
        );

    \I__5711\ : InMux
    port map (
            O => \N__26126\,
            I => \N__26115\
        );

    \I__5710\ : InMux
    port map (
            O => \N__26125\,
            I => \N__26115\
        );

    \I__5709\ : InMux
    port map (
            O => \N__26124\,
            I => \N__26112\
        );

    \I__5708\ : InMux
    port map (
            O => \N__26123\,
            I => \N__26107\
        );

    \I__5707\ : InMux
    port map (
            O => \N__26120\,
            I => \N__26107\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__26115\,
            I => \N__26102\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__26112\,
            I => \N__26099\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__26107\,
            I => \N__26096\
        );

    \I__5703\ : InMux
    port map (
            O => \N__26106\,
            I => \N__26091\
        );

    \I__5702\ : InMux
    port map (
            O => \N__26105\,
            I => \N__26091\
        );

    \I__5701\ : Span4Mux_h
    port map (
            O => \N__26102\,
            I => \N__26086\
        );

    \I__5700\ : Span4Mux_h
    port map (
            O => \N__26099\,
            I => \N__26086\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__26096\,
            I => \N__26083\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__26091\,
            I => \N_762\
        );

    \I__5697\ : Odrv4
    port map (
            O => \N__26086\,
            I => \N_762\
        );

    \I__5696\ : Odrv4
    port map (
            O => \N__26083\,
            I => \N_762\
        );

    \I__5695\ : CascadeMux
    port map (
            O => \N__26076\,
            I => \N__26073\
        );

    \I__5694\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26069\
        );

    \I__5693\ : CascadeMux
    port map (
            O => \N__26072\,
            I => \N__26066\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__26069\,
            I => \N__26062\
        );

    \I__5691\ : InMux
    port map (
            O => \N__26066\,
            I => \N__26059\
        );

    \I__5690\ : CascadeMux
    port map (
            O => \N__26065\,
            I => \N__26056\
        );

    \I__5689\ : Span4Mux_v
    port map (
            O => \N__26062\,
            I => \N__26050\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__26059\,
            I => \N__26050\
        );

    \I__5687\ : InMux
    port map (
            O => \N__26056\,
            I => \N__26047\
        );

    \I__5686\ : CascadeMux
    port map (
            O => \N__26055\,
            I => \N__26044\
        );

    \I__5685\ : Span4Mux_h
    port map (
            O => \N__26050\,
            I => \N__26036\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__26047\,
            I => \N__26036\
        );

    \I__5683\ : InMux
    port map (
            O => \N__26044\,
            I => \N__26033\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__26043\,
            I => \N__26030\
        );

    \I__5681\ : CascadeMux
    port map (
            O => \N__26042\,
            I => \N__26025\
        );

    \I__5680\ : CascadeMux
    port map (
            O => \N__26041\,
            I => \N__26021\
        );

    \I__5679\ : Span4Mux_v
    port map (
            O => \N__26036\,
            I => \N__26012\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__26033\,
            I => \N__26012\
        );

    \I__5677\ : InMux
    port map (
            O => \N__26030\,
            I => \N__26009\
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__26029\,
            I => \N__26006\
        );

    \I__5675\ : CascadeMux
    port map (
            O => \N__26028\,
            I => \N__26003\
        );

    \I__5674\ : InMux
    port map (
            O => \N__26025\,
            I => \N__26000\
        );

    \I__5673\ : CascadeMux
    port map (
            O => \N__26024\,
            I => \N__25997\
        );

    \I__5672\ : InMux
    port map (
            O => \N__26021\,
            I => \N__25994\
        );

    \I__5671\ : CascadeMux
    port map (
            O => \N__26020\,
            I => \N__25991\
        );

    \I__5670\ : CascadeMux
    port map (
            O => \N__26019\,
            I => \N__25987\
        );

    \I__5669\ : CascadeMux
    port map (
            O => \N__26018\,
            I => \N__25984\
        );

    \I__5668\ : CascadeMux
    port map (
            O => \N__26017\,
            I => \N__25981\
        );

    \I__5667\ : Span4Mux_h
    port map (
            O => \N__26012\,
            I => \N__25975\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__26009\,
            I => \N__25975\
        );

    \I__5665\ : InMux
    port map (
            O => \N__26006\,
            I => \N__25972\
        );

    \I__5664\ : InMux
    port map (
            O => \N__26003\,
            I => \N__25969\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__26000\,
            I => \N__25966\
        );

    \I__5662\ : InMux
    port map (
            O => \N__25997\,
            I => \N__25963\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__25994\,
            I => \N__25960\
        );

    \I__5660\ : InMux
    port map (
            O => \N__25991\,
            I => \N__25957\
        );

    \I__5659\ : CascadeMux
    port map (
            O => \N__25990\,
            I => \N__25954\
        );

    \I__5658\ : InMux
    port map (
            O => \N__25987\,
            I => \N__25948\
        );

    \I__5657\ : InMux
    port map (
            O => \N__25984\,
            I => \N__25945\
        );

    \I__5656\ : InMux
    port map (
            O => \N__25981\,
            I => \N__25942\
        );

    \I__5655\ : CascadeMux
    port map (
            O => \N__25980\,
            I => \N__25939\
        );

    \I__5654\ : Span4Mux_v
    port map (
            O => \N__25975\,
            I => \N__25934\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__25972\,
            I => \N__25934\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__25969\,
            I => \N__25931\
        );

    \I__5651\ : Span4Mux_v
    port map (
            O => \N__25966\,
            I => \N__25926\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__25963\,
            I => \N__25926\
        );

    \I__5649\ : Span4Mux_v
    port map (
            O => \N__25960\,
            I => \N__25921\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__25957\,
            I => \N__25921\
        );

    \I__5647\ : InMux
    port map (
            O => \N__25954\,
            I => \N__25918\
        );

    \I__5646\ : CascadeMux
    port map (
            O => \N__25953\,
            I => \N__25915\
        );

    \I__5645\ : InMux
    port map (
            O => \N__25952\,
            I => \N__25912\
        );

    \I__5644\ : InMux
    port map (
            O => \N__25951\,
            I => \N__25909\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__25948\,
            I => \N__25904\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__25945\,
            I => \N__25904\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__25942\,
            I => \N__25901\
        );

    \I__5640\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25898\
        );

    \I__5639\ : Span4Mux_h
    port map (
            O => \N__25934\,
            I => \N__25895\
        );

    \I__5638\ : Span4Mux_v
    port map (
            O => \N__25931\,
            I => \N__25890\
        );

    \I__5637\ : Span4Mux_v
    port map (
            O => \N__25926\,
            I => \N__25890\
        );

    \I__5636\ : Span4Mux_v
    port map (
            O => \N__25921\,
            I => \N__25885\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__25918\,
            I => \N__25885\
        );

    \I__5634\ : InMux
    port map (
            O => \N__25915\,
            I => \N__25882\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__25912\,
            I => \N__25879\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__25909\,
            I => \N__25876\
        );

    \I__5631\ : Span12Mux_v
    port map (
            O => \N__25904\,
            I => \N__25868\
        );

    \I__5630\ : Span12Mux_s8_v
    port map (
            O => \N__25901\,
            I => \N__25868\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__25898\,
            I => \N__25868\
        );

    \I__5628\ : Span4Mux_v
    port map (
            O => \N__25895\,
            I => \N__25861\
        );

    \I__5627\ : Span4Mux_h
    port map (
            O => \N__25890\,
            I => \N__25861\
        );

    \I__5626\ : Span4Mux_h
    port map (
            O => \N__25885\,
            I => \N__25861\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__25882\,
            I => \N__25854\
        );

    \I__5624\ : Span4Mux_h
    port map (
            O => \N__25879\,
            I => \N__25854\
        );

    \I__5623\ : Span4Mux_v
    port map (
            O => \N__25876\,
            I => \N__25854\
        );

    \I__5622\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25851\
        );

    \I__5621\ : Odrv12
    port map (
            O => \N__25868\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__25861\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__25854\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__25851\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__5617\ : CascadeMux
    port map (
            O => \N__25842\,
            I => \N_750_cascade_\
        );

    \I__5616\ : InMux
    port map (
            O => \N__25839\,
            I => \N__25836\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__25836\,
            I => \M_this_sprites_address_qc_9_0\
        );

    \I__5614\ : CascadeMux
    port map (
            O => \N__25833\,
            I => \N__25830\
        );

    \I__5613\ : InMux
    port map (
            O => \N__25830\,
            I => \N__25825\
        );

    \I__5612\ : InMux
    port map (
            O => \N__25829\,
            I => \N__25822\
        );

    \I__5611\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25819\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__25825\,
            I => \N__25810\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__25822\,
            I => \N__25810\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__25819\,
            I => \N__25807\
        );

    \I__5607\ : InMux
    port map (
            O => \N__25818\,
            I => \N__25804\
        );

    \I__5606\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25798\
        );

    \I__5605\ : InMux
    port map (
            O => \N__25816\,
            I => \N__25798\
        );

    \I__5604\ : InMux
    port map (
            O => \N__25815\,
            I => \N__25795\
        );

    \I__5603\ : Span4Mux_v
    port map (
            O => \N__25810\,
            I => \N__25790\
        );

    \I__5602\ : Span4Mux_h
    port map (
            O => \N__25807\,
            I => \N__25790\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__25804\,
            I => \N__25787\
        );

    \I__5600\ : InMux
    port map (
            O => \N__25803\,
            I => \N__25784\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__25798\,
            I => \N__25779\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__25795\,
            I => \N__25779\
        );

    \I__5597\ : Span4Mux_v
    port map (
            O => \N__25790\,
            I => \N__25776\
        );

    \I__5596\ : Span4Mux_h
    port map (
            O => \N__25787\,
            I => \N__25771\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__25784\,
            I => \N__25771\
        );

    \I__5594\ : Span12Mux_h
    port map (
            O => \N__25779\,
            I => \N__25768\
        );

    \I__5593\ : Span4Mux_v
    port map (
            O => \N__25776\,
            I => \N__25765\
        );

    \I__5592\ : Sp12to4
    port map (
            O => \N__25771\,
            I => \N__25762\
        );

    \I__5591\ : Odrv12
    port map (
            O => \N__25768\,
            I => port_address_in_0
        );

    \I__5590\ : Odrv4
    port map (
            O => \N__25765\,
            I => port_address_in_0
        );

    \I__5589\ : Odrv12
    port map (
            O => \N__25762\,
            I => port_address_in_0
        );

    \I__5588\ : InMux
    port map (
            O => \N__25755\,
            I => \N__25752\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__25752\,
            I => \N__25749\
        );

    \I__5586\ : Odrv4
    port map (
            O => \N__25749\,
            I => \this_vga_signals.N_648\
        );

    \I__5585\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25739\
        );

    \I__5584\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25736\
        );

    \I__5583\ : InMux
    port map (
            O => \N__25744\,
            I => \N__25733\
        );

    \I__5582\ : InMux
    port map (
            O => \N__25743\,
            I => \N__25730\
        );

    \I__5581\ : CascadeMux
    port map (
            O => \N__25742\,
            I => \N__25727\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__25739\,
            I => \N__25723\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__25736\,
            I => \N__25718\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__25733\,
            I => \N__25718\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__25730\,
            I => \N__25715\
        );

    \I__5576\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25712\
        );

    \I__5575\ : CascadeMux
    port map (
            O => \N__25726\,
            I => \N__25708\
        );

    \I__5574\ : Span4Mux_v
    port map (
            O => \N__25723\,
            I => \N__25704\
        );

    \I__5573\ : Span4Mux_v
    port map (
            O => \N__25718\,
            I => \N__25697\
        );

    \I__5572\ : Span4Mux_v
    port map (
            O => \N__25715\,
            I => \N__25697\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__25712\,
            I => \N__25697\
        );

    \I__5570\ : InMux
    port map (
            O => \N__25711\,
            I => \N__25694\
        );

    \I__5569\ : InMux
    port map (
            O => \N__25708\,
            I => \N__25689\
        );

    \I__5568\ : InMux
    port map (
            O => \N__25707\,
            I => \N__25689\
        );

    \I__5567\ : Span4Mux_h
    port map (
            O => \N__25704\,
            I => \N__25684\
        );

    \I__5566\ : Span4Mux_h
    port map (
            O => \N__25697\,
            I => \N__25684\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__25694\,
            I => \N__25679\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__25689\,
            I => \N__25679\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__25684\,
            I => \N__25676\
        );

    \I__5562\ : Span12Mux_h
    port map (
            O => \N__25679\,
            I => \N__25673\
        );

    \I__5561\ : Sp12to4
    port map (
            O => \N__25676\,
            I => \N__25670\
        );

    \I__5560\ : Odrv12
    port map (
            O => \N__25673\,
            I => port_address_in_1
        );

    \I__5559\ : Odrv12
    port map (
            O => \N__25670\,
            I => port_address_in_1
        );

    \I__5558\ : InMux
    port map (
            O => \N__25665\,
            I => \N__25659\
        );

    \I__5557\ : InMux
    port map (
            O => \N__25664\,
            I => \N__25655\
        );

    \I__5556\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25650\
        );

    \I__5555\ : InMux
    port map (
            O => \N__25662\,
            I => \N__25650\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__25659\,
            I => \N__25646\
        );

    \I__5553\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25643\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__25655\,
            I => \N__25640\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__25650\,
            I => \N__25637\
        );

    \I__5550\ : InMux
    port map (
            O => \N__25649\,
            I => \N__25634\
        );

    \I__5549\ : Span4Mux_h
    port map (
            O => \N__25646\,
            I => \N__25629\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__25643\,
            I => \N__25629\
        );

    \I__5547\ : Span4Mux_v
    port map (
            O => \N__25640\,
            I => \N__25622\
        );

    \I__5546\ : Span4Mux_h
    port map (
            O => \N__25637\,
            I => \N__25622\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__25634\,
            I => \N__25622\
        );

    \I__5544\ : Span4Mux_h
    port map (
            O => \N__25629\,
            I => \N__25619\
        );

    \I__5543\ : Span4Mux_h
    port map (
            O => \N__25622\,
            I => \N__25616\
        );

    \I__5542\ : Sp12to4
    port map (
            O => \N__25619\,
            I => \N__25613\
        );

    \I__5541\ : Span4Mux_v
    port map (
            O => \N__25616\,
            I => \N__25610\
        );

    \I__5540\ : Span12Mux_v
    port map (
            O => \N__25613\,
            I => \N__25607\
        );

    \I__5539\ : Span4Mux_v
    port map (
            O => \N__25610\,
            I => \N__25604\
        );

    \I__5538\ : Odrv12
    port map (
            O => \N__25607\,
            I => port_address_in_2
        );

    \I__5537\ : Odrv4
    port map (
            O => \N__25604\,
            I => port_address_in_2
        );

    \I__5536\ : InMux
    port map (
            O => \N__25599\,
            I => \N__25596\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__25596\,
            I => \N__25592\
        );

    \I__5534\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25589\
        );

    \I__5533\ : Span4Mux_v
    port map (
            O => \N__25592\,
            I => \N__25584\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__25589\,
            I => \N__25584\
        );

    \I__5531\ : Span4Mux_h
    port map (
            O => \N__25584\,
            I => \N__25581\
        );

    \I__5530\ : Sp12to4
    port map (
            O => \N__25581\,
            I => \N__25578\
        );

    \I__5529\ : Span12Mux_v
    port map (
            O => \N__25578\,
            I => \N__25575\
        );

    \I__5528\ : Span12Mux_v
    port map (
            O => \N__25575\,
            I => \N__25572\
        );

    \I__5527\ : Odrv12
    port map (
            O => \N__25572\,
            I => port_address_in_7
        );

    \I__5526\ : InMux
    port map (
            O => \N__25569\,
            I => \N__25565\
        );

    \I__5525\ : InMux
    port map (
            O => \N__25568\,
            I => \N__25562\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__25565\,
            I => \N__25559\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__25562\,
            I => \N__25556\
        );

    \I__5522\ : Span4Mux_h
    port map (
            O => \N__25559\,
            I => \N__25551\
        );

    \I__5521\ : Span4Mux_v
    port map (
            O => \N__25556\,
            I => \N__25551\
        );

    \I__5520\ : Sp12to4
    port map (
            O => \N__25551\,
            I => \N__25548\
        );

    \I__5519\ : Span12Mux_h
    port map (
            O => \N__25548\,
            I => \N__25544\
        );

    \I__5518\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25541\
        );

    \I__5517\ : Odrv12
    port map (
            O => \N__25544\,
            I => port_rw_in
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__25541\,
            I => port_rw_in
        );

    \I__5515\ : CascadeMux
    port map (
            O => \N__25536\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_5LZ0Z8_cascade_\
        );

    \I__5514\ : InMux
    port map (
            O => \N__25533\,
            I => \N__25530\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__25530\,
            I => \N__25527\
        );

    \I__5512\ : Span4Mux_h
    port map (
            O => \N__25527\,
            I => \N__25524\
        );

    \I__5511\ : Odrv4
    port map (
            O => \N__25524\,
            I => \M_this_substate_d_0_sqmuxa\
        );

    \I__5510\ : CascadeMux
    port map (
            O => \N__25521\,
            I => \M_this_substate_d_0_sqmuxa_cascade_\
        );

    \I__5509\ : InMux
    port map (
            O => \N__25518\,
            I => \N__25515\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__25515\,
            I => \N__25512\
        );

    \I__5507\ : Span4Mux_v
    port map (
            O => \N__25512\,
            I => \N__25509\
        );

    \I__5506\ : Odrv4
    port map (
            O => \N__25509\,
            I => dma_c4_1_0
        );

    \I__5505\ : InMux
    port map (
            O => \N__25506\,
            I => \N__25495\
        );

    \I__5504\ : InMux
    port map (
            O => \N__25505\,
            I => \N__25492\
        );

    \I__5503\ : InMux
    port map (
            O => \N__25504\,
            I => \N__25487\
        );

    \I__5502\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25487\
        );

    \I__5501\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25479\
        );

    \I__5500\ : InMux
    port map (
            O => \N__25501\,
            I => \N__25476\
        );

    \I__5499\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25473\
        );

    \I__5498\ : CascadeMux
    port map (
            O => \N__25499\,
            I => \N__25469\
        );

    \I__5497\ : InMux
    port map (
            O => \N__25498\,
            I => \N__25465\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__25495\,
            I => \N__25462\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__25492\,
            I => \N__25459\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__25487\,
            I => \N__25456\
        );

    \I__5493\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25451\
        );

    \I__5492\ : InMux
    port map (
            O => \N__25485\,
            I => \N__25451\
        );

    \I__5491\ : InMux
    port map (
            O => \N__25484\,
            I => \N__25448\
        );

    \I__5490\ : InMux
    port map (
            O => \N__25483\,
            I => \N__25443\
        );

    \I__5489\ : InMux
    port map (
            O => \N__25482\,
            I => \N__25443\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__25479\,
            I => \N__25436\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__25476\,
            I => \N__25436\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__25473\,
            I => \N__25436\
        );

    \I__5485\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25433\
        );

    \I__5484\ : InMux
    port map (
            O => \N__25469\,
            I => \N__25430\
        );

    \I__5483\ : InMux
    port map (
            O => \N__25468\,
            I => \N__25427\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__25465\,
            I => \N__25424\
        );

    \I__5481\ : Span4Mux_v
    port map (
            O => \N__25462\,
            I => \N__25419\
        );

    \I__5480\ : Span4Mux_v
    port map (
            O => \N__25459\,
            I => \N__25419\
        );

    \I__5479\ : Span4Mux_h
    port map (
            O => \N__25456\,
            I => \N__25408\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__25451\,
            I => \N__25408\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__25448\,
            I => \N__25408\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__25443\,
            I => \N__25408\
        );

    \I__5475\ : Span4Mux_v
    port map (
            O => \N__25436\,
            I => \N__25408\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__25433\,
            I => \N__25403\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__25430\,
            I => \N__25403\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__25427\,
            I => \this_vga_signals.N_732\
        );

    \I__5471\ : Odrv4
    port map (
            O => \N__25424\,
            I => \this_vga_signals.N_732\
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__25419\,
            I => \this_vga_signals.N_732\
        );

    \I__5469\ : Odrv4
    port map (
            O => \N__25408\,
            I => \this_vga_signals.N_732\
        );

    \I__5468\ : Odrv12
    port map (
            O => \N__25403\,
            I => \this_vga_signals.N_732\
        );

    \I__5467\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25386\
        );

    \I__5466\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25386\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__25386\,
            I => \un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0\
        );

    \I__5464\ : CascadeMux
    port map (
            O => \N__25383\,
            I => \N_622_cascade_\
        );

    \I__5463\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25377\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__25377\,
            I => \N_1278_tz_0\
        );

    \I__5461\ : CascadeMux
    port map (
            O => \N__25374\,
            I => \N__25371\
        );

    \I__5460\ : InMux
    port map (
            O => \N__25371\,
            I => \N__25368\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__25368\,
            I => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_12\
        );

    \I__5458\ : CascadeMux
    port map (
            O => \N__25365\,
            I => \N_460_0_cascade_\
        );

    \I__5457\ : CascadeMux
    port map (
            O => \N__25362\,
            I => \N__25359\
        );

    \I__5456\ : InMux
    port map (
            O => \N__25359\,
            I => \N__25354\
        );

    \I__5455\ : InMux
    port map (
            O => \N__25358\,
            I => \N__25341\
        );

    \I__5454\ : InMux
    port map (
            O => \N__25357\,
            I => \N__25341\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__25354\,
            I => \N__25338\
        );

    \I__5452\ : InMux
    port map (
            O => \N__25353\,
            I => \N__25329\
        );

    \I__5451\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25329\
        );

    \I__5450\ : InMux
    port map (
            O => \N__25351\,
            I => \N__25329\
        );

    \I__5449\ : InMux
    port map (
            O => \N__25350\,
            I => \N__25329\
        );

    \I__5448\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25320\
        );

    \I__5447\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25320\
        );

    \I__5446\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25320\
        );

    \I__5445\ : InMux
    port map (
            O => \N__25346\,
            I => \N__25320\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__25341\,
            I => \N__25317\
        );

    \I__5443\ : Span4Mux_v
    port map (
            O => \N__25338\,
            I => \N__25314\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__25329\,
            I => \N__25307\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__25320\,
            I => \N__25307\
        );

    \I__5440\ : Span12Mux_s5_v
    port map (
            O => \N__25317\,
            I => \N__25307\
        );

    \I__5439\ : Span4Mux_v
    port map (
            O => \N__25314\,
            I => \N__25304\
        );

    \I__5438\ : Odrv12
    port map (
            O => \N__25307\,
            I => \N_560\
        );

    \I__5437\ : Odrv4
    port map (
            O => \N__25304\,
            I => \N_560\
        );

    \I__5436\ : CEMux
    port map (
            O => \N__25299\,
            I => \N__25296\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__25296\,
            I => \N__25287\
        );

    \I__5434\ : InMux
    port map (
            O => \N__25295\,
            I => \N__25284\
        );

    \I__5433\ : InMux
    port map (
            O => \N__25294\,
            I => \N__25281\
        );

    \I__5432\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25278\
        );

    \I__5431\ : CEMux
    port map (
            O => \N__25292\,
            I => \N__25273\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__25291\,
            I => \N__25270\
        );

    \I__5429\ : InMux
    port map (
            O => \N__25290\,
            I => \N__25267\
        );

    \I__5428\ : Span4Mux_h
    port map (
            O => \N__25287\,
            I => \N__25259\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__25284\,
            I => \N__25259\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__25281\,
            I => \N__25259\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__25278\,
            I => \N__25256\
        );

    \I__5424\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25251\
        );

    \I__5423\ : InMux
    port map (
            O => \N__25276\,
            I => \N__25251\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__25273\,
            I => \N__25248\
        );

    \I__5421\ : InMux
    port map (
            O => \N__25270\,
            I => \N__25245\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__25267\,
            I => \N__25242\
        );

    \I__5419\ : InMux
    port map (
            O => \N__25266\,
            I => \N__25239\
        );

    \I__5418\ : Span4Mux_v
    port map (
            O => \N__25259\,
            I => \N__25236\
        );

    \I__5417\ : Span4Mux_v
    port map (
            O => \N__25256\,
            I => \N__25231\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__25251\,
            I => \N__25231\
        );

    \I__5415\ : Span4Mux_v
    port map (
            O => \N__25248\,
            I => \N__25224\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__25245\,
            I => \N__25224\
        );

    \I__5413\ : Span4Mux_h
    port map (
            O => \N__25242\,
            I => \N__25219\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__25239\,
            I => \N__25219\
        );

    \I__5411\ : Span4Mux_h
    port map (
            O => \N__25236\,
            I => \N__25214\
        );

    \I__5410\ : Span4Mux_v
    port map (
            O => \N__25231\,
            I => \N__25214\
        );

    \I__5409\ : InMux
    port map (
            O => \N__25230\,
            I => \N__25209\
        );

    \I__5408\ : InMux
    port map (
            O => \N__25229\,
            I => \N__25209\
        );

    \I__5407\ : Span4Mux_h
    port map (
            O => \N__25224\,
            I => \N__25206\
        );

    \I__5406\ : Span4Mux_h
    port map (
            O => \N__25219\,
            I => \N__25202\
        );

    \I__5405\ : Span4Mux_v
    port map (
            O => \N__25214\,
            I => \N__25199\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__25209\,
            I => \N__25194\
        );

    \I__5403\ : Sp12to4
    port map (
            O => \N__25206\,
            I => \N__25194\
        );

    \I__5402\ : InMux
    port map (
            O => \N__25205\,
            I => \N__25191\
        );

    \I__5401\ : Span4Mux_v
    port map (
            O => \N__25202\,
            I => \N__25188\
        );

    \I__5400\ : Sp12to4
    port map (
            O => \N__25199\,
            I => \N__25183\
        );

    \I__5399\ : Span12Mux_v
    port map (
            O => \N__25194\,
            I => \N__25183\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__25191\,
            I => \M_this_map_ram_write_en_0\
        );

    \I__5397\ : Odrv4
    port map (
            O => \N__25188\,
            I => \M_this_map_ram_write_en_0\
        );

    \I__5396\ : Odrv12
    port map (
            O => \N__25183\,
            I => \M_this_map_ram_write_en_0\
        );

    \I__5395\ : CascadeMux
    port map (
            O => \N__25176\,
            I => \N_888_0_cascade_\
        );

    \I__5394\ : CascadeMux
    port map (
            O => \N__25173\,
            I => \N__25170\
        );

    \I__5393\ : InMux
    port map (
            O => \N__25170\,
            I => \N__25167\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__25167\,
            I => \this_vga_signals.N_779\
        );

    \I__5391\ : InMux
    port map (
            O => \N__25164\,
            I => \N__25159\
        );

    \I__5390\ : InMux
    port map (
            O => \N__25163\,
            I => \N__25156\
        );

    \I__5389\ : InMux
    port map (
            O => \N__25162\,
            I => \N__25150\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__25159\,
            I => \N__25145\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__25156\,
            I => \N__25145\
        );

    \I__5386\ : InMux
    port map (
            O => \N__25155\,
            I => \N__25142\
        );

    \I__5385\ : InMux
    port map (
            O => \N__25154\,
            I => \N__25137\
        );

    \I__5384\ : InMux
    port map (
            O => \N__25153\,
            I => \N__25137\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__25150\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__5382\ : Odrv4
    port map (
            O => \N__25145\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__25142\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__25137\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__5379\ : CascadeMux
    port map (
            O => \N__25128\,
            I => \N__25123\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__25127\,
            I => \N__25120\
        );

    \I__5377\ : InMux
    port map (
            O => \N__25126\,
            I => \N__25112\
        );

    \I__5376\ : InMux
    port map (
            O => \N__25123\,
            I => \N__25112\
        );

    \I__5375\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25109\
        );

    \I__5374\ : InMux
    port map (
            O => \N__25119\,
            I => \N__25103\
        );

    \I__5373\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25103\
        );

    \I__5372\ : CascadeMux
    port map (
            O => \N__25117\,
            I => \N__25100\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__25112\,
            I => \N__25095\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__25109\,
            I => \N__25095\
        );

    \I__5369\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25092\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__25103\,
            I => \N__25089\
        );

    \I__5367\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25086\
        );

    \I__5366\ : Span4Mux_v
    port map (
            O => \N__25095\,
            I => \N__25083\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__25092\,
            I => \N__25080\
        );

    \I__5364\ : Span4Mux_h
    port map (
            O => \N__25089\,
            I => \N__25075\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__25086\,
            I => \N__25075\
        );

    \I__5362\ : Span4Mux_h
    port map (
            O => \N__25083\,
            I => \N__25072\
        );

    \I__5361\ : Span4Mux_v
    port map (
            O => \N__25080\,
            I => \N__25067\
        );

    \I__5360\ : Span4Mux_v
    port map (
            O => \N__25075\,
            I => \N__25067\
        );

    \I__5359\ : Sp12to4
    port map (
            O => \N__25072\,
            I => \N__25062\
        );

    \I__5358\ : Sp12to4
    port map (
            O => \N__25067\,
            I => \N__25062\
        );

    \I__5357\ : Span12Mux_h
    port map (
            O => \N__25062\,
            I => \N__25059\
        );

    \I__5356\ : Odrv12
    port map (
            O => \N__25059\,
            I => port_enb_c
        );

    \I__5355\ : InMux
    port map (
            O => \N__25056\,
            I => \N__25051\
        );

    \I__5354\ : InMux
    port map (
            O => \N__25055\,
            I => \N__25048\
        );

    \I__5353\ : InMux
    port map (
            O => \N__25054\,
            I => \N__25041\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__25051\,
            I => \N__25036\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__25048\,
            I => \N__25036\
        );

    \I__5350\ : InMux
    port map (
            O => \N__25047\,
            I => \N__25031\
        );

    \I__5349\ : InMux
    port map (
            O => \N__25046\,
            I => \N__25031\
        );

    \I__5348\ : InMux
    port map (
            O => \N__25045\,
            I => \N__25026\
        );

    \I__5347\ : InMux
    port map (
            O => \N__25044\,
            I => \N__25026\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__25041\,
            I => \M_this_delay_clk_out_0\
        );

    \I__5345\ : Odrv4
    port map (
            O => \N__25036\,
            I => \M_this_delay_clk_out_0\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__25031\,
            I => \M_this_delay_clk_out_0\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__25026\,
            I => \M_this_delay_clk_out_0\
        );

    \I__5342\ : IoInMux
    port map (
            O => \N__25017\,
            I => \N__25014\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__25014\,
            I => \N__25011\
        );

    \I__5340\ : IoSpan4Mux
    port map (
            O => \N__25011\,
            I => \N__25008\
        );

    \I__5339\ : Span4Mux_s2_v
    port map (
            O => \N__25008\,
            I => \N__25005\
        );

    \I__5338\ : Span4Mux_v
    port map (
            O => \N__25005\,
            I => \N__25002\
        );

    \I__5337\ : Span4Mux_v
    port map (
            O => \N__25002\,
            I => \N__24999\
        );

    \I__5336\ : Odrv4
    port map (
            O => \N__24999\,
            I => \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\
        );

    \I__5335\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24993\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__24993\,
            I => \N__24990\
        );

    \I__5333\ : Odrv4
    port map (
            O => \N__24990\,
            I => \M_this_state_q_RNI0A0EZ0Z_6\
        );

    \I__5332\ : CascadeMux
    port map (
            O => \N__24987\,
            I => \M_this_state_q_RNI244K2Z0Z_6_cascade_\
        );

    \I__5331\ : IoInMux
    port map (
            O => \N__24984\,
            I => \N__24981\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__24981\,
            I => \N__24976\
        );

    \I__5329\ : InMux
    port map (
            O => \N__24980\,
            I => \N__24973\
        );

    \I__5328\ : InMux
    port map (
            O => \N__24979\,
            I => \N__24970\
        );

    \I__5327\ : IoSpan4Mux
    port map (
            O => \N__24976\,
            I => \N__24967\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__24973\,
            I => \N__24964\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__24970\,
            I => \N__24961\
        );

    \I__5324\ : Span4Mux_s2_h
    port map (
            O => \N__24967\,
            I => \N__24958\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__24964\,
            I => \N__24955\
        );

    \I__5322\ : Span4Mux_v
    port map (
            O => \N__24961\,
            I => \N__24952\
        );

    \I__5321\ : Sp12to4
    port map (
            O => \N__24958\,
            I => \N__24948\
        );

    \I__5320\ : Span4Mux_v
    port map (
            O => \N__24955\,
            I => \N__24943\
        );

    \I__5319\ : Span4Mux_v
    port map (
            O => \N__24952\,
            I => \N__24943\
        );

    \I__5318\ : InMux
    port map (
            O => \N__24951\,
            I => \N__24940\
        );

    \I__5317\ : Span12Mux_h
    port map (
            O => \N__24948\,
            I => \N__24936\
        );

    \I__5316\ : Sp12to4
    port map (
            O => \N__24943\,
            I => \N__24933\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__24940\,
            I => \N__24930\
        );

    \I__5314\ : CascadeMux
    port map (
            O => \N__24939\,
            I => \N__24927\
        );

    \I__5313\ : Span12Mux_v
    port map (
            O => \N__24936\,
            I => \N__24922\
        );

    \I__5312\ : Span12Mux_h
    port map (
            O => \N__24933\,
            I => \N__24922\
        );

    \I__5311\ : Span4Mux_v
    port map (
            O => \N__24930\,
            I => \N__24919\
        );

    \I__5310\ : InMux
    port map (
            O => \N__24927\,
            I => \N__24916\
        );

    \I__5309\ : Odrv12
    port map (
            O => \N__24922\,
            I => dma_0
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__24919\,
            I => dma_0
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__24916\,
            I => dma_0
        );

    \I__5306\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24906\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__24906\,
            I => \N__24903\
        );

    \I__5304\ : Odrv4
    port map (
            O => \N__24903\,
            I => \M_this_state_q_fastZ0Z_9\
        );

    \I__5303\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24897\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__24897\,
            I => \N__24894\
        );

    \I__5301\ : Span4Mux_v
    port map (
            O => \N__24894\,
            I => \N__24891\
        );

    \I__5300\ : Odrv4
    port map (
            O => \N__24891\,
            I => \N_861\
        );

    \I__5299\ : CascadeMux
    port map (
            O => \N__24888\,
            I => \N_861_cascade_\
        );

    \I__5298\ : InMux
    port map (
            O => \N__24885\,
            I => \N__24882\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__24882\,
            I => dma_c4_1
        );

    \I__5296\ : CascadeMux
    port map (
            O => \N__24879\,
            I => \N__24876\
        );

    \I__5295\ : InMux
    port map (
            O => \N__24876\,
            I => \N__24873\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__24873\,
            I => this_vga_signals_un20_i_a2_4_a3_0_a4_2_1
        );

    \I__5293\ : InMux
    port map (
            O => \N__24870\,
            I => \N__24867\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__24867\,
            I => \this_ppu.un1_M_haddress_q_2_cry_7_THRU_CO\
        );

    \I__5291\ : CascadeMux
    port map (
            O => \N__24864\,
            I => \N__24861\
        );

    \I__5290\ : InMux
    port map (
            O => \N__24861\,
            I => \N__24858\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__24858\,
            I => \this_ppu.un1_M_haddress_q_cry_7_THRU_CO\
        );

    \I__5288\ : InMux
    port map (
            O => \N__24855\,
            I => \bfn_20_7_0_\
        );

    \I__5287\ : InMux
    port map (
            O => \N__24852\,
            I => \N__24849\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__24849\,
            I => \N__24845\
        );

    \I__5285\ : InMux
    port map (
            O => \N__24848\,
            I => \N__24842\
        );

    \I__5284\ : Span4Mux_v
    port map (
            O => \N__24845\,
            I => \N__24839\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__24842\,
            I => \N__24836\
        );

    \I__5282\ : Span4Mux_v
    port map (
            O => \N__24839\,
            I => \N__24833\
        );

    \I__5281\ : Span4Mux_v
    port map (
            O => \N__24836\,
            I => \N__24830\
        );

    \I__5280\ : Odrv4
    port map (
            O => \N__24833\,
            I => \this_ppu.vscroll8\
        );

    \I__5279\ : Odrv4
    port map (
            O => \N__24830\,
            I => \this_ppu.vscroll8\
        );

    \I__5278\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24822\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__24822\,
            I => \M_this_oam_ram_read_data_i_11\
        );

    \I__5276\ : InMux
    port map (
            O => \N__24819\,
            I => \N__24816\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__24816\,
            I => \this_ppu.un2_vscroll_axb_0\
        );

    \I__5274\ : CascadeMux
    port map (
            O => \N__24813\,
            I => \N__24805\
        );

    \I__5273\ : CascadeMux
    port map (
            O => \N__24812\,
            I => \N__24799\
        );

    \I__5272\ : CascadeMux
    port map (
            O => \N__24811\,
            I => \N__24796\
        );

    \I__5271\ : CascadeMux
    port map (
            O => \N__24810\,
            I => \N__24793\
        );

    \I__5270\ : CascadeMux
    port map (
            O => \N__24809\,
            I => \N__24790\
        );

    \I__5269\ : CascadeMux
    port map (
            O => \N__24808\,
            I => \N__24787\
        );

    \I__5268\ : InMux
    port map (
            O => \N__24805\,
            I => \N__24784\
        );

    \I__5267\ : CascadeMux
    port map (
            O => \N__24804\,
            I => \N__24781\
        );

    \I__5266\ : CascadeMux
    port map (
            O => \N__24803\,
            I => \N__24777\
        );

    \I__5265\ : CascadeMux
    port map (
            O => \N__24802\,
            I => \N__24769\
        );

    \I__5264\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24765\
        );

    \I__5263\ : InMux
    port map (
            O => \N__24796\,
            I => \N__24762\
        );

    \I__5262\ : InMux
    port map (
            O => \N__24793\,
            I => \N__24759\
        );

    \I__5261\ : InMux
    port map (
            O => \N__24790\,
            I => \N__24756\
        );

    \I__5260\ : InMux
    port map (
            O => \N__24787\,
            I => \N__24753\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__24784\,
            I => \N__24750\
        );

    \I__5258\ : InMux
    port map (
            O => \N__24781\,
            I => \N__24747\
        );

    \I__5257\ : CascadeMux
    port map (
            O => \N__24780\,
            I => \N__24744\
        );

    \I__5256\ : InMux
    port map (
            O => \N__24777\,
            I => \N__24741\
        );

    \I__5255\ : CascadeMux
    port map (
            O => \N__24776\,
            I => \N__24738\
        );

    \I__5254\ : CascadeMux
    port map (
            O => \N__24775\,
            I => \N__24735\
        );

    \I__5253\ : CascadeMux
    port map (
            O => \N__24774\,
            I => \N__24732\
        );

    \I__5252\ : CascadeMux
    port map (
            O => \N__24773\,
            I => \N__24729\
        );

    \I__5251\ : CascadeMux
    port map (
            O => \N__24772\,
            I => \N__24726\
        );

    \I__5250\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24723\
        );

    \I__5249\ : CascadeMux
    port map (
            O => \N__24768\,
            I => \N__24720\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__24765\,
            I => \N__24711\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__24762\,
            I => \N__24711\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__24759\,
            I => \N__24711\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__24756\,
            I => \N__24711\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__24753\,
            I => \N__24708\
        );

    \I__5243\ : Span4Mux_v
    port map (
            O => \N__24750\,
            I => \N__24703\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__24747\,
            I => \N__24703\
        );

    \I__5241\ : InMux
    port map (
            O => \N__24744\,
            I => \N__24700\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__24741\,
            I => \N__24697\
        );

    \I__5239\ : InMux
    port map (
            O => \N__24738\,
            I => \N__24694\
        );

    \I__5238\ : InMux
    port map (
            O => \N__24735\,
            I => \N__24691\
        );

    \I__5237\ : InMux
    port map (
            O => \N__24732\,
            I => \N__24688\
        );

    \I__5236\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24685\
        );

    \I__5235\ : InMux
    port map (
            O => \N__24726\,
            I => \N__24682\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__24723\,
            I => \N__24679\
        );

    \I__5233\ : InMux
    port map (
            O => \N__24720\,
            I => \N__24676\
        );

    \I__5232\ : Span12Mux_v
    port map (
            O => \N__24711\,
            I => \N__24673\
        );

    \I__5231\ : Span12Mux_s5_v
    port map (
            O => \N__24708\,
            I => \N__24658\
        );

    \I__5230\ : Sp12to4
    port map (
            O => \N__24703\,
            I => \N__24658\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__24700\,
            I => \N__24658\
        );

    \I__5228\ : Sp12to4
    port map (
            O => \N__24697\,
            I => \N__24658\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__24694\,
            I => \N__24658\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__24691\,
            I => \N__24658\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__24688\,
            I => \N__24658\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__24685\,
            I => \N__24653\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__24682\,
            I => \N__24653\
        );

    \I__5222\ : Span4Mux_h
    port map (
            O => \N__24679\,
            I => \N__24650\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__24676\,
            I => \N__24647\
        );

    \I__5220\ : Span12Mux_h
    port map (
            O => \N__24673\,
            I => \N__24644\
        );

    \I__5219\ : Span12Mux_v
    port map (
            O => \N__24658\,
            I => \N__24639\
        );

    \I__5218\ : Span12Mux_v
    port map (
            O => \N__24653\,
            I => \N__24639\
        );

    \I__5217\ : Span4Mux_v
    port map (
            O => \N__24650\,
            I => \N__24634\
        );

    \I__5216\ : Span4Mux_h
    port map (
            O => \N__24647\,
            I => \N__24634\
        );

    \I__5215\ : Odrv12
    port map (
            O => \N__24644\,
            I => \M_this_ppu_sprites_addr_3\
        );

    \I__5214\ : Odrv12
    port map (
            O => \N__24639\,
            I => \M_this_ppu_sprites_addr_3\
        );

    \I__5213\ : Odrv4
    port map (
            O => \N__24634\,
            I => \M_this_ppu_sprites_addr_3\
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__24627\,
            I => \N__24624\
        );

    \I__5211\ : InMux
    port map (
            O => \N__24624\,
            I => \N__24620\
        );

    \I__5210\ : CascadeMux
    port map (
            O => \N__24623\,
            I => \N__24617\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__24620\,
            I => \N__24612\
        );

    \I__5208\ : InMux
    port map (
            O => \N__24617\,
            I => \N__24609\
        );

    \I__5207\ : CascadeMux
    port map (
            O => \N__24616\,
            I => \N__24606\
        );

    \I__5206\ : CascadeMux
    port map (
            O => \N__24615\,
            I => \N__24602\
        );

    \I__5205\ : Span4Mux_v
    port map (
            O => \N__24612\,
            I => \N__24597\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__24609\,
            I => \N__24597\
        );

    \I__5203\ : InMux
    port map (
            O => \N__24606\,
            I => \N__24594\
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__24605\,
            I => \N__24590\
        );

    \I__5201\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24577\
        );

    \I__5200\ : Span4Mux_h
    port map (
            O => \N__24597\,
            I => \N__24572\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__24594\,
            I => \N__24572\
        );

    \I__5198\ : CascadeMux
    port map (
            O => \N__24593\,
            I => \N__24569\
        );

    \I__5197\ : InMux
    port map (
            O => \N__24590\,
            I => \N__24566\
        );

    \I__5196\ : CascadeMux
    port map (
            O => \N__24589\,
            I => \N__24563\
        );

    \I__5195\ : CascadeMux
    port map (
            O => \N__24588\,
            I => \N__24560\
        );

    \I__5194\ : CascadeMux
    port map (
            O => \N__24587\,
            I => \N__24557\
        );

    \I__5193\ : CascadeMux
    port map (
            O => \N__24586\,
            I => \N__24554\
        );

    \I__5192\ : CascadeMux
    port map (
            O => \N__24585\,
            I => \N__24551\
        );

    \I__5191\ : CascadeMux
    port map (
            O => \N__24584\,
            I => \N__24548\
        );

    \I__5190\ : CascadeMux
    port map (
            O => \N__24583\,
            I => \N__24545\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__24582\,
            I => \N__24542\
        );

    \I__5188\ : CascadeMux
    port map (
            O => \N__24581\,
            I => \N__24539\
        );

    \I__5187\ : CascadeMux
    port map (
            O => \N__24580\,
            I => \N__24536\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__24577\,
            I => \N__24533\
        );

    \I__5185\ : Span4Mux_v
    port map (
            O => \N__24572\,
            I => \N__24530\
        );

    \I__5184\ : InMux
    port map (
            O => \N__24569\,
            I => \N__24527\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__24566\,
            I => \N__24524\
        );

    \I__5182\ : InMux
    port map (
            O => \N__24563\,
            I => \N__24521\
        );

    \I__5181\ : InMux
    port map (
            O => \N__24560\,
            I => \N__24518\
        );

    \I__5180\ : InMux
    port map (
            O => \N__24557\,
            I => \N__24515\
        );

    \I__5179\ : InMux
    port map (
            O => \N__24554\,
            I => \N__24512\
        );

    \I__5178\ : InMux
    port map (
            O => \N__24551\,
            I => \N__24509\
        );

    \I__5177\ : InMux
    port map (
            O => \N__24548\,
            I => \N__24506\
        );

    \I__5176\ : InMux
    port map (
            O => \N__24545\,
            I => \N__24503\
        );

    \I__5175\ : InMux
    port map (
            O => \N__24542\,
            I => \N__24500\
        );

    \I__5174\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24497\
        );

    \I__5173\ : InMux
    port map (
            O => \N__24536\,
            I => \N__24494\
        );

    \I__5172\ : Span12Mux_h
    port map (
            O => \N__24533\,
            I => \N__24489\
        );

    \I__5171\ : Sp12to4
    port map (
            O => \N__24530\,
            I => \N__24484\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__24527\,
            I => \N__24484\
        );

    \I__5169\ : Span12Mux_v
    port map (
            O => \N__24524\,
            I => \N__24469\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__24521\,
            I => \N__24469\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__24518\,
            I => \N__24469\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__24515\,
            I => \N__24469\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__24512\,
            I => \N__24469\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__24509\,
            I => \N__24469\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__24506\,
            I => \N__24469\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__24503\,
            I => \N__24460\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__24500\,
            I => \N__24460\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__24497\,
            I => \N__24460\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__24494\,
            I => \N__24460\
        );

    \I__5158\ : CascadeMux
    port map (
            O => \N__24493\,
            I => \N__24456\
        );

    \I__5157\ : InMux
    port map (
            O => \N__24492\,
            I => \N__24452\
        );

    \I__5156\ : Span12Mux_v
    port map (
            O => \N__24489\,
            I => \N__24449\
        );

    \I__5155\ : Span12Mux_h
    port map (
            O => \N__24484\,
            I => \N__24446\
        );

    \I__5154\ : Span12Mux_v
    port map (
            O => \N__24469\,
            I => \N__24441\
        );

    \I__5153\ : Span12Mux_s7_v
    port map (
            O => \N__24460\,
            I => \N__24441\
        );

    \I__5152\ : InMux
    port map (
            O => \N__24459\,
            I => \N__24438\
        );

    \I__5151\ : InMux
    port map (
            O => \N__24456\,
            I => \N__24435\
        );

    \I__5150\ : InMux
    port map (
            O => \N__24455\,
            I => \N__24432\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__24452\,
            I => \N__24429\
        );

    \I__5148\ : Odrv12
    port map (
            O => \N__24449\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5147\ : Odrv12
    port map (
            O => \N__24446\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5146\ : Odrv12
    port map (
            O => \N__24441\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__24438\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__24435\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__24432\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__24429\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5141\ : InMux
    port map (
            O => \N__24414\,
            I => \N__24410\
        );

    \I__5140\ : InMux
    port map (
            O => \N__24413\,
            I => \N__24407\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__24410\,
            I => \N__24402\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__24407\,
            I => \N__24402\
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__24402\,
            I => \un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0\
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__24399\,
            I => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_10_cascade_\
        );

    \I__5135\ : InMux
    port map (
            O => \N__24396\,
            I => \N__24393\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__24393\,
            I => \N_612\
        );

    \I__5133\ : CascadeMux
    port map (
            O => \N__24390\,
            I => \N__24387\
        );

    \I__5132\ : InMux
    port map (
            O => \N__24387\,
            I => \N__24384\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__24384\,
            I => \N__24381\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__24381\,
            I => \this_ppu.un1_M_haddress_q_2_4\
        );

    \I__5129\ : InMux
    port map (
            O => \N__24378\,
            I => \N__24375\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__24375\,
            I => \N_627\
        );

    \I__5127\ : CascadeMux
    port map (
            O => \N__24372\,
            I => \N_509_0_cascade_\
        );

    \I__5126\ : CascadeMux
    port map (
            O => \N__24369\,
            I => \N__24363\
        );

    \I__5125\ : CascadeMux
    port map (
            O => \N__24368\,
            I => \N__24360\
        );

    \I__5124\ : CascadeMux
    port map (
            O => \N__24367\,
            I => \N__24355\
        );

    \I__5123\ : InMux
    port map (
            O => \N__24366\,
            I => \N__24352\
        );

    \I__5122\ : InMux
    port map (
            O => \N__24363\,
            I => \N__24349\
        );

    \I__5121\ : InMux
    port map (
            O => \N__24360\,
            I => \N__24346\
        );

    \I__5120\ : InMux
    port map (
            O => \N__24359\,
            I => \N__24342\
        );

    \I__5119\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24337\
        );

    \I__5118\ : InMux
    port map (
            O => \N__24355\,
            I => \N__24337\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__24352\,
            I => \N__24334\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__24349\,
            I => \N__24329\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__24346\,
            I => \N__24329\
        );

    \I__5114\ : InMux
    port map (
            O => \N__24345\,
            I => \N__24326\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__24342\,
            I => \N__24323\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__24337\,
            I => \N__24320\
        );

    \I__5111\ : Span4Mux_h
    port map (
            O => \N__24334\,
            I => \N__24313\
        );

    \I__5110\ : Span4Mux_v
    port map (
            O => \N__24329\,
            I => \N__24313\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__24326\,
            I => \N__24313\
        );

    \I__5108\ : Odrv4
    port map (
            O => \N__24323\,
            I => \this_vga_signals.N_415_0\
        );

    \I__5107\ : Odrv4
    port map (
            O => \N__24320\,
            I => \this_vga_signals.N_415_0\
        );

    \I__5106\ : Odrv4
    port map (
            O => \N__24313\,
            I => \this_vga_signals.N_415_0\
        );

    \I__5105\ : InMux
    port map (
            O => \N__24306\,
            I => \N__24300\
        );

    \I__5104\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24300\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__24300\,
            I => \N__24297\
        );

    \I__5102\ : Odrv4
    port map (
            O => \N__24297\,
            I => \un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0\
        );

    \I__5101\ : InMux
    port map (
            O => \N__24294\,
            I => \N__24291\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__24291\,
            I => \M_this_sprites_address_q_0_0_i_472\
        );

    \I__5099\ : InMux
    port map (
            O => \N__24288\,
            I => \N__24285\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__24285\,
            I => \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_6\
        );

    \I__5097\ : InMux
    port map (
            O => \N__24282\,
            I => \N__24276\
        );

    \I__5096\ : CascadeMux
    port map (
            O => \N__24281\,
            I => \N__24272\
        );

    \I__5095\ : CascadeMux
    port map (
            O => \N__24280\,
            I => \N__24269\
        );

    \I__5094\ : InMux
    port map (
            O => \N__24279\,
            I => \N__24265\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__24276\,
            I => \N__24262\
        );

    \I__5092\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24259\
        );

    \I__5091\ : InMux
    port map (
            O => \N__24272\,
            I => \N__24254\
        );

    \I__5090\ : InMux
    port map (
            O => \N__24269\,
            I => \N__24254\
        );

    \I__5089\ : InMux
    port map (
            O => \N__24268\,
            I => \N__24251\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__24265\,
            I => \N_773\
        );

    \I__5087\ : Odrv4
    port map (
            O => \N__24262\,
            I => \N_773\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__24259\,
            I => \N_773\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__24254\,
            I => \N_773\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__24251\,
            I => \N_773\
        );

    \I__5083\ : CascadeMux
    port map (
            O => \N__24240\,
            I => \N__24229\
        );

    \I__5082\ : CascadeMux
    port map (
            O => \N__24239\,
            I => \N__24226\
        );

    \I__5081\ : CascadeMux
    port map (
            O => \N__24238\,
            I => \N__24219\
        );

    \I__5080\ : CascadeMux
    port map (
            O => \N__24237\,
            I => \N__24216\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__24236\,
            I => \N__24213\
        );

    \I__5078\ : CascadeMux
    port map (
            O => \N__24235\,
            I => \N__24210\
        );

    \I__5077\ : CascadeMux
    port map (
            O => \N__24234\,
            I => \N__24207\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__24233\,
            I => \N__24202\
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__24232\,
            I => \N__24199\
        );

    \I__5074\ : InMux
    port map (
            O => \N__24229\,
            I => \N__24196\
        );

    \I__5073\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24193\
        );

    \I__5072\ : CascadeMux
    port map (
            O => \N__24225\,
            I => \N__24190\
        );

    \I__5071\ : CascadeMux
    port map (
            O => \N__24224\,
            I => \N__24187\
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__24223\,
            I => \N__24184\
        );

    \I__5069\ : CascadeMux
    port map (
            O => \N__24222\,
            I => \N__24181\
        );

    \I__5068\ : InMux
    port map (
            O => \N__24219\,
            I => \N__24178\
        );

    \I__5067\ : InMux
    port map (
            O => \N__24216\,
            I => \N__24175\
        );

    \I__5066\ : InMux
    port map (
            O => \N__24213\,
            I => \N__24172\
        );

    \I__5065\ : InMux
    port map (
            O => \N__24210\,
            I => \N__24169\
        );

    \I__5064\ : InMux
    port map (
            O => \N__24207\,
            I => \N__24166\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__24206\,
            I => \N__24163\
        );

    \I__5062\ : CascadeMux
    port map (
            O => \N__24205\,
            I => \N__24160\
        );

    \I__5061\ : InMux
    port map (
            O => \N__24202\,
            I => \N__24157\
        );

    \I__5060\ : InMux
    port map (
            O => \N__24199\,
            I => \N__24154\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__24196\,
            I => \N__24150\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__24193\,
            I => \N__24146\
        );

    \I__5057\ : InMux
    port map (
            O => \N__24190\,
            I => \N__24143\
        );

    \I__5056\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24140\
        );

    \I__5055\ : InMux
    port map (
            O => \N__24184\,
            I => \N__24137\
        );

    \I__5054\ : InMux
    port map (
            O => \N__24181\,
            I => \N__24134\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__24178\,
            I => \N__24129\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__24175\,
            I => \N__24129\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__24172\,
            I => \N__24126\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__24169\,
            I => \N__24121\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__24166\,
            I => \N__24121\
        );

    \I__5048\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24118\
        );

    \I__5047\ : InMux
    port map (
            O => \N__24160\,
            I => \N__24115\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__24157\,
            I => \N__24110\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__24154\,
            I => \N__24110\
        );

    \I__5044\ : CascadeMux
    port map (
            O => \N__24153\,
            I => \N__24105\
        );

    \I__5043\ : Span4Mux_h
    port map (
            O => \N__24150\,
            I => \N__24102\
        );

    \I__5042\ : CascadeMux
    port map (
            O => \N__24149\,
            I => \N__24099\
        );

    \I__5041\ : Span4Mux_v
    port map (
            O => \N__24146\,
            I => \N__24092\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__24143\,
            I => \N__24092\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__24140\,
            I => \N__24092\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__24137\,
            I => \N__24089\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__24134\,
            I => \N__24086\
        );

    \I__5036\ : Span4Mux_v
    port map (
            O => \N__24129\,
            I => \N__24081\
        );

    \I__5035\ : Span4Mux_v
    port map (
            O => \N__24126\,
            I => \N__24081\
        );

    \I__5034\ : Span4Mux_v
    port map (
            O => \N__24121\,
            I => \N__24072\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__24118\,
            I => \N__24072\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__24115\,
            I => \N__24072\
        );

    \I__5031\ : Span4Mux_v
    port map (
            O => \N__24110\,
            I => \N__24072\
        );

    \I__5030\ : CascadeMux
    port map (
            O => \N__24109\,
            I => \N__24068\
        );

    \I__5029\ : InMux
    port map (
            O => \N__24108\,
            I => \N__24063\
        );

    \I__5028\ : InMux
    port map (
            O => \N__24105\,
            I => \N__24063\
        );

    \I__5027\ : Span4Mux_h
    port map (
            O => \N__24102\,
            I => \N__24060\
        );

    \I__5026\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24057\
        );

    \I__5025\ : Sp12to4
    port map (
            O => \N__24092\,
            I => \N__24050\
        );

    \I__5024\ : Sp12to4
    port map (
            O => \N__24089\,
            I => \N__24050\
        );

    \I__5023\ : Sp12to4
    port map (
            O => \N__24086\,
            I => \N__24050\
        );

    \I__5022\ : Sp12to4
    port map (
            O => \N__24081\,
            I => \N__24047\
        );

    \I__5021\ : Sp12to4
    port map (
            O => \N__24072\,
            I => \N__24044\
        );

    \I__5020\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24041\
        );

    \I__5019\ : InMux
    port map (
            O => \N__24068\,
            I => \N__24038\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__24063\,
            I => \N__24035\
        );

    \I__5017\ : Span4Mux_h
    port map (
            O => \N__24060\,
            I => \N__24032\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__24057\,
            I => \N__24023\
        );

    \I__5015\ : Span12Mux_s8_v
    port map (
            O => \N__24050\,
            I => \N__24023\
        );

    \I__5014\ : Span12Mux_h
    port map (
            O => \N__24047\,
            I => \N__24023\
        );

    \I__5013\ : Span12Mux_v
    port map (
            O => \N__24044\,
            I => \N__24023\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__24041\,
            I => \N__24020\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__24038\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__5010\ : Odrv4
    port map (
            O => \N__24035\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__5009\ : Odrv4
    port map (
            O => \N__24032\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__5008\ : Odrv12
    port map (
            O => \N__24023\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__24020\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__5006\ : InMux
    port map (
            O => \N__24009\,
            I => \N__24006\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__24006\,
            I => \M_this_sprites_address_qc_6_0\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__24003\,
            I => \N__24000\
        );

    \I__5003\ : InMux
    port map (
            O => \N__24000\,
            I => \N__23997\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__23997\,
            I => \N__23994\
        );

    \I__5001\ : Odrv4
    port map (
            O => \N__23994\,
            I => \N_1282_tz_0\
        );

    \I__5000\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23987\
        );

    \I__4999\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23984\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__23987\,
            I => \un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__23984\,
            I => \un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0\
        );

    \I__4996\ : CascadeMux
    port map (
            O => \N__23979\,
            I => \N_1290_tz_0_cascade_\
        );

    \I__4995\ : InMux
    port map (
            O => \N__23976\,
            I => \N__23973\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__23973\,
            I => \N_607\
        );

    \I__4993\ : CascadeMux
    port map (
            O => \N__23970\,
            I => \N__23965\
        );

    \I__4992\ : CascadeMux
    port map (
            O => \N__23969\,
            I => \N__23958\
        );

    \I__4991\ : CascadeMux
    port map (
            O => \N__23968\,
            I => \N__23955\
        );

    \I__4990\ : InMux
    port map (
            O => \N__23965\,
            I => \N__23951\
        );

    \I__4989\ : CascadeMux
    port map (
            O => \N__23964\,
            I => \N__23948\
        );

    \I__4988\ : CascadeMux
    port map (
            O => \N__23963\,
            I => \N__23943\
        );

    \I__4987\ : CascadeMux
    port map (
            O => \N__23962\,
            I => \N__23939\
        );

    \I__4986\ : CascadeMux
    port map (
            O => \N__23961\,
            I => \N__23934\
        );

    \I__4985\ : InMux
    port map (
            O => \N__23958\,
            I => \N__23931\
        );

    \I__4984\ : InMux
    port map (
            O => \N__23955\,
            I => \N__23928\
        );

    \I__4983\ : CascadeMux
    port map (
            O => \N__23954\,
            I => \N__23925\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__23951\,
            I => \N__23922\
        );

    \I__4981\ : InMux
    port map (
            O => \N__23948\,
            I => \N__23919\
        );

    \I__4980\ : CascadeMux
    port map (
            O => \N__23947\,
            I => \N__23916\
        );

    \I__4979\ : CascadeMux
    port map (
            O => \N__23946\,
            I => \N__23913\
        );

    \I__4978\ : InMux
    port map (
            O => \N__23943\,
            I => \N__23910\
        );

    \I__4977\ : CascadeMux
    port map (
            O => \N__23942\,
            I => \N__23907\
        );

    \I__4976\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23903\
        );

    \I__4975\ : CascadeMux
    port map (
            O => \N__23938\,
            I => \N__23900\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__23937\,
            I => \N__23897\
        );

    \I__4973\ : InMux
    port map (
            O => \N__23934\,
            I => \N__23894\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__23931\,
            I => \N__23890\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__23928\,
            I => \N__23887\
        );

    \I__4970\ : InMux
    port map (
            O => \N__23925\,
            I => \N__23884\
        );

    \I__4969\ : Span4Mux_h
    port map (
            O => \N__23922\,
            I => \N__23880\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__23919\,
            I => \N__23877\
        );

    \I__4967\ : InMux
    port map (
            O => \N__23916\,
            I => \N__23874\
        );

    \I__4966\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23871\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__23910\,
            I => \N__23868\
        );

    \I__4964\ : InMux
    port map (
            O => \N__23907\,
            I => \N__23865\
        );

    \I__4963\ : CascadeMux
    port map (
            O => \N__23906\,
            I => \N__23862\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__23903\,
            I => \N__23859\
        );

    \I__4961\ : InMux
    port map (
            O => \N__23900\,
            I => \N__23856\
        );

    \I__4960\ : InMux
    port map (
            O => \N__23897\,
            I => \N__23853\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__23894\,
            I => \N__23850\
        );

    \I__4958\ : CascadeMux
    port map (
            O => \N__23893\,
            I => \N__23847\
        );

    \I__4957\ : Span4Mux_s2_v
    port map (
            O => \N__23890\,
            I => \N__23840\
        );

    \I__4956\ : Span4Mux_h
    port map (
            O => \N__23887\,
            I => \N__23840\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__23884\,
            I => \N__23840\
        );

    \I__4954\ : CascadeMux
    port map (
            O => \N__23883\,
            I => \N__23837\
        );

    \I__4953\ : Span4Mux_v
    port map (
            O => \N__23880\,
            I => \N__23832\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__23877\,
            I => \N__23832\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__23874\,
            I => \N__23829\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__23871\,
            I => \N__23826\
        );

    \I__4949\ : Span4Mux_h
    port map (
            O => \N__23868\,
            I => \N__23821\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__23865\,
            I => \N__23821\
        );

    \I__4947\ : InMux
    port map (
            O => \N__23862\,
            I => \N__23818\
        );

    \I__4946\ : Span4Mux_h
    port map (
            O => \N__23859\,
            I => \N__23815\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__23856\,
            I => \N__23812\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__23853\,
            I => \N__23808\
        );

    \I__4943\ : Span4Mux_v
    port map (
            O => \N__23850\,
            I => \N__23805\
        );

    \I__4942\ : InMux
    port map (
            O => \N__23847\,
            I => \N__23802\
        );

    \I__4941\ : Span4Mux_v
    port map (
            O => \N__23840\,
            I => \N__23799\
        );

    \I__4940\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23796\
        );

    \I__4939\ : Span4Mux_v
    port map (
            O => \N__23832\,
            I => \N__23791\
        );

    \I__4938\ : Span4Mux_h
    port map (
            O => \N__23829\,
            I => \N__23791\
        );

    \I__4937\ : Span4Mux_v
    port map (
            O => \N__23826\,
            I => \N__23784\
        );

    \I__4936\ : Span4Mux_v
    port map (
            O => \N__23821\,
            I => \N__23784\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__23818\,
            I => \N__23784\
        );

    \I__4934\ : Span4Mux_v
    port map (
            O => \N__23815\,
            I => \N__23777\
        );

    \I__4933\ : Span4Mux_h
    port map (
            O => \N__23812\,
            I => \N__23777\
        );

    \I__4932\ : InMux
    port map (
            O => \N__23811\,
            I => \N__23774\
        );

    \I__4931\ : Span12Mux_h
    port map (
            O => \N__23808\,
            I => \N__23771\
        );

    \I__4930\ : Sp12to4
    port map (
            O => \N__23805\,
            I => \N__23766\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__23802\,
            I => \N__23766\
        );

    \I__4928\ : Sp12to4
    port map (
            O => \N__23799\,
            I => \N__23761\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__23796\,
            I => \N__23761\
        );

    \I__4926\ : Span4Mux_h
    port map (
            O => \N__23791\,
            I => \N__23758\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__23784\,
            I => \N__23755\
        );

    \I__4924\ : CascadeMux
    port map (
            O => \N__23783\,
            I => \N__23752\
        );

    \I__4923\ : CascadeMux
    port map (
            O => \N__23782\,
            I => \N__23749\
        );

    \I__4922\ : Span4Mux_h
    port map (
            O => \N__23777\,
            I => \N__23743\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__23774\,
            I => \N__23743\
        );

    \I__4920\ : Span12Mux_v
    port map (
            O => \N__23771\,
            I => \N__23740\
        );

    \I__4919\ : Span12Mux_h
    port map (
            O => \N__23766\,
            I => \N__23735\
        );

    \I__4918\ : Span12Mux_h
    port map (
            O => \N__23761\,
            I => \N__23735\
        );

    \I__4917\ : Span4Mux_h
    port map (
            O => \N__23758\,
            I => \N__23730\
        );

    \I__4916\ : Span4Mux_h
    port map (
            O => \N__23755\,
            I => \N__23730\
        );

    \I__4915\ : InMux
    port map (
            O => \N__23752\,
            I => \N__23725\
        );

    \I__4914\ : InMux
    port map (
            O => \N__23749\,
            I => \N__23725\
        );

    \I__4913\ : InMux
    port map (
            O => \N__23748\,
            I => \N__23722\
        );

    \I__4912\ : Span4Mux_h
    port map (
            O => \N__23743\,
            I => \N__23719\
        );

    \I__4911\ : Odrv12
    port map (
            O => \N__23740\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__4910\ : Odrv12
    port map (
            O => \N__23735\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__23730\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__23725\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__23722\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__4906\ : Odrv4
    port map (
            O => \N__23719\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__4905\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23700\
        );

    \I__4904\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23700\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__23700\,
            I => \N__23697\
        );

    \I__4902\ : Span4Mux_h
    port map (
            O => \N__23697\,
            I => \N__23694\
        );

    \I__4901\ : Odrv4
    port map (
            O => \N__23694\,
            I => \un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0\
        );

    \I__4900\ : InMux
    port map (
            O => \N__23691\,
            I => \un1_M_this_sprites_address_q_cry_6\
        );

    \I__4899\ : CascadeMux
    port map (
            O => \N__23688\,
            I => \N__23684\
        );

    \I__4898\ : CascadeMux
    port map (
            O => \N__23687\,
            I => \N__23678\
        );

    \I__4897\ : InMux
    port map (
            O => \N__23684\,
            I => \N__23674\
        );

    \I__4896\ : CascadeMux
    port map (
            O => \N__23683\,
            I => \N__23671\
        );

    \I__4895\ : CascadeMux
    port map (
            O => \N__23682\,
            I => \N__23668\
        );

    \I__4894\ : CascadeMux
    port map (
            O => \N__23681\,
            I => \N__23661\
        );

    \I__4893\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23658\
        );

    \I__4892\ : CascadeMux
    port map (
            O => \N__23677\,
            I => \N__23655\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__23674\,
            I => \N__23650\
        );

    \I__4890\ : InMux
    port map (
            O => \N__23671\,
            I => \N__23647\
        );

    \I__4889\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23644\
        );

    \I__4888\ : CascadeMux
    port map (
            O => \N__23667\,
            I => \N__23641\
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__23666\,
            I => \N__23638\
        );

    \I__4886\ : CascadeMux
    port map (
            O => \N__23665\,
            I => \N__23633\
        );

    \I__4885\ : CascadeMux
    port map (
            O => \N__23664\,
            I => \N__23630\
        );

    \I__4884\ : InMux
    port map (
            O => \N__23661\,
            I => \N__23625\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__23658\,
            I => \N__23622\
        );

    \I__4882\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23619\
        );

    \I__4881\ : CascadeMux
    port map (
            O => \N__23654\,
            I => \N__23616\
        );

    \I__4880\ : CascadeMux
    port map (
            O => \N__23653\,
            I => \N__23613\
        );

    \I__4879\ : Span4Mux_v
    port map (
            O => \N__23650\,
            I => \N__23606\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__23647\,
            I => \N__23606\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__23644\,
            I => \N__23606\
        );

    \I__4876\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23603\
        );

    \I__4875\ : InMux
    port map (
            O => \N__23638\,
            I => \N__23600\
        );

    \I__4874\ : CascadeMux
    port map (
            O => \N__23637\,
            I => \N__23597\
        );

    \I__4873\ : CascadeMux
    port map (
            O => \N__23636\,
            I => \N__23594\
        );

    \I__4872\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23591\
        );

    \I__4871\ : InMux
    port map (
            O => \N__23630\,
            I => \N__23588\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__23629\,
            I => \N__23585\
        );

    \I__4869\ : CascadeMux
    port map (
            O => \N__23628\,
            I => \N__23582\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__23625\,
            I => \N__23579\
        );

    \I__4867\ : Span4Mux_h
    port map (
            O => \N__23622\,
            I => \N__23574\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__23619\,
            I => \N__23574\
        );

    \I__4865\ : InMux
    port map (
            O => \N__23616\,
            I => \N__23571\
        );

    \I__4864\ : InMux
    port map (
            O => \N__23613\,
            I => \N__23568\
        );

    \I__4863\ : Span4Mux_v
    port map (
            O => \N__23606\,
            I => \N__23561\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__23603\,
            I => \N__23561\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__23600\,
            I => \N__23561\
        );

    \I__4860\ : InMux
    port map (
            O => \N__23597\,
            I => \N__23558\
        );

    \I__4859\ : InMux
    port map (
            O => \N__23594\,
            I => \N__23555\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__23591\,
            I => \N__23550\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__23588\,
            I => \N__23550\
        );

    \I__4856\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23547\
        );

    \I__4855\ : InMux
    port map (
            O => \N__23582\,
            I => \N__23544\
        );

    \I__4854\ : Span4Mux_v
    port map (
            O => \N__23579\,
            I => \N__23537\
        );

    \I__4853\ : Span4Mux_v
    port map (
            O => \N__23574\,
            I => \N__23537\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__23571\,
            I => \N__23537\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__23568\,
            I => \N__23533\
        );

    \I__4850\ : Span4Mux_v
    port map (
            O => \N__23561\,
            I => \N__23526\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__23558\,
            I => \N__23526\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__23555\,
            I => \N__23526\
        );

    \I__4847\ : Span4Mux_v
    port map (
            O => \N__23550\,
            I => \N__23519\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__23547\,
            I => \N__23519\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__23544\,
            I => \N__23519\
        );

    \I__4844\ : Span4Mux_h
    port map (
            O => \N__23537\,
            I => \N__23514\
        );

    \I__4843\ : CascadeMux
    port map (
            O => \N__23536\,
            I => \N__23511\
        );

    \I__4842\ : Sp12to4
    port map (
            O => \N__23533\,
            I => \N__23507\
        );

    \I__4841\ : Span4Mux_v
    port map (
            O => \N__23526\,
            I => \N__23502\
        );

    \I__4840\ : Span4Mux_v
    port map (
            O => \N__23519\,
            I => \N__23502\
        );

    \I__4839\ : InMux
    port map (
            O => \N__23518\,
            I => \N__23499\
        );

    \I__4838\ : InMux
    port map (
            O => \N__23517\,
            I => \N__23496\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__23514\,
            I => \N__23493\
        );

    \I__4836\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23490\
        );

    \I__4835\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23487\
        );

    \I__4834\ : Span12Mux_s9_v
    port map (
            O => \N__23507\,
            I => \N__23478\
        );

    \I__4833\ : Sp12to4
    port map (
            O => \N__23502\,
            I => \N__23478\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__23499\,
            I => \N__23478\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__23496\,
            I => \N__23478\
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__23493\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__23490\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__23487\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__4827\ : Odrv12
    port map (
            O => \N__23478\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__4826\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23463\
        );

    \I__4825\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23463\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__23463\,
            I => \N__23460\
        );

    \I__4823\ : Odrv12
    port map (
            O => \N__23460\,
            I => \un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0\
        );

    \I__4822\ : InMux
    port map (
            O => \N__23457\,
            I => \bfn_19_23_0_\
        );

    \I__4821\ : InMux
    port map (
            O => \N__23454\,
            I => \un1_M_this_sprites_address_q_cry_8\
        );

    \I__4820\ : InMux
    port map (
            O => \N__23451\,
            I => \un1_M_this_sprites_address_q_cry_9\
        );

    \I__4819\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23445\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__23445\,
            I => \N__23441\
        );

    \I__4817\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23438\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__23441\,
            I => \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__23438\,
            I => \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\
        );

    \I__4814\ : InMux
    port map (
            O => \N__23433\,
            I => \un1_M_this_sprites_address_q_cry_10\
        );

    \I__4813\ : InMux
    port map (
            O => \N__23430\,
            I => \un1_M_this_sprites_address_q_cry_11\
        );

    \I__4812\ : InMux
    port map (
            O => \N__23427\,
            I => \un1_M_this_sprites_address_q_cry_12\
        );

    \I__4811\ : CascadeMux
    port map (
            O => \N__23424\,
            I => \N__23421\
        );

    \I__4810\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23418\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__23418\,
            I => \N__23415\
        );

    \I__4808\ : Span4Mux_v
    port map (
            O => \N__23415\,
            I => \N__23412\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__23412\,
            I => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_9\
        );

    \I__4806\ : CascadeMux
    port map (
            O => \N__23409\,
            I => \N__23406\
        );

    \I__4805\ : InMux
    port map (
            O => \N__23406\,
            I => \N__23403\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__23403\,
            I => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_13\
        );

    \I__4803\ : InMux
    port map (
            O => \N__23400\,
            I => \N__23396\
        );

    \I__4802\ : InMux
    port map (
            O => \N__23399\,
            I => \N__23393\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__23396\,
            I => \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__23393\,
            I => \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\
        );

    \I__4799\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23385\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__23385\,
            I => \this_vga_signals.N_459_0\
        );

    \I__4797\ : InMux
    port map (
            O => \N__23382\,
            I => \N__23378\
        );

    \I__4796\ : CascadeMux
    port map (
            O => \N__23381\,
            I => \N__23374\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__23378\,
            I => \N__23371\
        );

    \I__4794\ : InMux
    port map (
            O => \N__23377\,
            I => \N__23368\
        );

    \I__4793\ : InMux
    port map (
            O => \N__23374\,
            I => \N__23365\
        );

    \I__4792\ : Span4Mux_v
    port map (
            O => \N__23371\,
            I => \N__23362\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__23368\,
            I => \N_440_0\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__23365\,
            I => \N_440_0\
        );

    \I__4789\ : Odrv4
    port map (
            O => \N__23362\,
            I => \N_440_0\
        );

    \I__4788\ : CascadeMux
    port map (
            O => \N__23355\,
            I => \N__23348\
        );

    \I__4787\ : CascadeMux
    port map (
            O => \N__23354\,
            I => \N__23345\
        );

    \I__4786\ : CascadeMux
    port map (
            O => \N__23353\,
            I => \N__23342\
        );

    \I__4785\ : CascadeMux
    port map (
            O => \N__23352\,
            I => \N__23338\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__23351\,
            I => \N__23331\
        );

    \I__4783\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23324\
        );

    \I__4782\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23321\
        );

    \I__4781\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23318\
        );

    \I__4780\ : CascadeMux
    port map (
            O => \N__23341\,
            I => \N__23314\
        );

    \I__4779\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23311\
        );

    \I__4778\ : CascadeMux
    port map (
            O => \N__23337\,
            I => \N__23308\
        );

    \I__4777\ : CascadeMux
    port map (
            O => \N__23336\,
            I => \N__23304\
        );

    \I__4776\ : CascadeMux
    port map (
            O => \N__23335\,
            I => \N__23301\
        );

    \I__4775\ : CascadeMux
    port map (
            O => \N__23334\,
            I => \N__23298\
        );

    \I__4774\ : InMux
    port map (
            O => \N__23331\,
            I => \N__23295\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__23330\,
            I => \N__23292\
        );

    \I__4772\ : CascadeMux
    port map (
            O => \N__23329\,
            I => \N__23289\
        );

    \I__4771\ : CascadeMux
    port map (
            O => \N__23328\,
            I => \N__23286\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__23327\,
            I => \N__23283\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__23324\,
            I => \N__23280\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__23321\,
            I => \N__23275\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__23318\,
            I => \N__23275\
        );

    \I__4766\ : CascadeMux
    port map (
            O => \N__23317\,
            I => \N__23272\
        );

    \I__4765\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23269\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__23311\,
            I => \N__23266\
        );

    \I__4763\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23263\
        );

    \I__4762\ : CascadeMux
    port map (
            O => \N__23307\,
            I => \N__23260\
        );

    \I__4761\ : InMux
    port map (
            O => \N__23304\,
            I => \N__23257\
        );

    \I__4760\ : InMux
    port map (
            O => \N__23301\,
            I => \N__23254\
        );

    \I__4759\ : InMux
    port map (
            O => \N__23298\,
            I => \N__23251\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__23295\,
            I => \N__23248\
        );

    \I__4757\ : InMux
    port map (
            O => \N__23292\,
            I => \N__23245\
        );

    \I__4756\ : InMux
    port map (
            O => \N__23289\,
            I => \N__23242\
        );

    \I__4755\ : InMux
    port map (
            O => \N__23286\,
            I => \N__23239\
        );

    \I__4754\ : InMux
    port map (
            O => \N__23283\,
            I => \N__23236\
        );

    \I__4753\ : Span4Mux_v
    port map (
            O => \N__23280\,
            I => \N__23231\
        );

    \I__4752\ : Span4Mux_v
    port map (
            O => \N__23275\,
            I => \N__23231\
        );

    \I__4751\ : InMux
    port map (
            O => \N__23272\,
            I => \N__23228\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__23269\,
            I => \N__23225\
        );

    \I__4749\ : Span4Mux_h
    port map (
            O => \N__23266\,
            I => \N__23220\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__23263\,
            I => \N__23220\
        );

    \I__4747\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23217\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__23257\,
            I => \N__23210\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__23254\,
            I => \N__23210\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23210\
        );

    \I__4743\ : Span12Mux_s7_h
    port map (
            O => \N__23248\,
            I => \N__23199\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__23245\,
            I => \N__23199\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__23242\,
            I => \N__23199\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__23239\,
            I => \N__23199\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__23236\,
            I => \N__23199\
        );

    \I__4738\ : Span4Mux_h
    port map (
            O => \N__23231\,
            I => \N__23196\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__23228\,
            I => \N__23193\
        );

    \I__4736\ : Span4Mux_v
    port map (
            O => \N__23225\,
            I => \N__23186\
        );

    \I__4735\ : Span4Mux_v
    port map (
            O => \N__23220\,
            I => \N__23186\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__23217\,
            I => \N__23186\
        );

    \I__4733\ : Span12Mux_s10_v
    port map (
            O => \N__23210\,
            I => \N__23172\
        );

    \I__4732\ : Span12Mux_v
    port map (
            O => \N__23199\,
            I => \N__23172\
        );

    \I__4731\ : Sp12to4
    port map (
            O => \N__23196\,
            I => \N__23172\
        );

    \I__4730\ : Span12Mux_h
    port map (
            O => \N__23193\,
            I => \N__23172\
        );

    \I__4729\ : Span4Mux_h
    port map (
            O => \N__23186\,
            I => \N__23169\
        );

    \I__4728\ : InMux
    port map (
            O => \N__23185\,
            I => \N__23166\
        );

    \I__4727\ : InMux
    port map (
            O => \N__23184\,
            I => \N__23163\
        );

    \I__4726\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23158\
        );

    \I__4725\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23158\
        );

    \I__4724\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23155\
        );

    \I__4723\ : Odrv12
    port map (
            O => \N__23172\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__4722\ : Odrv4
    port map (
            O => \N__23169\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__23166\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__23163\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__23158\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__23155\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__4717\ : CascadeMux
    port map (
            O => \N__23142\,
            I => \N__23138\
        );

    \I__4716\ : InMux
    port map (
            O => \N__23141\,
            I => \N__23135\
        );

    \I__4715\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23132\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__23135\,
            I => \un1_M_this_state_q_6_0\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__23132\,
            I => \un1_M_this_state_q_6_0\
        );

    \I__4712\ : InMux
    port map (
            O => \N__23127\,
            I => \N__23124\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__23124\,
            I => \N__23120\
        );

    \I__4710\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23117\
        );

    \I__4709\ : Odrv4
    port map (
            O => \N__23120\,
            I => \M_this_sprites_address_q_RNIRO0N6Z0Z_0\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__23117\,
            I => \M_this_sprites_address_q_RNIRO0N6Z0Z_0\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__23112\,
            I => \N__23105\
        );

    \I__4706\ : CascadeMux
    port map (
            O => \N__23111\,
            I => \N__23102\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__23110\,
            I => \N__23098\
        );

    \I__4704\ : CascadeMux
    port map (
            O => \N__23109\,
            I => \N__23095\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__23108\,
            I => \N__23090\
        );

    \I__4702\ : InMux
    port map (
            O => \N__23105\,
            I => \N__23084\
        );

    \I__4701\ : InMux
    port map (
            O => \N__23102\,
            I => \N__23081\
        );

    \I__4700\ : CascadeMux
    port map (
            O => \N__23101\,
            I => \N__23078\
        );

    \I__4699\ : InMux
    port map (
            O => \N__23098\,
            I => \N__23075\
        );

    \I__4698\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23072\
        );

    \I__4697\ : CascadeMux
    port map (
            O => \N__23094\,
            I => \N__23069\
        );

    \I__4696\ : CascadeMux
    port map (
            O => \N__23093\,
            I => \N__23066\
        );

    \I__4695\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23062\
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__23089\,
            I => \N__23059\
        );

    \I__4693\ : CascadeMux
    port map (
            O => \N__23088\,
            I => \N__23056\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__23087\,
            I => \N__23051\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__23084\,
            I => \N__23048\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__23081\,
            I => \N__23045\
        );

    \I__4689\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23042\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__23075\,
            I => \N__23039\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__23072\,
            I => \N__23036\
        );

    \I__4686\ : InMux
    port map (
            O => \N__23069\,
            I => \N__23033\
        );

    \I__4685\ : InMux
    port map (
            O => \N__23066\,
            I => \N__23030\
        );

    \I__4684\ : CascadeMux
    port map (
            O => \N__23065\,
            I => \N__23027\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__23062\,
            I => \N__23024\
        );

    \I__4682\ : InMux
    port map (
            O => \N__23059\,
            I => \N__23021\
        );

    \I__4681\ : InMux
    port map (
            O => \N__23056\,
            I => \N__23018\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__23055\,
            I => \N__23015\
        );

    \I__4679\ : CascadeMux
    port map (
            O => \N__23054\,
            I => \N__23012\
        );

    \I__4678\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23008\
        );

    \I__4677\ : Span4Mux_h
    port map (
            O => \N__23048\,
            I => \N__23001\
        );

    \I__4676\ : Span4Mux_v
    port map (
            O => \N__23045\,
            I => \N__23001\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__23042\,
            I => \N__23001\
        );

    \I__4674\ : Span4Mux_v
    port map (
            O => \N__23039\,
            I => \N__22994\
        );

    \I__4673\ : Span4Mux_h
    port map (
            O => \N__23036\,
            I => \N__22994\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__23033\,
            I => \N__22994\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__23030\,
            I => \N__22991\
        );

    \I__4670\ : InMux
    port map (
            O => \N__23027\,
            I => \N__22988\
        );

    \I__4669\ : Span4Mux_s2_v
    port map (
            O => \N__23024\,
            I => \N__22981\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__23021\,
            I => \N__22981\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__23018\,
            I => \N__22981\
        );

    \I__4666\ : InMux
    port map (
            O => \N__23015\,
            I => \N__22978\
        );

    \I__4665\ : InMux
    port map (
            O => \N__23012\,
            I => \N__22975\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__23011\,
            I => \N__22971\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__23008\,
            I => \N__22968\
        );

    \I__4662\ : Span4Mux_v
    port map (
            O => \N__23001\,
            I => \N__22965\
        );

    \I__4661\ : Span4Mux_v
    port map (
            O => \N__22994\,
            I => \N__22958\
        );

    \I__4660\ : Span4Mux_h
    port map (
            O => \N__22991\,
            I => \N__22958\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__22988\,
            I => \N__22958\
        );

    \I__4658\ : Span4Mux_v
    port map (
            O => \N__22981\,
            I => \N__22951\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__22978\,
            I => \N__22951\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__22975\,
            I => \N__22951\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__22974\,
            I => \N__22948\
        );

    \I__4654\ : InMux
    port map (
            O => \N__22971\,
            I => \N__22944\
        );

    \I__4653\ : Span12Mux_h
    port map (
            O => \N__22968\,
            I => \N__22941\
        );

    \I__4652\ : Sp12to4
    port map (
            O => \N__22965\,
            I => \N__22938\
        );

    \I__4651\ : Span4Mux_v
    port map (
            O => \N__22958\,
            I => \N__22933\
        );

    \I__4650\ : Span4Mux_v
    port map (
            O => \N__22951\,
            I => \N__22933\
        );

    \I__4649\ : InMux
    port map (
            O => \N__22948\,
            I => \N__22930\
        );

    \I__4648\ : InMux
    port map (
            O => \N__22947\,
            I => \N__22927\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__22944\,
            I => \N__22921\
        );

    \I__4646\ : Span12Mux_v
    port map (
            O => \N__22941\,
            I => \N__22912\
        );

    \I__4645\ : Span12Mux_h
    port map (
            O => \N__22938\,
            I => \N__22912\
        );

    \I__4644\ : Sp12to4
    port map (
            O => \N__22933\,
            I => \N__22912\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__22930\,
            I => \N__22912\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__22927\,
            I => \N__22909\
        );

    \I__4641\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22906\
        );

    \I__4640\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22903\
        );

    \I__4639\ : InMux
    port map (
            O => \N__22924\,
            I => \N__22900\
        );

    \I__4638\ : Odrv12
    port map (
            O => \N__22921\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__4637\ : Odrv12
    port map (
            O => \N__22912\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__22909\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__22906\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__22903\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__22900\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__4632\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22884\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__22884\,
            I => \N__22880\
        );

    \I__4630\ : InMux
    port map (
            O => \N__22883\,
            I => \N__22877\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__22880\,
            I => \un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__22877\,
            I => \un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0\
        );

    \I__4627\ : InMux
    port map (
            O => \N__22872\,
            I => \un1_M_this_sprites_address_q_cry_0\
        );

    \I__4626\ : CascadeMux
    port map (
            O => \N__22869\,
            I => \N__22865\
        );

    \I__4625\ : CascadeMux
    port map (
            O => \N__22868\,
            I => \N__22860\
        );

    \I__4624\ : InMux
    port map (
            O => \N__22865\,
            I => \N__22849\
        );

    \I__4623\ : CascadeMux
    port map (
            O => \N__22864\,
            I => \N__22846\
        );

    \I__4622\ : CascadeMux
    port map (
            O => \N__22863\,
            I => \N__22842\
        );

    \I__4621\ : InMux
    port map (
            O => \N__22860\,
            I => \N__22839\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__22859\,
            I => \N__22836\
        );

    \I__4619\ : CascadeMux
    port map (
            O => \N__22858\,
            I => \N__22833\
        );

    \I__4618\ : CascadeMux
    port map (
            O => \N__22857\,
            I => \N__22830\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__22856\,
            I => \N__22827\
        );

    \I__4616\ : CascadeMux
    port map (
            O => \N__22855\,
            I => \N__22824\
        );

    \I__4615\ : CascadeMux
    port map (
            O => \N__22854\,
            I => \N__22821\
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__22853\,
            I => \N__22818\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__22852\,
            I => \N__22814\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__22849\,
            I => \N__22811\
        );

    \I__4611\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22808\
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__22845\,
            I => \N__22805\
        );

    \I__4609\ : InMux
    port map (
            O => \N__22842\,
            I => \N__22802\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__22839\,
            I => \N__22797\
        );

    \I__4607\ : InMux
    port map (
            O => \N__22836\,
            I => \N__22794\
        );

    \I__4606\ : InMux
    port map (
            O => \N__22833\,
            I => \N__22791\
        );

    \I__4605\ : InMux
    port map (
            O => \N__22830\,
            I => \N__22788\
        );

    \I__4604\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22785\
        );

    \I__4603\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22782\
        );

    \I__4602\ : InMux
    port map (
            O => \N__22821\,
            I => \N__22779\
        );

    \I__4601\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22776\
        );

    \I__4600\ : CascadeMux
    port map (
            O => \N__22817\,
            I => \N__22772\
        );

    \I__4599\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22769\
        );

    \I__4598\ : Span4Mux_v
    port map (
            O => \N__22811\,
            I => \N__22764\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__22808\,
            I => \N__22764\
        );

    \I__4596\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22761\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__22802\,
            I => \N__22758\
        );

    \I__4594\ : CascadeMux
    port map (
            O => \N__22801\,
            I => \N__22755\
        );

    \I__4593\ : CascadeMux
    port map (
            O => \N__22800\,
            I => \N__22752\
        );

    \I__4592\ : Span4Mux_v
    port map (
            O => \N__22797\,
            I => \N__22745\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__22794\,
            I => \N__22745\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__22791\,
            I => \N__22745\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__22788\,
            I => \N__22742\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__22785\,
            I => \N__22737\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__22782\,
            I => \N__22737\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__22779\,
            I => \N__22732\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__22776\,
            I => \N__22732\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__22775\,
            I => \N__22729\
        );

    \I__4583\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22726\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__22769\,
            I => \N__22719\
        );

    \I__4581\ : Span4Mux_v
    port map (
            O => \N__22764\,
            I => \N__22719\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__22761\,
            I => \N__22719\
        );

    \I__4579\ : Span4Mux_v
    port map (
            O => \N__22758\,
            I => \N__22716\
        );

    \I__4578\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22713\
        );

    \I__4577\ : InMux
    port map (
            O => \N__22752\,
            I => \N__22710\
        );

    \I__4576\ : Span4Mux_v
    port map (
            O => \N__22745\,
            I => \N__22707\
        );

    \I__4575\ : Span4Mux_v
    port map (
            O => \N__22742\,
            I => \N__22704\
        );

    \I__4574\ : Span4Mux_v
    port map (
            O => \N__22737\,
            I => \N__22698\
        );

    \I__4573\ : Span4Mux_v
    port map (
            O => \N__22732\,
            I => \N__22698\
        );

    \I__4572\ : InMux
    port map (
            O => \N__22729\,
            I => \N__22695\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__22726\,
            I => \N__22692\
        );

    \I__4570\ : Span4Mux_v
    port map (
            O => \N__22719\,
            I => \N__22687\
        );

    \I__4569\ : Span4Mux_h
    port map (
            O => \N__22716\,
            I => \N__22684\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__22713\,
            I => \N__22681\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__22710\,
            I => \N__22674\
        );

    \I__4566\ : Sp12to4
    port map (
            O => \N__22707\,
            I => \N__22674\
        );

    \I__4565\ : Sp12to4
    port map (
            O => \N__22704\,
            I => \N__22674\
        );

    \I__4564\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22671\
        );

    \I__4563\ : Span4Mux_h
    port map (
            O => \N__22698\,
            I => \N__22668\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__22695\,
            I => \N__22665\
        );

    \I__4561\ : Span12Mux_h
    port map (
            O => \N__22692\,
            I => \N__22662\
        );

    \I__4560\ : InMux
    port map (
            O => \N__22691\,
            I => \N__22659\
        );

    \I__4559\ : InMux
    port map (
            O => \N__22690\,
            I => \N__22656\
        );

    \I__4558\ : Span4Mux_h
    port map (
            O => \N__22687\,
            I => \N__22651\
        );

    \I__4557\ : Span4Mux_v
    port map (
            O => \N__22684\,
            I => \N__22651\
        );

    \I__4556\ : Span12Mux_h
    port map (
            O => \N__22681\,
            I => \N__22646\
        );

    \I__4555\ : Span12Mux_h
    port map (
            O => \N__22674\,
            I => \N__22646\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__22671\,
            I => \N__22639\
        );

    \I__4553\ : Span4Mux_h
    port map (
            O => \N__22668\,
            I => \N__22639\
        );

    \I__4552\ : Span4Mux_v
    port map (
            O => \N__22665\,
            I => \N__22639\
        );

    \I__4551\ : Odrv12
    port map (
            O => \N__22662\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__22659\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__22656\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4548\ : Odrv4
    port map (
            O => \N__22651\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4547\ : Odrv12
    port map (
            O => \N__22646\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4546\ : Odrv4
    port map (
            O => \N__22639\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__4545\ : InMux
    port map (
            O => \N__22626\,
            I => \N__22620\
        );

    \I__4544\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22620\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__22620\,
            I => \N__22617\
        );

    \I__4542\ : Span4Mux_h
    port map (
            O => \N__22617\,
            I => \N__22614\
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__22614\,
            I => \un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0\
        );

    \I__4540\ : InMux
    port map (
            O => \N__22611\,
            I => \un1_M_this_sprites_address_q_cry_1\
        );

    \I__4539\ : CascadeMux
    port map (
            O => \N__22608\,
            I => \N__22605\
        );

    \I__4538\ : InMux
    port map (
            O => \N__22605\,
            I => \N__22599\
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__22604\,
            I => \N__22596\
        );

    \I__4536\ : CascadeMux
    port map (
            O => \N__22603\,
            I => \N__22593\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__22602\,
            I => \N__22588\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__22599\,
            I => \N__22583\
        );

    \I__4533\ : InMux
    port map (
            O => \N__22596\,
            I => \N__22580\
        );

    \I__4532\ : InMux
    port map (
            O => \N__22593\,
            I => \N__22577\
        );

    \I__4531\ : CascadeMux
    port map (
            O => \N__22592\,
            I => \N__22574\
        );

    \I__4530\ : CascadeMux
    port map (
            O => \N__22591\,
            I => \N__22571\
        );

    \I__4529\ : InMux
    port map (
            O => \N__22588\,
            I => \N__22566\
        );

    \I__4528\ : CascadeMux
    port map (
            O => \N__22587\,
            I => \N__22563\
        );

    \I__4527\ : CascadeMux
    port map (
            O => \N__22586\,
            I => \N__22560\
        );

    \I__4526\ : Span4Mux_h
    port map (
            O => \N__22583\,
            I => \N__22549\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__22580\,
            I => \N__22549\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__22577\,
            I => \N__22546\
        );

    \I__4523\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22543\
        );

    \I__4522\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22540\
        );

    \I__4521\ : CascadeMux
    port map (
            O => \N__22570\,
            I => \N__22537\
        );

    \I__4520\ : CascadeMux
    port map (
            O => \N__22569\,
            I => \N__22534\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__22566\,
            I => \N__22531\
        );

    \I__4518\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22528\
        );

    \I__4517\ : InMux
    port map (
            O => \N__22560\,
            I => \N__22525\
        );

    \I__4516\ : CascadeMux
    port map (
            O => \N__22559\,
            I => \N__22522\
        );

    \I__4515\ : CascadeMux
    port map (
            O => \N__22558\,
            I => \N__22519\
        );

    \I__4514\ : CascadeMux
    port map (
            O => \N__22557\,
            I => \N__22516\
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__22556\,
            I => \N__22513\
        );

    \I__4512\ : CascadeMux
    port map (
            O => \N__22555\,
            I => \N__22510\
        );

    \I__4511\ : CascadeMux
    port map (
            O => \N__22554\,
            I => \N__22507\
        );

    \I__4510\ : Span4Mux_v
    port map (
            O => \N__22549\,
            I => \N__22500\
        );

    \I__4509\ : Span4Mux_h
    port map (
            O => \N__22546\,
            I => \N__22500\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__22543\,
            I => \N__22500\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__22540\,
            I => \N__22497\
        );

    \I__4506\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22494\
        );

    \I__4505\ : InMux
    port map (
            O => \N__22534\,
            I => \N__22491\
        );

    \I__4504\ : Span4Mux_s2_v
    port map (
            O => \N__22531\,
            I => \N__22484\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__22528\,
            I => \N__22484\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__22525\,
            I => \N__22484\
        );

    \I__4501\ : InMux
    port map (
            O => \N__22522\,
            I => \N__22481\
        );

    \I__4500\ : InMux
    port map (
            O => \N__22519\,
            I => \N__22478\
        );

    \I__4499\ : InMux
    port map (
            O => \N__22516\,
            I => \N__22475\
        );

    \I__4498\ : InMux
    port map (
            O => \N__22513\,
            I => \N__22472\
        );

    \I__4497\ : InMux
    port map (
            O => \N__22510\,
            I => \N__22469\
        );

    \I__4496\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22466\
        );

    \I__4495\ : Span4Mux_v
    port map (
            O => \N__22500\,
            I => \N__22459\
        );

    \I__4494\ : Span4Mux_h
    port map (
            O => \N__22497\,
            I => \N__22459\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__22494\,
            I => \N__22459\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__22491\,
            I => \N__22456\
        );

    \I__4491\ : Span4Mux_v
    port map (
            O => \N__22484\,
            I => \N__22449\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__22481\,
            I => \N__22449\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__22478\,
            I => \N__22449\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__22475\,
            I => \N__22443\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__22472\,
            I => \N__22443\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__22469\,
            I => \N__22438\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__22466\,
            I => \N__22438\
        );

    \I__4484\ : Span4Mux_v
    port map (
            O => \N__22459\,
            I => \N__22431\
        );

    \I__4483\ : Span4Mux_h
    port map (
            O => \N__22456\,
            I => \N__22431\
        );

    \I__4482\ : Span4Mux_v
    port map (
            O => \N__22449\,
            I => \N__22431\
        );

    \I__4481\ : InMux
    port map (
            O => \N__22448\,
            I => \N__22428\
        );

    \I__4480\ : Span4Mux_v
    port map (
            O => \N__22443\,
            I => \N__22423\
        );

    \I__4479\ : Span4Mux_v
    port map (
            O => \N__22438\,
            I => \N__22423\
        );

    \I__4478\ : Span4Mux_h
    port map (
            O => \N__22431\,
            I => \N__22415\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__22428\,
            I => \N__22415\
        );

    \I__4476\ : Sp12to4
    port map (
            O => \N__22423\,
            I => \N__22412\
        );

    \I__4475\ : InMux
    port map (
            O => \N__22422\,
            I => \N__22407\
        );

    \I__4474\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22407\
        );

    \I__4473\ : InMux
    port map (
            O => \N__22420\,
            I => \N__22404\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__22415\,
            I => \N__22401\
        );

    \I__4471\ : Odrv12
    port map (
            O => \N__22412\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__22407\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__22404\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__22401\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__22392\,
            I => \N__22389\
        );

    \I__4466\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22386\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__22386\,
            I => \N__22382\
        );

    \I__4464\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22379\
        );

    \I__4463\ : Span4Mux_h
    port map (
            O => \N__22382\,
            I => \N__22376\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__22379\,
            I => \un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__22376\,
            I => \un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0\
        );

    \I__4460\ : InMux
    port map (
            O => \N__22371\,
            I => \un1_M_this_sprites_address_q_cry_2\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__22368\,
            I => \N__22362\
        );

    \I__4458\ : CascadeMux
    port map (
            O => \N__22367\,
            I => \N__22359\
        );

    \I__4457\ : CascadeMux
    port map (
            O => \N__22366\,
            I => \N__22353\
        );

    \I__4456\ : CascadeMux
    port map (
            O => \N__22365\,
            I => \N__22349\
        );

    \I__4455\ : InMux
    port map (
            O => \N__22362\,
            I => \N__22342\
        );

    \I__4454\ : InMux
    port map (
            O => \N__22359\,
            I => \N__22339\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__22358\,
            I => \N__22336\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__22357\,
            I => \N__22331\
        );

    \I__4451\ : CascadeMux
    port map (
            O => \N__22356\,
            I => \N__22328\
        );

    \I__4450\ : InMux
    port map (
            O => \N__22353\,
            I => \N__22325\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__22352\,
            I => \N__22322\
        );

    \I__4448\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22319\
        );

    \I__4447\ : CascadeMux
    port map (
            O => \N__22348\,
            I => \N__22316\
        );

    \I__4446\ : CascadeMux
    port map (
            O => \N__22347\,
            I => \N__22313\
        );

    \I__4445\ : CascadeMux
    port map (
            O => \N__22346\,
            I => \N__22310\
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__22345\,
            I => \N__22306\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__22342\,
            I => \N__22301\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__22339\,
            I => \N__22301\
        );

    \I__4441\ : InMux
    port map (
            O => \N__22336\,
            I => \N__22298\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__22335\,
            I => \N__22295\
        );

    \I__4439\ : CascadeMux
    port map (
            O => \N__22334\,
            I => \N__22292\
        );

    \I__4438\ : InMux
    port map (
            O => \N__22331\,
            I => \N__22289\
        );

    \I__4437\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22286\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__22325\,
            I => \N__22283\
        );

    \I__4435\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22280\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__22319\,
            I => \N__22276\
        );

    \I__4433\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22273\
        );

    \I__4432\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22270\
        );

    \I__4431\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22267\
        );

    \I__4430\ : CascadeMux
    port map (
            O => \N__22309\,
            I => \N__22264\
        );

    \I__4429\ : InMux
    port map (
            O => \N__22306\,
            I => \N__22261\
        );

    \I__4428\ : Span4Mux_v
    port map (
            O => \N__22301\,
            I => \N__22256\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__22298\,
            I => \N__22256\
        );

    \I__4426\ : InMux
    port map (
            O => \N__22295\,
            I => \N__22253\
        );

    \I__4425\ : InMux
    port map (
            O => \N__22292\,
            I => \N__22250\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__22289\,
            I => \N__22247\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__22286\,
            I => \N__22242\
        );

    \I__4422\ : Span4Mux_h
    port map (
            O => \N__22283\,
            I => \N__22242\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__22280\,
            I => \N__22239\
        );

    \I__4420\ : CascadeMux
    port map (
            O => \N__22279\,
            I => \N__22236\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__22276\,
            I => \N__22231\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__22273\,
            I => \N__22231\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22226\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__22267\,
            I => \N__22226\
        );

    \I__4415\ : InMux
    port map (
            O => \N__22264\,
            I => \N__22223\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__22261\,
            I => \N__22220\
        );

    \I__4413\ : Span4Mux_h
    port map (
            O => \N__22256\,
            I => \N__22217\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__22253\,
            I => \N__22212\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__22250\,
            I => \N__22212\
        );

    \I__4410\ : Span4Mux_v
    port map (
            O => \N__22247\,
            I => \N__22205\
        );

    \I__4409\ : Span4Mux_v
    port map (
            O => \N__22242\,
            I => \N__22205\
        );

    \I__4408\ : Span4Mux_h
    port map (
            O => \N__22239\,
            I => \N__22205\
        );

    \I__4407\ : InMux
    port map (
            O => \N__22236\,
            I => \N__22199\
        );

    \I__4406\ : Span4Mux_s2_v
    port map (
            O => \N__22231\,
            I => \N__22196\
        );

    \I__4405\ : Span4Mux_v
    port map (
            O => \N__22226\,
            I => \N__22189\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__22223\,
            I => \N__22189\
        );

    \I__4403\ : Span4Mux_v
    port map (
            O => \N__22220\,
            I => \N__22189\
        );

    \I__4402\ : Span4Mux_v
    port map (
            O => \N__22217\,
            I => \N__22186\
        );

    \I__4401\ : Span4Mux_v
    port map (
            O => \N__22212\,
            I => \N__22183\
        );

    \I__4400\ : Span4Mux_h
    port map (
            O => \N__22205\,
            I => \N__22180\
        );

    \I__4399\ : InMux
    port map (
            O => \N__22204\,
            I => \N__22177\
        );

    \I__4398\ : CascadeMux
    port map (
            O => \N__22203\,
            I => \N__22174\
        );

    \I__4397\ : CascadeMux
    port map (
            O => \N__22202\,
            I => \N__22171\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__22199\,
            I => \N__22165\
        );

    \I__4395\ : Sp12to4
    port map (
            O => \N__22196\,
            I => \N__22165\
        );

    \I__4394\ : Span4Mux_h
    port map (
            O => \N__22189\,
            I => \N__22160\
        );

    \I__4393\ : Span4Mux_v
    port map (
            O => \N__22186\,
            I => \N__22160\
        );

    \I__4392\ : Span4Mux_h
    port map (
            O => \N__22183\,
            I => \N__22153\
        );

    \I__4391\ : Span4Mux_h
    port map (
            O => \N__22180\,
            I => \N__22153\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__22177\,
            I => \N__22153\
        );

    \I__4389\ : InMux
    port map (
            O => \N__22174\,
            I => \N__22146\
        );

    \I__4388\ : InMux
    port map (
            O => \N__22171\,
            I => \N__22146\
        );

    \I__4387\ : InMux
    port map (
            O => \N__22170\,
            I => \N__22146\
        );

    \I__4386\ : Span12Mux_h
    port map (
            O => \N__22165\,
            I => \N__22143\
        );

    \I__4385\ : Span4Mux_h
    port map (
            O => \N__22160\,
            I => \N__22140\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__22153\,
            I => \N__22137\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__22146\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__4382\ : Odrv12
    port map (
            O => \N__22143\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__22140\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__22137\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__4379\ : InMux
    port map (
            O => \N__22128\,
            I => \N__22122\
        );

    \I__4378\ : InMux
    port map (
            O => \N__22127\,
            I => \N__22122\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__22122\,
            I => \N__22119\
        );

    \I__4376\ : Span4Mux_h
    port map (
            O => \N__22119\,
            I => \N__22116\
        );

    \I__4375\ : Odrv4
    port map (
            O => \N__22116\,
            I => \un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0\
        );

    \I__4374\ : InMux
    port map (
            O => \N__22113\,
            I => \un1_M_this_sprites_address_q_cry_3\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__22110\,
            I => \N__22107\
        );

    \I__4372\ : InMux
    port map (
            O => \N__22107\,
            I => \N__22103\
        );

    \I__4371\ : CascadeMux
    port map (
            O => \N__22106\,
            I => \N__22100\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__22103\,
            I => \N__22095\
        );

    \I__4369\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22092\
        );

    \I__4368\ : CascadeMux
    port map (
            O => \N__22099\,
            I => \N__22089\
        );

    \I__4367\ : CascadeMux
    port map (
            O => \N__22098\,
            I => \N__22085\
        );

    \I__4366\ : Span4Mux_h
    port map (
            O => \N__22095\,
            I => \N__22078\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__22092\,
            I => \N__22078\
        );

    \I__4364\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22075\
        );

    \I__4363\ : CascadeMux
    port map (
            O => \N__22088\,
            I => \N__22072\
        );

    \I__4362\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22067\
        );

    \I__4361\ : CascadeMux
    port map (
            O => \N__22084\,
            I => \N__22064\
        );

    \I__4360\ : CascadeMux
    port map (
            O => \N__22083\,
            I => \N__22061\
        );

    \I__4359\ : Span4Mux_v
    port map (
            O => \N__22078\,
            I => \N__22054\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__22075\,
            I => \N__22054\
        );

    \I__4357\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22051\
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__22071\,
            I => \N__22048\
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__22070\,
            I => \N__22043\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__22067\,
            I => \N__22038\
        );

    \I__4353\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22035\
        );

    \I__4352\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22032\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__22060\,
            I => \N__22029\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__22059\,
            I => \N__22026\
        );

    \I__4349\ : Span4Mux_h
    port map (
            O => \N__22054\,
            I => \N__22021\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__22051\,
            I => \N__22021\
        );

    \I__4347\ : InMux
    port map (
            O => \N__22048\,
            I => \N__22018\
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__22047\,
            I => \N__22015\
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__22046\,
            I => \N__22011\
        );

    \I__4344\ : InMux
    port map (
            O => \N__22043\,
            I => \N__22008\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__22042\,
            I => \N__22005\
        );

    \I__4342\ : CascadeMux
    port map (
            O => \N__22041\,
            I => \N__22002\
        );

    \I__4341\ : Span4Mux_s2_v
    port map (
            O => \N__22038\,
            I => \N__21997\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__22035\,
            I => \N__21997\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__22032\,
            I => \N__21994\
        );

    \I__4338\ : InMux
    port map (
            O => \N__22029\,
            I => \N__21991\
        );

    \I__4337\ : InMux
    port map (
            O => \N__22026\,
            I => \N__21988\
        );

    \I__4336\ : Span4Mux_v
    port map (
            O => \N__22021\,
            I => \N__21983\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__22018\,
            I => \N__21983\
        );

    \I__4334\ : InMux
    port map (
            O => \N__22015\,
            I => \N__21980\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__22014\,
            I => \N__21977\
        );

    \I__4332\ : InMux
    port map (
            O => \N__22011\,
            I => \N__21974\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__22008\,
            I => \N__21971\
        );

    \I__4330\ : InMux
    port map (
            O => \N__22005\,
            I => \N__21968\
        );

    \I__4329\ : InMux
    port map (
            O => \N__22002\,
            I => \N__21965\
        );

    \I__4328\ : Span4Mux_v
    port map (
            O => \N__21997\,
            I => \N__21956\
        );

    \I__4327\ : Span4Mux_v
    port map (
            O => \N__21994\,
            I => \N__21956\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__21991\,
            I => \N__21956\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__21988\,
            I => \N__21956\
        );

    \I__4324\ : Span4Mux_h
    port map (
            O => \N__21983\,
            I => \N__21951\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__21980\,
            I => \N__21951\
        );

    \I__4322\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21948\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__21974\,
            I => \N__21944\
        );

    \I__4320\ : Span4Mux_v
    port map (
            O => \N__21971\,
            I => \N__21937\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__21968\,
            I => \N__21937\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__21965\,
            I => \N__21937\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__21956\,
            I => \N__21928\
        );

    \I__4316\ : Span4Mux_v
    port map (
            O => \N__21951\,
            I => \N__21928\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__21948\,
            I => \N__21928\
        );

    \I__4314\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21925\
        );

    \I__4313\ : Span4Mux_v
    port map (
            O => \N__21944\,
            I => \N__21920\
        );

    \I__4312\ : Span4Mux_v
    port map (
            O => \N__21937\,
            I => \N__21920\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__21936\,
            I => \N__21916\
        );

    \I__4310\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21913\
        );

    \I__4309\ : Span4Mux_h
    port map (
            O => \N__21928\,
            I => \N__21908\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__21925\,
            I => \N__21908\
        );

    \I__4307\ : Sp12to4
    port map (
            O => \N__21920\,
            I => \N__21905\
        );

    \I__4306\ : InMux
    port map (
            O => \N__21919\,
            I => \N__21902\
        );

    \I__4305\ : InMux
    port map (
            O => \N__21916\,
            I => \N__21899\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__21913\,
            I => \N__21894\
        );

    \I__4303\ : Span4Mux_h
    port map (
            O => \N__21908\,
            I => \N__21894\
        );

    \I__4302\ : Odrv12
    port map (
            O => \N__21905\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__21902\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__21899\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__4299\ : Odrv4
    port map (
            O => \N__21894\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__4298\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21879\
        );

    \I__4297\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21879\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__21879\,
            I => \un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0\
        );

    \I__4295\ : InMux
    port map (
            O => \N__21876\,
            I => \un1_M_this_sprites_address_q_cry_4\
        );

    \I__4294\ : InMux
    port map (
            O => \N__21873\,
            I => \un1_M_this_sprites_address_q_cry_5\
        );

    \I__4293\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21867\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__21867\,
            I => \N__21864\
        );

    \I__4291\ : Odrv4
    port map (
            O => \N__21864\,
            I => \this_delay_clk.M_pipe_qZ0Z_3\
        );

    \I__4290\ : InMux
    port map (
            O => \N__21861\,
            I => \N__21858\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__21858\,
            I => \N__21855\
        );

    \I__4288\ : Span4Mux_h
    port map (
            O => \N__21855\,
            I => \N__21852\
        );

    \I__4287\ : Span4Mux_h
    port map (
            O => \N__21852\,
            I => \N__21849\
        );

    \I__4286\ : Odrv4
    port map (
            O => \N__21849\,
            I => \this_sprites_ram.mem_out_bus6_3\
        );

    \I__4285\ : InMux
    port map (
            O => \N__21846\,
            I => \N__21843\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__21843\,
            I => \N__21840\
        );

    \I__4283\ : Span4Mux_v
    port map (
            O => \N__21840\,
            I => \N__21837\
        );

    \I__4282\ : Sp12to4
    port map (
            O => \N__21837\,
            I => \N__21834\
        );

    \I__4281\ : Odrv12
    port map (
            O => \N__21834\,
            I => \this_sprites_ram.mem_out_bus2_3\
        );

    \I__4280\ : InMux
    port map (
            O => \N__21831\,
            I => \N__21828\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__21828\,
            I => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__21825\,
            I => \this_vga_signals.N_746_cascade_\
        );

    \I__4277\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21819\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__21819\,
            I => \this_vga_signals.N_505\
        );

    \I__4275\ : CascadeMux
    port map (
            O => \N__21816\,
            I => \N__21813\
        );

    \I__4274\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21810\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__21810\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_i_a4_2Z0Z_0\
        );

    \I__4272\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21804\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__21804\,
            I => \N__21801\
        );

    \I__4270\ : Span4Mux_h
    port map (
            O => \N__21801\,
            I => \N__21798\
        );

    \I__4269\ : Span4Mux_h
    port map (
            O => \N__21798\,
            I => \N__21795\
        );

    \I__4268\ : Sp12to4
    port map (
            O => \N__21795\,
            I => \N__21792\
        );

    \I__4267\ : Odrv12
    port map (
            O => \N__21792\,
            I => \this_sprites_ram.mem_out_bus4_1\
        );

    \I__4266\ : InMux
    port map (
            O => \N__21789\,
            I => \N__21786\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__21786\,
            I => \N__21783\
        );

    \I__4264\ : Span4Mux_h
    port map (
            O => \N__21783\,
            I => \N__21780\
        );

    \I__4263\ : Sp12to4
    port map (
            O => \N__21780\,
            I => \N__21777\
        );

    \I__4262\ : Span12Mux_v
    port map (
            O => \N__21777\,
            I => \N__21774\
        );

    \I__4261\ : Odrv12
    port map (
            O => \N__21774\,
            I => \this_sprites_ram.mem_out_bus0_1\
        );

    \I__4260\ : CascadeMux
    port map (
            O => \N__21771\,
            I => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0_cascade_\
        );

    \I__4259\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21758\
        );

    \I__4258\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21758\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__21766\,
            I => \N__21754\
        );

    \I__4256\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21750\
        );

    \I__4255\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21745\
        );

    \I__4254\ : InMux
    port map (
            O => \N__21763\,
            I => \N__21745\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21742\
        );

    \I__4252\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21739\
        );

    \I__4251\ : InMux
    port map (
            O => \N__21754\,
            I => \N__21734\
        );

    \I__4250\ : InMux
    port map (
            O => \N__21753\,
            I => \N__21734\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__21750\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__21745\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__21742\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__21739\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__21734\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__4244\ : CascadeMux
    port map (
            O => \N__21723\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\
        );

    \I__4243\ : InMux
    port map (
            O => \N__21720\,
            I => \N__21717\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__21717\,
            I => \N__21713\
        );

    \I__4241\ : InMux
    port map (
            O => \N__21716\,
            I => \N__21710\
        );

    \I__4240\ : Span12Mux_h
    port map (
            O => \N__21713\,
            I => \N__21707\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__21710\,
            I => \N__21704\
        );

    \I__4238\ : Odrv12
    port map (
            O => \N__21707\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__4237\ : Odrv4
    port map (
            O => \N__21704\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__4236\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21696\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__21696\,
            I => \N__21693\
        );

    \I__4234\ : Span12Mux_h
    port map (
            O => \N__21693\,
            I => \N__21690\
        );

    \I__4233\ : Span12Mux_v
    port map (
            O => \N__21690\,
            I => \N__21687\
        );

    \I__4232\ : Odrv12
    port map (
            O => \N__21687\,
            I => \M_this_oam_ram_read_data_6\
        );

    \I__4231\ : InMux
    port map (
            O => \N__21684\,
            I => \N__21681\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__21681\,
            I => \N__21678\
        );

    \I__4229\ : Sp12to4
    port map (
            O => \N__21678\,
            I => \N__21675\
        );

    \I__4228\ : Span12Mux_v
    port map (
            O => \N__21675\,
            I => \N__21672\
        );

    \I__4227\ : Span12Mux_h
    port map (
            O => \N__21672\,
            I => \N__21669\
        );

    \I__4226\ : Odrv12
    port map (
            O => \N__21669\,
            I => \M_this_map_ram_read_data_6\
        );

    \I__4225\ : CascadeMux
    port map (
            O => \N__21666\,
            I => \N__21663\
        );

    \I__4224\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21657\
        );

    \I__4223\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21654\
        );

    \I__4222\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21651\
        );

    \I__4221\ : InMux
    port map (
            O => \N__21660\,
            I => \N__21648\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__21657\,
            I => \N__21645\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__21654\,
            I => \N__21642\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__21651\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__21648\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__4216\ : Odrv4
    port map (
            O => \N__21645\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__4215\ : Odrv4
    port map (
            O => \N__21642\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__4214\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21630\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__21630\,
            I => \N__21627\
        );

    \I__4212\ : Span4Mux_h
    port map (
            O => \N__21627\,
            I => \N__21624\
        );

    \I__4211\ : Span4Mux_h
    port map (
            O => \N__21624\,
            I => \N__21621\
        );

    \I__4210\ : Odrv4
    port map (
            O => \N__21621\,
            I => \this_sprites_ram.mem_out_bus6_1\
        );

    \I__4209\ : InMux
    port map (
            O => \N__21618\,
            I => \N__21615\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__21615\,
            I => \N__21612\
        );

    \I__4207\ : Odrv12
    port map (
            O => \N__21612\,
            I => \this_sprites_ram.mem_out_bus2_1\
        );

    \I__4206\ : InMux
    port map (
            O => \N__21609\,
            I => \N__21606\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__21606\,
            I => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\
        );

    \I__4204\ : InMux
    port map (
            O => \N__21603\,
            I => \N__21600\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__21600\,
            I => \N__21597\
        );

    \I__4202\ : Span4Mux_h
    port map (
            O => \N__21597\,
            I => \N__21594\
        );

    \I__4201\ : Span4Mux_h
    port map (
            O => \N__21594\,
            I => \N__21591\
        );

    \I__4200\ : Span4Mux_v
    port map (
            O => \N__21591\,
            I => \N__21588\
        );

    \I__4199\ : Odrv4
    port map (
            O => \N__21588\,
            I => \this_sprites_ram.mem_out_bus5_1\
        );

    \I__4198\ : InMux
    port map (
            O => \N__21585\,
            I => \N__21582\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__21582\,
            I => \N__21579\
        );

    \I__4196\ : Span4Mux_h
    port map (
            O => \N__21579\,
            I => \N__21576\
        );

    \I__4195\ : Span4Mux_h
    port map (
            O => \N__21576\,
            I => \N__21573\
        );

    \I__4194\ : Span4Mux_v
    port map (
            O => \N__21573\,
            I => \N__21570\
        );

    \I__4193\ : Odrv4
    port map (
            O => \N__21570\,
            I => \this_sprites_ram.mem_out_bus1_1\
        );

    \I__4192\ : InMux
    port map (
            O => \N__21567\,
            I => \N__21564\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__21564\,
            I => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\
        );

    \I__4190\ : InMux
    port map (
            O => \N__21561\,
            I => \N__21558\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__21558\,
            I => \N__21555\
        );

    \I__4188\ : Odrv12
    port map (
            O => \N__21555\,
            I => \this_sprites_ram.mem_out_bus7_1\
        );

    \I__4187\ : InMux
    port map (
            O => \N__21552\,
            I => \N__21549\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__21549\,
            I => \N__21546\
        );

    \I__4185\ : Span4Mux_h
    port map (
            O => \N__21546\,
            I => \N__21543\
        );

    \I__4184\ : Span4Mux_h
    port map (
            O => \N__21543\,
            I => \N__21540\
        );

    \I__4183\ : Span4Mux_h
    port map (
            O => \N__21540\,
            I => \N__21537\
        );

    \I__4182\ : Odrv4
    port map (
            O => \N__21537\,
            I => \this_sprites_ram.mem_out_bus3_1\
        );

    \I__4181\ : InMux
    port map (
            O => \N__21534\,
            I => \N__21531\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__21531\,
            I => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\
        );

    \I__4179\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21525\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__21525\,
            I => \N__21520\
        );

    \I__4177\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21516\
        );

    \I__4176\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21513\
        );

    \I__4175\ : Span4Mux_h
    port map (
            O => \N__21520\,
            I => \N__21510\
        );

    \I__4174\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21507\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__21516\,
            I => \N__21504\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__21513\,
            I => \this_ppu.M_count_d_0_sqmuxa\
        );

    \I__4171\ : Odrv4
    port map (
            O => \N__21510\,
            I => \this_ppu.M_count_d_0_sqmuxa\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__21507\,
            I => \this_ppu.M_count_d_0_sqmuxa\
        );

    \I__4169\ : Odrv12
    port map (
            O => \N__21504\,
            I => \this_ppu.M_count_d_0_sqmuxa\
        );

    \I__4168\ : SRMux
    port map (
            O => \N__21495\,
            I => \N__21491\
        );

    \I__4167\ : SRMux
    port map (
            O => \N__21494\,
            I => \N__21488\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__21491\,
            I => \N__21485\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__21488\,
            I => \N__21481\
        );

    \I__4164\ : Span4Mux_v
    port map (
            O => \N__21485\,
            I => \N__21478\
        );

    \I__4163\ : SRMux
    port map (
            O => \N__21484\,
            I => \N__21475\
        );

    \I__4162\ : Span4Mux_h
    port map (
            O => \N__21481\,
            I => \N__21471\
        );

    \I__4161\ : Span4Mux_h
    port map (
            O => \N__21478\,
            I => \N__21466\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__21475\,
            I => \N__21466\
        );

    \I__4159\ : SRMux
    port map (
            O => \N__21474\,
            I => \N__21463\
        );

    \I__4158\ : Span4Mux_h
    port map (
            O => \N__21471\,
            I => \N__21460\
        );

    \I__4157\ : Span4Mux_h
    port map (
            O => \N__21466\,
            I => \N__21457\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__21463\,
            I => \N__21454\
        );

    \I__4155\ : Odrv4
    port map (
            O => \N__21460\,
            I => \this_ppu.M_last_q_RNIQRTEB\
        );

    \I__4154\ : Odrv4
    port map (
            O => \N__21457\,
            I => \this_ppu.M_last_q_RNIQRTEB\
        );

    \I__4153\ : Odrv12
    port map (
            O => \N__21454\,
            I => \this_ppu.M_last_q_RNIQRTEB\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__21447\,
            I => \N__21443\
        );

    \I__4151\ : CascadeMux
    port map (
            O => \N__21446\,
            I => \N__21440\
        );

    \I__4150\ : CascadeBuf
    port map (
            O => \N__21443\,
            I => \N__21437\
        );

    \I__4149\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21434\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__21437\,
            I => \N__21431\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__21434\,
            I => \N__21428\
        );

    \I__4146\ : InMux
    port map (
            O => \N__21431\,
            I => \N__21425\
        );

    \I__4145\ : Span4Mux_v
    port map (
            O => \N__21428\,
            I => \N__21421\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__21425\,
            I => \N__21418\
        );

    \I__4143\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21413\
        );

    \I__4142\ : Sp12to4
    port map (
            O => \N__21421\,
            I => \N__21410\
        );

    \I__4141\ : Span12Mux_h
    port map (
            O => \N__21418\,
            I => \N__21407\
        );

    \I__4140\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21404\
        );

    \I__4139\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21401\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__21413\,
            I => \N__21398\
        );

    \I__4137\ : Span12Mux_h
    port map (
            O => \N__21410\,
            I => \N__21393\
        );

    \I__4136\ : Span12Mux_v
    port map (
            O => \N__21407\,
            I => \N__21393\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__21404\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__21401\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4133\ : Odrv12
    port map (
            O => \N__21398\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4132\ : Odrv12
    port map (
            O => \N__21393\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4131\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21378\
        );

    \I__4130\ : InMux
    port map (
            O => \N__21383\,
            I => \N__21378\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__21378\,
            I => \this_ppu.un1_M_haddress_q_3_c2\
        );

    \I__4128\ : CascadeMux
    port map (
            O => \N__21375\,
            I => \N__21371\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__21374\,
            I => \N__21368\
        );

    \I__4126\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21365\
        );

    \I__4125\ : CascadeBuf
    port map (
            O => \N__21368\,
            I => \N__21362\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__21365\,
            I => \N__21358\
        );

    \I__4123\ : CascadeMux
    port map (
            O => \N__21362\,
            I => \N__21355\
        );

    \I__4122\ : InMux
    port map (
            O => \N__21361\,
            I => \N__21352\
        );

    \I__4121\ : Span4Mux_h
    port map (
            O => \N__21358\,
            I => \N__21349\
        );

    \I__4120\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21346\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__21352\,
            I => \N__21343\
        );

    \I__4118\ : Span4Mux_h
    port map (
            O => \N__21349\,
            I => \N__21340\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__21346\,
            I => \N__21337\
        );

    \I__4116\ : Span4Mux_v
    port map (
            O => \N__21343\,
            I => \N__21331\
        );

    \I__4115\ : Sp12to4
    port map (
            O => \N__21340\,
            I => \N__21326\
        );

    \I__4114\ : Span12Mux_h
    port map (
            O => \N__21337\,
            I => \N__21326\
        );

    \I__4113\ : InMux
    port map (
            O => \N__21336\,
            I => \N__21321\
        );

    \I__4112\ : InMux
    port map (
            O => \N__21335\,
            I => \N__21321\
        );

    \I__4111\ : InMux
    port map (
            O => \N__21334\,
            I => \N__21318\
        );

    \I__4110\ : Span4Mux_v
    port map (
            O => \N__21331\,
            I => \N__21315\
        );

    \I__4109\ : Span12Mux_v
    port map (
            O => \N__21326\,
            I => \N__21312\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__21321\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__21318\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__4106\ : Odrv4
    port map (
            O => \N__21315\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__4105\ : Odrv12
    port map (
            O => \N__21312\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__4104\ : CascadeMux
    port map (
            O => \N__21303\,
            I => \N__21300\
        );

    \I__4103\ : CascadeBuf
    port map (
            O => \N__21300\,
            I => \N__21297\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__21297\,
            I => \N__21294\
        );

    \I__4101\ : InMux
    port map (
            O => \N__21294\,
            I => \N__21291\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__21291\,
            I => \N__21287\
        );

    \I__4099\ : InMux
    port map (
            O => \N__21290\,
            I => \N__21284\
        );

    \I__4098\ : Span12Mux_h
    port map (
            O => \N__21287\,
            I => \N__21281\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__21284\,
            I => \N__21277\
        );

    \I__4096\ : Span12Mux_h
    port map (
            O => \N__21281\,
            I => \N__21274\
        );

    \I__4095\ : InMux
    port map (
            O => \N__21280\,
            I => \N__21271\
        );

    \I__4094\ : Span12Mux_h
    port map (
            O => \N__21277\,
            I => \N__21268\
        );

    \I__4093\ : Span12Mux_v
    port map (
            O => \N__21274\,
            I => \N__21265\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__21271\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__4091\ : Odrv12
    port map (
            O => \N__21268\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__4090\ : Odrv12
    port map (
            O => \N__21265\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__4089\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21249\
        );

    \I__4088\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21249\
        );

    \I__4087\ : InMux
    port map (
            O => \N__21256\,
            I => \N__21249\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__21249\,
            I => \this_ppu.un1_M_haddress_q_3_c5\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__21246\,
            I => \N__21242\
        );

    \I__4084\ : CascadeMux
    port map (
            O => \N__21245\,
            I => \N__21239\
        );

    \I__4083\ : CascadeBuf
    port map (
            O => \N__21242\,
            I => \N__21236\
        );

    \I__4082\ : InMux
    port map (
            O => \N__21239\,
            I => \N__21232\
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__21236\,
            I => \N__21229\
        );

    \I__4080\ : InMux
    port map (
            O => \N__21235\,
            I => \N__21226\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__21232\,
            I => \N__21223\
        );

    \I__4078\ : InMux
    port map (
            O => \N__21229\,
            I => \N__21220\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__21226\,
            I => \N__21215\
        );

    \I__4076\ : Span4Mux_h
    port map (
            O => \N__21223\,
            I => \N__21212\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__21220\,
            I => \N__21209\
        );

    \I__4074\ : CascadeMux
    port map (
            O => \N__21219\,
            I => \N__21206\
        );

    \I__4073\ : CascadeMux
    port map (
            O => \N__21218\,
            I => \N__21203\
        );

    \I__4072\ : Span4Mux_v
    port map (
            O => \N__21215\,
            I => \N__21199\
        );

    \I__4071\ : Sp12to4
    port map (
            O => \N__21212\,
            I => \N__21194\
        );

    \I__4070\ : Span12Mux_s11_h
    port map (
            O => \N__21209\,
            I => \N__21194\
        );

    \I__4069\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21187\
        );

    \I__4068\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21187\
        );

    \I__4067\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21187\
        );

    \I__4066\ : Span4Mux_v
    port map (
            O => \N__21199\,
            I => \N__21184\
        );

    \I__4065\ : Span12Mux_v
    port map (
            O => \N__21194\,
            I => \N__21181\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__21187\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__21184\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__4062\ : Odrv12
    port map (
            O => \N__21181\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__4061\ : CascadeMux
    port map (
            O => \N__21174\,
            I => \N__21171\
        );

    \I__4060\ : CascadeBuf
    port map (
            O => \N__21171\,
            I => \N__21167\
        );

    \I__4059\ : CascadeMux
    port map (
            O => \N__21170\,
            I => \N__21164\
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__21167\,
            I => \N__21161\
        );

    \I__4057\ : InMux
    port map (
            O => \N__21164\,
            I => \N__21157\
        );

    \I__4056\ : InMux
    port map (
            O => \N__21161\,
            I => \N__21154\
        );

    \I__4055\ : InMux
    port map (
            O => \N__21160\,
            I => \N__21151\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__21157\,
            I => \N__21148\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__21154\,
            I => \N__21145\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__21151\,
            I => \N__21142\
        );

    \I__4051\ : Span4Mux_v
    port map (
            O => \N__21148\,
            I => \N__21139\
        );

    \I__4050\ : Sp12to4
    port map (
            O => \N__21145\,
            I => \N__21136\
        );

    \I__4049\ : Span4Mux_v
    port map (
            O => \N__21142\,
            I => \N__21131\
        );

    \I__4048\ : Span4Mux_h
    port map (
            O => \N__21139\,
            I => \N__21128\
        );

    \I__4047\ : Span12Mux_h
    port map (
            O => \N__21136\,
            I => \N__21125\
        );

    \I__4046\ : InMux
    port map (
            O => \N__21135\,
            I => \N__21120\
        );

    \I__4045\ : InMux
    port map (
            O => \N__21134\,
            I => \N__21120\
        );

    \I__4044\ : Span4Mux_v
    port map (
            O => \N__21131\,
            I => \N__21117\
        );

    \I__4043\ : Span4Mux_h
    port map (
            O => \N__21128\,
            I => \N__21114\
        );

    \I__4042\ : Span12Mux_v
    port map (
            O => \N__21125\,
            I => \N__21111\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__21120\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__4040\ : Odrv4
    port map (
            O => \N__21117\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__4039\ : Odrv4
    port map (
            O => \N__21114\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__4038\ : Odrv12
    port map (
            O => \N__21111\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__4037\ : CEMux
    port map (
            O => \N__21102\,
            I => \N__21099\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__21099\,
            I => \N__21096\
        );

    \I__4035\ : Span4Mux_v
    port map (
            O => \N__21096\,
            I => \N__21093\
        );

    \I__4034\ : Span4Mux_h
    port map (
            O => \N__21093\,
            I => \N__21089\
        );

    \I__4033\ : InMux
    port map (
            O => \N__21092\,
            I => \N__21086\
        );

    \I__4032\ : Span4Mux_h
    port map (
            O => \N__21089\,
            I => \N__21082\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__21086\,
            I => \N__21079\
        );

    \I__4030\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21076\
        );

    \I__4029\ : Odrv4
    port map (
            O => \N__21082\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4028\ : Odrv4
    port map (
            O => \N__21079\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__21076\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4026\ : SRMux
    port map (
            O => \N__21069\,
            I => \N__21064\
        );

    \I__4025\ : SRMux
    port map (
            O => \N__21068\,
            I => \N__21061\
        );

    \I__4024\ : SRMux
    port map (
            O => \N__21067\,
            I => \N__21058\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__21064\,
            I => \N__21055\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__21061\,
            I => \N__21052\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__21058\,
            I => \N__21049\
        );

    \I__4020\ : Span4Mux_v
    port map (
            O => \N__21055\,
            I => \N__21046\
        );

    \I__4019\ : Span4Mux_v
    port map (
            O => \N__21052\,
            I => \N__21041\
        );

    \I__4018\ : Span4Mux_h
    port map (
            O => \N__21049\,
            I => \N__21041\
        );

    \I__4017\ : Odrv4
    port map (
            O => \N__21046\,
            I => \this_ppu.M_last_q_RNI3BB75\
        );

    \I__4016\ : Odrv4
    port map (
            O => \N__21041\,
            I => \this_ppu.M_last_q_RNI3BB75\
        );

    \I__4015\ : InMux
    port map (
            O => \N__21036\,
            I => \N__21033\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__21033\,
            I => \N__21030\
        );

    \I__4013\ : Span4Mux_v
    port map (
            O => \N__21030\,
            I => \N__21027\
        );

    \I__4012\ : Span4Mux_h
    port map (
            O => \N__21027\,
            I => \N__21024\
        );

    \I__4011\ : Sp12to4
    port map (
            O => \N__21024\,
            I => \N__21021\
        );

    \I__4010\ : Span12Mux_v
    port map (
            O => \N__21021\,
            I => \N__21018\
        );

    \I__4009\ : Odrv12
    port map (
            O => \N__21018\,
            I => \M_this_oam_ram_read_data_1\
        );

    \I__4008\ : InMux
    port map (
            O => \N__21015\,
            I => \N__21012\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__21012\,
            I => \N__21009\
        );

    \I__4006\ : Span4Mux_v
    port map (
            O => \N__21009\,
            I => \N__21006\
        );

    \I__4005\ : Sp12to4
    port map (
            O => \N__21006\,
            I => \N__21003\
        );

    \I__4004\ : Span12Mux_h
    port map (
            O => \N__21003\,
            I => \N__21000\
        );

    \I__4003\ : Odrv12
    port map (
            O => \N__21000\,
            I => \M_this_map_ram_read_data_1\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__20997\,
            I => \N__20989\
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__20996\,
            I => \N__20984\
        );

    \I__4000\ : CascadeMux
    port map (
            O => \N__20995\,
            I => \N__20981\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__20994\,
            I => \N__20977\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__20993\,
            I => \N__20973\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__20992\,
            I => \N__20969\
        );

    \I__3996\ : InMux
    port map (
            O => \N__20989\,
            I => \N__20966\
        );

    \I__3995\ : CascadeMux
    port map (
            O => \N__20988\,
            I => \N__20963\
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__20987\,
            I => \N__20958\
        );

    \I__3993\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20953\
        );

    \I__3992\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20950\
        );

    \I__3991\ : CascadeMux
    port map (
            O => \N__20980\,
            I => \N__20947\
        );

    \I__3990\ : InMux
    port map (
            O => \N__20977\,
            I => \N__20944\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__20976\,
            I => \N__20941\
        );

    \I__3988\ : InMux
    port map (
            O => \N__20973\,
            I => \N__20938\
        );

    \I__3987\ : CascadeMux
    port map (
            O => \N__20972\,
            I => \N__20935\
        );

    \I__3986\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20932\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__20966\,
            I => \N__20929\
        );

    \I__3984\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20926\
        );

    \I__3983\ : CascadeMux
    port map (
            O => \N__20962\,
            I => \N__20923\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__20961\,
            I => \N__20920\
        );

    \I__3981\ : InMux
    port map (
            O => \N__20958\,
            I => \N__20917\
        );

    \I__3980\ : CascadeMux
    port map (
            O => \N__20957\,
            I => \N__20913\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__20956\,
            I => \N__20910\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__20953\,
            I => \N__20907\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__20950\,
            I => \N__20904\
        );

    \I__3976\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20901\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__20944\,
            I => \N__20898\
        );

    \I__3974\ : InMux
    port map (
            O => \N__20941\,
            I => \N__20895\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__20938\,
            I => \N__20892\
        );

    \I__3972\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20889\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__20932\,
            I => \N__20886\
        );

    \I__3970\ : Span4Mux_h
    port map (
            O => \N__20929\,
            I => \N__20883\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__20926\,
            I => \N__20880\
        );

    \I__3968\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20877\
        );

    \I__3967\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20874\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__20917\,
            I => \N__20871\
        );

    \I__3965\ : CascadeMux
    port map (
            O => \N__20916\,
            I => \N__20868\
        );

    \I__3964\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20865\
        );

    \I__3963\ : InMux
    port map (
            O => \N__20910\,
            I => \N__20862\
        );

    \I__3962\ : Span4Mux_h
    port map (
            O => \N__20907\,
            I => \N__20859\
        );

    \I__3961\ : Span4Mux_h
    port map (
            O => \N__20904\,
            I => \N__20856\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__20901\,
            I => \N__20853\
        );

    \I__3959\ : Span4Mux_h
    port map (
            O => \N__20898\,
            I => \N__20850\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__20895\,
            I => \N__20847\
        );

    \I__3957\ : Span4Mux_h
    port map (
            O => \N__20892\,
            I => \N__20844\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__20889\,
            I => \N__20841\
        );

    \I__3955\ : Span4Mux_h
    port map (
            O => \N__20886\,
            I => \N__20836\
        );

    \I__3954\ : Span4Mux_v
    port map (
            O => \N__20883\,
            I => \N__20836\
        );

    \I__3953\ : Span4Mux_h
    port map (
            O => \N__20880\,
            I => \N__20833\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__20877\,
            I => \N__20830\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__20874\,
            I => \N__20827\
        );

    \I__3950\ : Span4Mux_h
    port map (
            O => \N__20871\,
            I => \N__20824\
        );

    \I__3949\ : InMux
    port map (
            O => \N__20868\,
            I => \N__20821\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__20865\,
            I => \N__20818\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__20862\,
            I => \N__20815\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__20859\,
            I => \N__20810\
        );

    \I__3945\ : Span4Mux_h
    port map (
            O => \N__20856\,
            I => \N__20810\
        );

    \I__3944\ : Span4Mux_h
    port map (
            O => \N__20853\,
            I => \N__20807\
        );

    \I__3943\ : Span4Mux_h
    port map (
            O => \N__20850\,
            I => \N__20804\
        );

    \I__3942\ : Span4Mux_h
    port map (
            O => \N__20847\,
            I => \N__20801\
        );

    \I__3941\ : Span4Mux_h
    port map (
            O => \N__20844\,
            I => \N__20798\
        );

    \I__3940\ : Span4Mux_h
    port map (
            O => \N__20841\,
            I => \N__20793\
        );

    \I__3939\ : Span4Mux_v
    port map (
            O => \N__20836\,
            I => \N__20793\
        );

    \I__3938\ : Span4Mux_h
    port map (
            O => \N__20833\,
            I => \N__20790\
        );

    \I__3937\ : Span4Mux_h
    port map (
            O => \N__20830\,
            I => \N__20787\
        );

    \I__3936\ : Span4Mux_h
    port map (
            O => \N__20827\,
            I => \N__20782\
        );

    \I__3935\ : Span4Mux_v
    port map (
            O => \N__20824\,
            I => \N__20782\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__20821\,
            I => \N__20775\
        );

    \I__3933\ : Span4Mux_v
    port map (
            O => \N__20818\,
            I => \N__20775\
        );

    \I__3932\ : Span4Mux_v
    port map (
            O => \N__20815\,
            I => \N__20775\
        );

    \I__3931\ : Span4Mux_h
    port map (
            O => \N__20810\,
            I => \N__20768\
        );

    \I__3930\ : Span4Mux_h
    port map (
            O => \N__20807\,
            I => \N__20768\
        );

    \I__3929\ : Span4Mux_h
    port map (
            O => \N__20804\,
            I => \N__20768\
        );

    \I__3928\ : Span4Mux_h
    port map (
            O => \N__20801\,
            I => \N__20759\
        );

    \I__3927\ : Span4Mux_h
    port map (
            O => \N__20798\,
            I => \N__20759\
        );

    \I__3926\ : Span4Mux_h
    port map (
            O => \N__20793\,
            I => \N__20759\
        );

    \I__3925\ : Span4Mux_h
    port map (
            O => \N__20790\,
            I => \N__20759\
        );

    \I__3924\ : Span4Mux_h
    port map (
            O => \N__20787\,
            I => \N__20754\
        );

    \I__3923\ : Span4Mux_h
    port map (
            O => \N__20782\,
            I => \N__20754\
        );

    \I__3922\ : Sp12to4
    port map (
            O => \N__20775\,
            I => \N__20751\
        );

    \I__3921\ : Sp12to4
    port map (
            O => \N__20768\,
            I => \N__20742\
        );

    \I__3920\ : Sp12to4
    port map (
            O => \N__20759\,
            I => \N__20742\
        );

    \I__3919\ : Sp12to4
    port map (
            O => \N__20754\,
            I => \N__20742\
        );

    \I__3918\ : Span12Mux_h
    port map (
            O => \N__20751\,
            I => \N__20742\
        );

    \I__3917\ : Odrv12
    port map (
            O => \N__20742\,
            I => \M_this_ppu_sprites_addr_7\
        );

    \I__3916\ : CascadeMux
    port map (
            O => \N__20739\,
            I => \N__20736\
        );

    \I__3915\ : InMux
    port map (
            O => \N__20736\,
            I => \N__20732\
        );

    \I__3914\ : CascadeMux
    port map (
            O => \N__20735\,
            I => \N__20729\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__20732\,
            I => \N__20726\
        );

    \I__3912\ : InMux
    port map (
            O => \N__20729\,
            I => \N__20723\
        );

    \I__3911\ : Odrv4
    port map (
            O => \N__20726\,
            I => \this_ppu.M_this_ppu_map_addr_i_3\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__20723\,
            I => \this_ppu.M_this_ppu_map_addr_i_3\
        );

    \I__3909\ : CascadeMux
    port map (
            O => \N__20718\,
            I => \N__20715\
        );

    \I__3908\ : InMux
    port map (
            O => \N__20715\,
            I => \N__20711\
        );

    \I__3907\ : CascadeMux
    port map (
            O => \N__20714\,
            I => \N__20708\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__20711\,
            I => \N__20705\
        );

    \I__3905\ : InMux
    port map (
            O => \N__20708\,
            I => \N__20702\
        );

    \I__3904\ : Odrv4
    port map (
            O => \N__20705\,
            I => \this_ppu.M_this_ppu_map_addr_i_4\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__20702\,
            I => \this_ppu.M_this_ppu_map_addr_i_4\
        );

    \I__3902\ : InMux
    port map (
            O => \N__20697\,
            I => \bfn_19_8_0_\
        );

    \I__3901\ : InMux
    port map (
            O => \N__20694\,
            I => \N__20691\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__20691\,
            I => \N__20688\
        );

    \I__3899\ : Span4Mux_h
    port map (
            O => \N__20688\,
            I => \N__20683\
        );

    \I__3898\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20680\
        );

    \I__3897\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20677\
        );

    \I__3896\ : Odrv4
    port map (
            O => \N__20683\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__20680\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__20677\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__3893\ : InMux
    port map (
            O => \N__20670\,
            I => \N__20666\
        );

    \I__3892\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20662\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__20666\,
            I => \N__20659\
        );

    \I__3890\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20656\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__20662\,
            I => \N__20651\
        );

    \I__3888\ : Span4Mux_v
    port map (
            O => \N__20659\,
            I => \N__20651\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__20656\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__3886\ : Odrv4
    port map (
            O => \N__20651\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__3885\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20643\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__20643\,
            I => \N__20639\
        );

    \I__3883\ : CascadeMux
    port map (
            O => \N__20642\,
            I => \N__20636\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__20639\,
            I => \N__20633\
        );

    \I__3881\ : InMux
    port map (
            O => \N__20636\,
            I => \N__20630\
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__20633\,
            I => \this_ppu.N_122\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__20630\,
            I => \this_ppu.N_122\
        );

    \I__3878\ : InMux
    port map (
            O => \N__20625\,
            I => \N__20622\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__20622\,
            I => \N__20617\
        );

    \I__3876\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20612\
        );

    \I__3875\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20612\
        );

    \I__3874\ : Span4Mux_v
    port map (
            O => \N__20617\,
            I => \N__20607\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__20612\,
            I => \N__20607\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__20607\,
            I => \this_ppu.un1_M_vaddress_q_2_c2\
        );

    \I__3871\ : InMux
    port map (
            O => \N__20604\,
            I => \N__20600\
        );

    \I__3870\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20597\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__20600\,
            I => \N__20594\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__20597\,
            I => \N__20590\
        );

    \I__3867\ : Span4Mux_h
    port map (
            O => \N__20594\,
            I => \N__20586\
        );

    \I__3866\ : InMux
    port map (
            O => \N__20593\,
            I => \N__20582\
        );

    \I__3865\ : Span4Mux_v
    port map (
            O => \N__20590\,
            I => \N__20579\
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__20589\,
            I => \N__20576\
        );

    \I__3863\ : Sp12to4
    port map (
            O => \N__20586\,
            I => \N__20573\
        );

    \I__3862\ : InMux
    port map (
            O => \N__20585\,
            I => \N__20570\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__20582\,
            I => \N__20567\
        );

    \I__3860\ : Sp12to4
    port map (
            O => \N__20579\,
            I => \N__20564\
        );

    \I__3859\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20561\
        );

    \I__3858\ : Span12Mux_v
    port map (
            O => \N__20573\,
            I => \N__20558\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__20570\,
            I => \N__20555\
        );

    \I__3856\ : Span4Mux_v
    port map (
            O => \N__20567\,
            I => \N__20552\
        );

    \I__3855\ : Span12Mux_s11_h
    port map (
            O => \N__20564\,
            I => \N__20547\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__20561\,
            I => \N__20547\
        );

    \I__3853\ : Odrv12
    port map (
            O => \N__20558\,
            I => this_vga_signals_vvisibility
        );

    \I__3852\ : Odrv12
    port map (
            O => \N__20555\,
            I => this_vga_signals_vvisibility
        );

    \I__3851\ : Odrv4
    port map (
            O => \N__20552\,
            I => this_vga_signals_vvisibility
        );

    \I__3850\ : Odrv12
    port map (
            O => \N__20547\,
            I => this_vga_signals_vvisibility
        );

    \I__3849\ : InMux
    port map (
            O => \N__20538\,
            I => \bfn_19_6_0_\
        );

    \I__3848\ : CascadeMux
    port map (
            O => \N__20535\,
            I => \N__20532\
        );

    \I__3847\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20528\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__20531\,
            I => \N__20525\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__20528\,
            I => \N__20522\
        );

    \I__3844\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20519\
        );

    \I__3843\ : Odrv4
    port map (
            O => \N__20522\,
            I => \this_ppu.M_this_ppu_vram_addr_i_0\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__20519\,
            I => \this_ppu.M_this_ppu_vram_addr_i_0\
        );

    \I__3841\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20510\
        );

    \I__3840\ : CascadeMux
    port map (
            O => \N__20513\,
            I => \N__20507\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__20510\,
            I => \N__20504\
        );

    \I__3838\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20501\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__20504\,
            I => \this_ppu.M_this_ppu_vram_addr_i_1\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__20501\,
            I => \this_ppu.M_this_ppu_vram_addr_i_1\
        );

    \I__3835\ : InMux
    port map (
            O => \N__20496\,
            I => \N__20493\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__20493\,
            I => \N__20489\
        );

    \I__3833\ : InMux
    port map (
            O => \N__20492\,
            I => \N__20486\
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__20489\,
            I => \this_ppu.M_this_ppu_vram_addr_i_2\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__20486\,
            I => \this_ppu.M_this_ppu_vram_addr_i_2\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__20481\,
            I => \N__20478\
        );

    \I__3829\ : InMux
    port map (
            O => \N__20478\,
            I => \N__20474\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__20477\,
            I => \N__20471\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__20474\,
            I => \N__20468\
        );

    \I__3826\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20465\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__20468\,
            I => \this_ppu.M_this_ppu_map_addr_i_0\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__20465\,
            I => \this_ppu.M_this_ppu_map_addr_i_0\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__20460\,
            I => \N__20457\
        );

    \I__3822\ : InMux
    port map (
            O => \N__20457\,
            I => \N__20454\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__20454\,
            I => \N__20450\
        );

    \I__3820\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20447\
        );

    \I__3819\ : Odrv4
    port map (
            O => \N__20450\,
            I => \this_ppu.M_this_ppu_map_addr_i_1\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__20447\,
            I => \this_ppu.M_this_ppu_map_addr_i_1\
        );

    \I__3817\ : CascadeMux
    port map (
            O => \N__20442\,
            I => \N__20439\
        );

    \I__3816\ : InMux
    port map (
            O => \N__20439\,
            I => \N__20435\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__20438\,
            I => \N__20432\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__20435\,
            I => \N__20429\
        );

    \I__3813\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20426\
        );

    \I__3812\ : Odrv4
    port map (
            O => \N__20429\,
            I => \this_ppu.M_this_ppu_map_addr_i_2\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__20426\,
            I => \this_ppu.M_this_ppu_map_addr_i_2\
        );

    \I__3810\ : InMux
    port map (
            O => \N__20421\,
            I => \N__20418\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__20418\,
            I => \N_617\
        );

    \I__3808\ : InMux
    port map (
            O => \N__20415\,
            I => \N__20412\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__20412\,
            I => \M_this_sprites_address_qc_11_0\
        );

    \I__3806\ : InMux
    port map (
            O => \N__20409\,
            I => \N__20406\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__20406\,
            I => \N_896_0\
        );

    \I__3804\ : InMux
    port map (
            O => \N__20403\,
            I => \N__20400\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__20400\,
            I => \N_512_0\
        );

    \I__3802\ : CascadeMux
    port map (
            O => \N__20397\,
            I => \N__20394\
        );

    \I__3801\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20391\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__20391\,
            I => \N__20388\
        );

    \I__3799\ : Odrv4
    port map (
            O => \N__20388\,
            I => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_8\
        );

    \I__3798\ : InMux
    port map (
            O => \N__20385\,
            I => \N__20382\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__20382\,
            I => \N__20379\
        );

    \I__3796\ : Span4Mux_v
    port map (
            O => \N__20379\,
            I => \N__20376\
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__20376\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1Z0Z_5\
        );

    \I__3794\ : CascadeMux
    port map (
            O => \N__20373\,
            I => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_11_cascade_\
        );

    \I__3793\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20367\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__20367\,
            I => \N__20364\
        );

    \I__3791\ : Odrv4
    port map (
            O => \N__20364\,
            I => \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_1\
        );

    \I__3790\ : InMux
    port map (
            O => \N__20361\,
            I => \N__20358\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__20358\,
            I => \M_this_sprites_address_qc_10_0\
        );

    \I__3788\ : CascadeMux
    port map (
            O => \N__20355\,
            I => \N_1286_tz_0_cascade_\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__20352\,
            I => \N_562_cascade_\
        );

    \I__3786\ : InMux
    port map (
            O => \N__20349\,
            I => \N__20346\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__20346\,
            I => \M_this_sprites_address_q_0_0_i_476\
        );

    \I__3784\ : CascadeMux
    port map (
            O => \N__20343\,
            I => \M_this_sprites_address_q_0_0_i_496_cascade_\
        );

    \I__3783\ : InMux
    port map (
            O => \N__20340\,
            I => \N__20337\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__20337\,
            I => \M_this_sprites_address_qc_0_1\
        );

    \I__3781\ : CascadeMux
    port map (
            O => \N__20334\,
            I => \N__20331\
        );

    \I__3780\ : InMux
    port map (
            O => \N__20331\,
            I => \N__20328\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__20328\,
            I => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_0\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__20325\,
            I => \N_773_cascade_\
        );

    \I__3777\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20319\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__20319\,
            I => \M_this_sprites_address_q_0_0_i_492\
        );

    \I__3775\ : CascadeMux
    port map (
            O => \N__20316\,
            I => \M_this_sprites_address_qc_1_0_cascade_\
        );

    \I__3774\ : CascadeMux
    port map (
            O => \N__20313\,
            I => \this_vga_signals.N_419_0_cascade_\
        );

    \I__3773\ : CascadeMux
    port map (
            O => \N__20310\,
            I => \N_440_0_cascade_\
        );

    \I__3772\ : CascadeMux
    port map (
            O => \N__20307\,
            I => \this_vga_signals.N_467_0_cascade_\
        );

    \I__3771\ : InMux
    port map (
            O => \N__20304\,
            I => \N__20301\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__20301\,
            I => \this_vga_signals.N_467_0\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__20298\,
            I => \N__20295\
        );

    \I__3768\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20292\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__20292\,
            I => \N__20289\
        );

    \I__3766\ : Span4Mux_v
    port map (
            O => \N__20289\,
            I => \N__20286\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__20286\,
            I => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0Z0Z_6\
        );

    \I__3764\ : InMux
    port map (
            O => \N__20283\,
            I => \N__20280\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__20280\,
            I => \N_510_0\
        );

    \I__3762\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20274\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__20274\,
            I => \N__20271\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__20271\,
            I => \M_this_sprites_address_qc_5_0\
        );

    \I__3759\ : InMux
    port map (
            O => \N__20268\,
            I => \N__20265\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__20265\,
            I => \N__20262\
        );

    \I__3757\ : Span4Mux_v
    port map (
            O => \N__20262\,
            I => \N__20259\
        );

    \I__3756\ : Span4Mux_h
    port map (
            O => \N__20259\,
            I => \N__20256\
        );

    \I__3755\ : Span4Mux_h
    port map (
            O => \N__20256\,
            I => \N__20253\
        );

    \I__3754\ : Odrv4
    port map (
            O => \N__20253\,
            I => \this_sprites_ram.mem_out_bus5_2\
        );

    \I__3753\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20247\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__20247\,
            I => \N__20244\
        );

    \I__3751\ : Span4Mux_h
    port map (
            O => \N__20244\,
            I => \N__20241\
        );

    \I__3750\ : Span4Mux_h
    port map (
            O => \N__20241\,
            I => \N__20238\
        );

    \I__3749\ : Odrv4
    port map (
            O => \N__20238\,
            I => \this_sprites_ram.mem_out_bus1_2\
        );

    \I__3748\ : InMux
    port map (
            O => \N__20235\,
            I => \N__20232\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__20232\,
            I => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\
        );

    \I__3746\ : IoInMux
    port map (
            O => \N__20229\,
            I => \N__20225\
        );

    \I__3745\ : IoInMux
    port map (
            O => \N__20228\,
            I => \N__20222\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__20225\,
            I => \N__20216\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__20222\,
            I => \N__20216\
        );

    \I__3742\ : IoInMux
    port map (
            O => \N__20221\,
            I => \N__20208\
        );

    \I__3741\ : IoSpan4Mux
    port map (
            O => \N__20216\,
            I => \N__20205\
        );

    \I__3740\ : IoInMux
    port map (
            O => \N__20215\,
            I => \N__20202\
        );

    \I__3739\ : IoInMux
    port map (
            O => \N__20214\,
            I => \N__20199\
        );

    \I__3738\ : IoInMux
    port map (
            O => \N__20213\,
            I => \N__20196\
        );

    \I__3737\ : IoInMux
    port map (
            O => \N__20212\,
            I => \N__20193\
        );

    \I__3736\ : IoInMux
    port map (
            O => \N__20211\,
            I => \N__20189\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__20208\,
            I => \N__20184\
        );

    \I__3734\ : IoSpan4Mux
    port map (
            O => \N__20205\,
            I => \N__20181\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__20202\,
            I => \N__20172\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__20199\,
            I => \N__20172\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__20196\,
            I => \N__20172\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__20193\,
            I => \N__20172\
        );

    \I__3729\ : IoInMux
    port map (
            O => \N__20192\,
            I => \N__20169\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__20189\,
            I => \N__20166\
        );

    \I__3727\ : IoInMux
    port map (
            O => \N__20188\,
            I => \N__20163\
        );

    \I__3726\ : IoInMux
    port map (
            O => \N__20187\,
            I => \N__20160\
        );

    \I__3725\ : Span4Mux_s1_h
    port map (
            O => \N__20184\,
            I => \N__20152\
        );

    \I__3724\ : IoSpan4Mux
    port map (
            O => \N__20181\,
            I => \N__20144\
        );

    \I__3723\ : IoSpan4Mux
    port map (
            O => \N__20172\,
            I => \N__20144\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__20169\,
            I => \N__20144\
        );

    \I__3721\ : IoSpan4Mux
    port map (
            O => \N__20166\,
            I => \N__20139\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__20163\,
            I => \N__20139\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__20160\,
            I => \N__20136\
        );

    \I__3718\ : IoInMux
    port map (
            O => \N__20159\,
            I => \N__20133\
        );

    \I__3717\ : IoInMux
    port map (
            O => \N__20158\,
            I => \N__20130\
        );

    \I__3716\ : IoInMux
    port map (
            O => \N__20157\,
            I => \N__20127\
        );

    \I__3715\ : IoInMux
    port map (
            O => \N__20156\,
            I => \N__20124\
        );

    \I__3714\ : IoInMux
    port map (
            O => \N__20155\,
            I => \N__20121\
        );

    \I__3713\ : Span4Mux_h
    port map (
            O => \N__20152\,
            I => \N__20118\
        );

    \I__3712\ : IoInMux
    port map (
            O => \N__20151\,
            I => \N__20115\
        );

    \I__3711\ : IoSpan4Mux
    port map (
            O => \N__20144\,
            I => \N__20112\
        );

    \I__3710\ : IoSpan4Mux
    port map (
            O => \N__20139\,
            I => \N__20105\
        );

    \I__3709\ : IoSpan4Mux
    port map (
            O => \N__20136\,
            I => \N__20105\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__20133\,
            I => \N__20105\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__20130\,
            I => \N__20100\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__20127\,
            I => \N__20100\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__20124\,
            I => \N__20097\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__20121\,
            I => \N__20094\
        );

    \I__3703\ : Sp12to4
    port map (
            O => \N__20118\,
            I => \N__20091\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__20115\,
            I => \N__20088\
        );

    \I__3701\ : Span4Mux_s0_h
    port map (
            O => \N__20112\,
            I => \N__20085\
        );

    \I__3700\ : IoSpan4Mux
    port map (
            O => \N__20105\,
            I => \N__20080\
        );

    \I__3699\ : IoSpan4Mux
    port map (
            O => \N__20100\,
            I => \N__20080\
        );

    \I__3698\ : Span12Mux_s4_v
    port map (
            O => \N__20097\,
            I => \N__20075\
        );

    \I__3697\ : Span12Mux_s2_h
    port map (
            O => \N__20094\,
            I => \N__20075\
        );

    \I__3696\ : Span12Mux_v
    port map (
            O => \N__20091\,
            I => \N__20072\
        );

    \I__3695\ : Span12Mux_s2_h
    port map (
            O => \N__20088\,
            I => \N__20067\
        );

    \I__3694\ : Sp12to4
    port map (
            O => \N__20085\,
            I => \N__20067\
        );

    \I__3693\ : Span4Mux_s3_v
    port map (
            O => \N__20080\,
            I => \N__20064\
        );

    \I__3692\ : Span12Mux_h
    port map (
            O => \N__20075\,
            I => \N__20055\
        );

    \I__3691\ : Span12Mux_h
    port map (
            O => \N__20072\,
            I => \N__20055\
        );

    \I__3690\ : Span12Mux_h
    port map (
            O => \N__20067\,
            I => \N__20055\
        );

    \I__3689\ : Sp12to4
    port map (
            O => \N__20064\,
            I => \N__20055\
        );

    \I__3688\ : Odrv12
    port map (
            O => \N__20055\,
            I => dma_0_i
        );

    \I__3687\ : InMux
    port map (
            O => \N__20052\,
            I => \N__20049\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__20049\,
            I => \N__20046\
        );

    \I__3685\ : Span12Mux_h
    port map (
            O => \N__20046\,
            I => \N__20043\
        );

    \I__3684\ : Span12Mux_v
    port map (
            O => \N__20043\,
            I => \N__20040\
        );

    \I__3683\ : Odrv12
    port map (
            O => \N__20040\,
            I => \this_sprites_ram.mem_out_bus4_3\
        );

    \I__3682\ : InMux
    port map (
            O => \N__20037\,
            I => \N__20034\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__20034\,
            I => \N__20031\
        );

    \I__3680\ : Span4Mux_v
    port map (
            O => \N__20031\,
            I => \N__20028\
        );

    \I__3679\ : Span4Mux_h
    port map (
            O => \N__20028\,
            I => \N__20025\
        );

    \I__3678\ : Span4Mux_v
    port map (
            O => \N__20025\,
            I => \N__20022\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__20022\,
            I => \this_sprites_ram.mem_out_bus0_3\
        );

    \I__3676\ : CascadeMux
    port map (
            O => \N__20019\,
            I => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0_cascade_\
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__20016\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\
        );

    \I__3674\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20010\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__20010\,
            I => \N__20007\
        );

    \I__3672\ : Span4Mux_h
    port map (
            O => \N__20007\,
            I => \N__20003\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__20006\,
            I => \N__20000\
        );

    \I__3670\ : Span4Mux_h
    port map (
            O => \N__20003\,
            I => \N__19997\
        );

    \I__3669\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19994\
        );

    \I__3668\ : Span4Mux_h
    port map (
            O => \N__19997\,
            I => \N__19991\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__19994\,
            I => \N__19988\
        );

    \I__3666\ : Odrv4
    port map (
            O => \N__19991\,
            I => \M_this_ppu_vram_data_3\
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__19988\,
            I => \M_this_ppu_vram_data_3\
        );

    \I__3664\ : InMux
    port map (
            O => \N__19983\,
            I => \N__19980\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__19980\,
            I => \N__19977\
        );

    \I__3662\ : Span4Mux_h
    port map (
            O => \N__19977\,
            I => \N__19974\
        );

    \I__3661\ : Span4Mux_v
    port map (
            O => \N__19974\,
            I => \N__19971\
        );

    \I__3660\ : Span4Mux_h
    port map (
            O => \N__19971\,
            I => \N__19968\
        );

    \I__3659\ : Odrv4
    port map (
            O => \N__19968\,
            I => \this_sprites_ram.mem_out_bus5_3\
        );

    \I__3658\ : InMux
    port map (
            O => \N__19965\,
            I => \N__19962\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__19962\,
            I => \N__19959\
        );

    \I__3656\ : Span4Mux_v
    port map (
            O => \N__19959\,
            I => \N__19956\
        );

    \I__3655\ : Span4Mux_h
    port map (
            O => \N__19956\,
            I => \N__19953\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__19953\,
            I => \this_sprites_ram.mem_out_bus1_3\
        );

    \I__3653\ : InMux
    port map (
            O => \N__19950\,
            I => \N__19947\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__19947\,
            I => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\
        );

    \I__3651\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19941\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__19941\,
            I => \N__19938\
        );

    \I__3649\ : Span4Mux_h
    port map (
            O => \N__19938\,
            I => \N__19935\
        );

    \I__3648\ : Span4Mux_h
    port map (
            O => \N__19935\,
            I => \N__19932\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__19932\,
            I => \this_sprites_ram.mem_out_bus7_3\
        );

    \I__3646\ : InMux
    port map (
            O => \N__19929\,
            I => \N__19926\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__19926\,
            I => \N__19923\
        );

    \I__3644\ : Span4Mux_v
    port map (
            O => \N__19923\,
            I => \N__19920\
        );

    \I__3643\ : Span4Mux_v
    port map (
            O => \N__19920\,
            I => \N__19917\
        );

    \I__3642\ : Sp12to4
    port map (
            O => \N__19917\,
            I => \N__19914\
        );

    \I__3641\ : Odrv12
    port map (
            O => \N__19914\,
            I => \this_sprites_ram.mem_out_bus3_3\
        );

    \I__3640\ : InMux
    port map (
            O => \N__19911\,
            I => \N__19908\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__19908\,
            I => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\
        );

    \I__3638\ : InMux
    port map (
            O => \N__19905\,
            I => \N__19901\
        );

    \I__3637\ : InMux
    port map (
            O => \N__19904\,
            I => \N__19898\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__19901\,
            I => \N__19891\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__19898\,
            I => \N__19891\
        );

    \I__3634\ : InMux
    port map (
            O => \N__19897\,
            I => \N__19886\
        );

    \I__3633\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19886\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__19891\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__19886\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__3630\ : InMux
    port map (
            O => \N__19881\,
            I => \N__19878\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__19878\,
            I => \N__19875\
        );

    \I__3628\ : Span4Mux_v
    port map (
            O => \N__19875\,
            I => \N__19872\
        );

    \I__3627\ : Sp12to4
    port map (
            O => \N__19872\,
            I => \N__19869\
        );

    \I__3626\ : Span12Mux_h
    port map (
            O => \N__19869\,
            I => \N__19866\
        );

    \I__3625\ : Span12Mux_v
    port map (
            O => \N__19866\,
            I => \N__19863\
        );

    \I__3624\ : Odrv12
    port map (
            O => \N__19863\,
            I => \this_sprites_ram.mem_out_bus4_0\
        );

    \I__3623\ : InMux
    port map (
            O => \N__19860\,
            I => \N__19857\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__19857\,
            I => \N__19854\
        );

    \I__3621\ : Span4Mux_h
    port map (
            O => \N__19854\,
            I => \N__19851\
        );

    \I__3620\ : Span4Mux_h
    port map (
            O => \N__19851\,
            I => \N__19848\
        );

    \I__3619\ : Span4Mux_v
    port map (
            O => \N__19848\,
            I => \N__19845\
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__19845\,
            I => \this_sprites_ram.mem_out_bus0_0\
        );

    \I__3617\ : InMux
    port map (
            O => \N__19842\,
            I => \N__19838\
        );

    \I__3616\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19835\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__19838\,
            I => \N__19832\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__19835\,
            I => \N__19829\
        );

    \I__3613\ : Odrv12
    port map (
            O => \N__19832\,
            I => \this_ppu.vram_en_i_a2Z0Z_0\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__19829\,
            I => \this_ppu.vram_en_i_a2Z0Z_0\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__19824\,
            I => \this_ppu.vram_en_i_a2Z0Z_0_cascade_\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__19821\,
            I => \M_this_ppu_vram_en_0_cascade_\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__19818\,
            I => \this_ppu.un1_M_haddress_q_3_c2_cascade_\
        );

    \I__3608\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19812\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__19812\,
            I => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\
        );

    \I__3606\ : InMux
    port map (
            O => \N__19809\,
            I => \N__19806\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__19806\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2\
        );

    \I__3604\ : InMux
    port map (
            O => \N__19803\,
            I => \N__19800\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__19800\,
            I => \N__19797\
        );

    \I__3602\ : Span12Mux_h
    port map (
            O => \N__19797\,
            I => \N__19793\
        );

    \I__3601\ : InMux
    port map (
            O => \N__19796\,
            I => \N__19790\
        );

    \I__3600\ : Odrv12
    port map (
            O => \N__19793\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__19790\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__3598\ : InMux
    port map (
            O => \N__19785\,
            I => \N__19782\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__19782\,
            I => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0\
        );

    \I__3596\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19776\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__19776\,
            I => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\
        );

    \I__3594\ : InMux
    port map (
            O => \N__19773\,
            I => \N__19770\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__19770\,
            I => \N__19767\
        );

    \I__3592\ : Span4Mux_h
    port map (
            O => \N__19767\,
            I => \N__19764\
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__19764\,
            I => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__19761\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0_cascade_\
        );

    \I__3589\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__19755\,
            I => \N__19752\
        );

    \I__3587\ : Span12Mux_h
    port map (
            O => \N__19752\,
            I => \N__19748\
        );

    \I__3586\ : InMux
    port map (
            O => \N__19751\,
            I => \N__19745\
        );

    \I__3585\ : Odrv12
    port map (
            O => \N__19748\,
            I => \M_this_ppu_vram_data_0\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__19745\,
            I => \M_this_ppu_vram_data_0\
        );

    \I__3583\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19737\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__19737\,
            I => \this_ppu.N_124\
        );

    \I__3581\ : CascadeMux
    port map (
            O => \N__19734\,
            I => \this_ppu.N_124_cascade_\
        );

    \I__3580\ : CascadeMux
    port map (
            O => \N__19731\,
            I => \this_ppu.un1_M_vaddress_q_2_c5_cascade_\
        );

    \I__3579\ : InMux
    port map (
            O => \N__19728\,
            I => \N__19724\
        );

    \I__3578\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19721\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__19724\,
            I => \this_ppu.un1_M_vaddress_q_2_c5\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__19721\,
            I => \this_ppu.un1_M_vaddress_q_2_c5\
        );

    \I__3575\ : InMux
    port map (
            O => \N__19716\,
            I => \N__19712\
        );

    \I__3574\ : InMux
    port map (
            O => \N__19715\,
            I => \N__19706\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__19712\,
            I => \N__19703\
        );

    \I__3572\ : InMux
    port map (
            O => \N__19711\,
            I => \N__19696\
        );

    \I__3571\ : InMux
    port map (
            O => \N__19710\,
            I => \N__19696\
        );

    \I__3570\ : InMux
    port map (
            O => \N__19709\,
            I => \N__19696\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__19706\,
            I => \this_ppu.M_last_q\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__19703\,
            I => \this_ppu.M_last_q\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__19696\,
            I => \this_ppu.M_last_q\
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__19689\,
            I => \N__19685\
        );

    \I__3565\ : CascadeMux
    port map (
            O => \N__19688\,
            I => \N__19680\
        );

    \I__3564\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19677\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__19684\,
            I => \N__19674\
        );

    \I__3562\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19665\
        );

    \I__3561\ : InMux
    port map (
            O => \N__19680\,
            I => \N__19665\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__19677\,
            I => \N__19662\
        );

    \I__3559\ : InMux
    port map (
            O => \N__19674\,
            I => \N__19655\
        );

    \I__3558\ : InMux
    port map (
            O => \N__19673\,
            I => \N__19655\
        );

    \I__3557\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19655\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__19671\,
            I => \N__19652\
        );

    \I__3555\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19649\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__19665\,
            I => \N__19642\
        );

    \I__3553\ : Span4Mux_h
    port map (
            O => \N__19662\,
            I => \N__19642\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__19655\,
            I => \N__19642\
        );

    \I__3551\ : InMux
    port map (
            O => \N__19652\,
            I => \N__19639\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__19649\,
            I => \N__19636\
        );

    \I__3549\ : Span4Mux_h
    port map (
            O => \N__19642\,
            I => \N__19633\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__19639\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__3547\ : Odrv12
    port map (
            O => \N__19636\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__3546\ : Odrv4
    port map (
            O => \N__19633\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__3545\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19623\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__19623\,
            I => \N__19620\
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__19620\,
            I => \N_1318_tz_0\
        );

    \I__3542\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19614\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__19614\,
            I => \this_ppu.M_this_oam_ram_read_data_i_16\
        );

    \I__3540\ : InMux
    port map (
            O => \N__19611\,
            I => \N__19608\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__19608\,
            I => \N__19605\
        );

    \I__3538\ : Odrv4
    port map (
            O => \N__19605\,
            I => \this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0\
        );

    \I__3537\ : InMux
    port map (
            O => \N__19602\,
            I => \this_ppu.un2_vscroll_cry_0\
        );

    \I__3536\ : InMux
    port map (
            O => \N__19599\,
            I => \this_ppu.un2_vscroll_cry_1\
        );

    \I__3535\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19593\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__19593\,
            I => \this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0\
        );

    \I__3533\ : InMux
    port map (
            O => \N__19590\,
            I => \N__19587\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__19587\,
            I => \M_this_oam_ram_read_data_i_17\
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__19584\,
            I => \N__19581\
        );

    \I__3530\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19578\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__19578\,
            I => \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_5\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__19575\,
            I => \this_vga_signals.N_659_cascade_\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__19572\,
            I => \N_572_cascade_\
        );

    \I__3526\ : InMux
    port map (
            O => \N__19569\,
            I => \N__19566\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__19566\,
            I => \M_this_sprites_address_qc_2_0\
        );

    \I__3524\ : CascadeMux
    port map (
            O => \N__19563\,
            I => \N__19560\
        );

    \I__3523\ : InMux
    port map (
            O => \N__19560\,
            I => \N__19557\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__19557\,
            I => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_2\
        );

    \I__3521\ : InMux
    port map (
            O => \N__19554\,
            I => \N__19551\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__19551\,
            I => \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_3\
        );

    \I__3519\ : InMux
    port map (
            O => \N__19548\,
            I => \N__19545\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__19545\,
            I => \M_this_sprites_address_q_0_0_i_484\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__19542\,
            I => \M_this_sprites_address_qc_3_0_cascade_\
        );

    \I__3516\ : CascadeMux
    port map (
            O => \N__19539\,
            I => \N__19536\
        );

    \I__3515\ : InMux
    port map (
            O => \N__19536\,
            I => \N__19533\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__19533\,
            I => \M_this_substate_q_s_1\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__19530\,
            I => \M_this_sprites_address_q_0_0_i_480_cascade_\
        );

    \I__3512\ : InMux
    port map (
            O => \N__19527\,
            I => \N__19524\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__19524\,
            I => \M_this_sprites_address_qc_4_0\
        );

    \I__3510\ : InMux
    port map (
            O => \N__19521\,
            I => \N__19518\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__19518\,
            I => \N_511_1\
        );

    \I__3508\ : InMux
    port map (
            O => \N__19515\,
            I => \N__19512\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__19512\,
            I => \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_4\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__19509\,
            I => \N__19502\
        );

    \I__3505\ : InMux
    port map (
            O => \N__19508\,
            I => \N__19492\
        );

    \I__3504\ : InMux
    port map (
            O => \N__19507\,
            I => \N__19492\
        );

    \I__3503\ : InMux
    port map (
            O => \N__19506\,
            I => \N__19492\
        );

    \I__3502\ : InMux
    port map (
            O => \N__19505\,
            I => \N__19492\
        );

    \I__3501\ : InMux
    port map (
            O => \N__19502\,
            I => \N__19487\
        );

    \I__3500\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19487\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__19492\,
            I => \N__19481\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__19487\,
            I => \N__19478\
        );

    \I__3497\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19475\
        );

    \I__3496\ : InMux
    port map (
            O => \N__19485\,
            I => \N__19470\
        );

    \I__3495\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19470\
        );

    \I__3494\ : Span12Mux_v
    port map (
            O => \N__19481\,
            I => \N__19462\
        );

    \I__3493\ : Sp12to4
    port map (
            O => \N__19478\,
            I => \N__19462\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__19475\,
            I => \N__19462\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__19470\,
            I => \N__19459\
        );

    \I__3490\ : InMux
    port map (
            O => \N__19469\,
            I => \N__19456\
        );

    \I__3489\ : Span12Mux_v
    port map (
            O => \N__19462\,
            I => \N__19453\
        );

    \I__3488\ : Span12Mux_v
    port map (
            O => \N__19459\,
            I => \N__19450\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__19456\,
            I => \N__19447\
        );

    \I__3486\ : Odrv12
    port map (
            O => \N__19453\,
            I => rst_n_c
        );

    \I__3485\ : Odrv12
    port map (
            O => \N__19450\,
            I => rst_n_c
        );

    \I__3484\ : Odrv12
    port map (
            O => \N__19447\,
            I => rst_n_c
        );

    \I__3483\ : InMux
    port map (
            O => \N__19440\,
            I => \N__19437\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__19437\,
            I => \this_reset_cond.M_stage_qZ0Z_4\
        );

    \I__3481\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19431\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__19431\,
            I => \this_reset_cond.M_stage_qZ0Z_5\
        );

    \I__3479\ : InMux
    port map (
            O => \N__19428\,
            I => \N__19425\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__19425\,
            I => \N__19422\
        );

    \I__3477\ : Span4Mux_h
    port map (
            O => \N__19422\,
            I => \N__19419\
        );

    \I__3476\ : Span4Mux_v
    port map (
            O => \N__19419\,
            I => \N__19416\
        );

    \I__3475\ : Span4Mux_h
    port map (
            O => \N__19416\,
            I => \N__19413\
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__19413\,
            I => \this_sprites_ram.mem_out_bus6_0\
        );

    \I__3473\ : InMux
    port map (
            O => \N__19410\,
            I => \N__19407\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__19407\,
            I => \N__19404\
        );

    \I__3471\ : Span4Mux_v
    port map (
            O => \N__19404\,
            I => \N__19401\
        );

    \I__3470\ : Sp12to4
    port map (
            O => \N__19401\,
            I => \N__19398\
        );

    \I__3469\ : Odrv12
    port map (
            O => \N__19398\,
            I => \this_sprites_ram.mem_out_bus2_0\
        );

    \I__3468\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19392\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__19392\,
            I => \N__19389\
        );

    \I__3466\ : Span4Mux_v
    port map (
            O => \N__19389\,
            I => \N__19386\
        );

    \I__3465\ : Span4Mux_v
    port map (
            O => \N__19386\,
            I => \N__19383\
        );

    \I__3464\ : Span4Mux_h
    port map (
            O => \N__19383\,
            I => \N__19380\
        );

    \I__3463\ : Span4Mux_h
    port map (
            O => \N__19380\,
            I => \N__19377\
        );

    \I__3462\ : Odrv4
    port map (
            O => \N__19377\,
            I => \M_this_map_ram_read_data_5\
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__19374\,
            I => \N__19371\
        );

    \I__3460\ : InMux
    port map (
            O => \N__19371\,
            I => \N__19368\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__19368\,
            I => \N__19365\
        );

    \I__3458\ : Span4Mux_v
    port map (
            O => \N__19365\,
            I => \N__19362\
        );

    \I__3457\ : Sp12to4
    port map (
            O => \N__19362\,
            I => \N__19359\
        );

    \I__3456\ : Span12Mux_h
    port map (
            O => \N__19359\,
            I => \N__19356\
        );

    \I__3455\ : Odrv12
    port map (
            O => \N__19356\,
            I => \M_this_oam_ram_read_data_5\
        );

    \I__3454\ : InMux
    port map (
            O => \N__19353\,
            I => \N__19350\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__19350\,
            I => \N__19347\
        );

    \I__3452\ : Span4Mux_h
    port map (
            O => \N__19347\,
            I => \N__19344\
        );

    \I__3451\ : Sp12to4
    port map (
            O => \N__19344\,
            I => \N__19341\
        );

    \I__3450\ : Span12Mux_v
    port map (
            O => \N__19341\,
            I => \N__19338\
        );

    \I__3449\ : Odrv12
    port map (
            O => \N__19338\,
            I => \M_this_map_ram_read_data_7\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__19335\,
            I => \N__19332\
        );

    \I__3447\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19329\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__19329\,
            I => \N__19326\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__19326\,
            I => \N__19323\
        );

    \I__3444\ : Span4Mux_h
    port map (
            O => \N__19323\,
            I => \N__19320\
        );

    \I__3443\ : Sp12to4
    port map (
            O => \N__19320\,
            I => \N__19317\
        );

    \I__3442\ : Span12Mux_v
    port map (
            O => \N__19317\,
            I => \N__19314\
        );

    \I__3441\ : Odrv12
    port map (
            O => \N__19314\,
            I => \M_this_oam_ram_read_data_7\
        );

    \I__3440\ : InMux
    port map (
            O => \N__19311\,
            I => \N__19308\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__19308\,
            I => \N__19305\
        );

    \I__3438\ : Sp12to4
    port map (
            O => \N__19305\,
            I => \N__19302\
        );

    \I__3437\ : Span12Mux_v
    port map (
            O => \N__19302\,
            I => \N__19299\
        );

    \I__3436\ : Odrv12
    port map (
            O => \N__19299\,
            I => \this_sprites_ram.mem_out_bus4_2\
        );

    \I__3435\ : InMux
    port map (
            O => \N__19296\,
            I => \N__19293\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__19293\,
            I => \N__19290\
        );

    \I__3433\ : Span12Mux_v
    port map (
            O => \N__19290\,
            I => \N__19287\
        );

    \I__3432\ : Odrv12
    port map (
            O => \N__19287\,
            I => \this_sprites_ram.mem_out_bus0_2\
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__19284\,
            I => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_\
        );

    \I__3430\ : InMux
    port map (
            O => \N__19281\,
            I => \N__19278\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__19278\,
            I => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0\
        );

    \I__3428\ : InMux
    port map (
            O => \N__19275\,
            I => \N__19272\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__19272\,
            I => \N__19269\
        );

    \I__3426\ : Span4Mux_v
    port map (
            O => \N__19269\,
            I => \N__19266\
        );

    \I__3425\ : Span4Mux_h
    port map (
            O => \N__19266\,
            I => \N__19263\
        );

    \I__3424\ : Span4Mux_h
    port map (
            O => \N__19263\,
            I => \N__19260\
        );

    \I__3423\ : Span4Mux_v
    port map (
            O => \N__19260\,
            I => \N__19257\
        );

    \I__3422\ : Span4Mux_v
    port map (
            O => \N__19257\,
            I => \N__19254\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__19254\,
            I => \M_this_oam_ram_read_data_3\
        );

    \I__3420\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19248\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__19248\,
            I => \N__19245\
        );

    \I__3418\ : Span4Mux_v
    port map (
            O => \N__19245\,
            I => \N__19242\
        );

    \I__3417\ : Sp12to4
    port map (
            O => \N__19242\,
            I => \N__19239\
        );

    \I__3416\ : Span12Mux_h
    port map (
            O => \N__19239\,
            I => \N__19236\
        );

    \I__3415\ : Odrv12
    port map (
            O => \N__19236\,
            I => \M_this_map_ram_read_data_3\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__19233\,
            I => \N__19225\
        );

    \I__3413\ : CascadeMux
    port map (
            O => \N__19232\,
            I => \N__19222\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__19231\,
            I => \N__19219\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__19230\,
            I => \N__19216\
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__19229\,
            I => \N__19209\
        );

    \I__3409\ : CascadeMux
    port map (
            O => \N__19228\,
            I => \N__19206\
        );

    \I__3408\ : InMux
    port map (
            O => \N__19225\,
            I => \N__19203\
        );

    \I__3407\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19200\
        );

    \I__3406\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19197\
        );

    \I__3405\ : InMux
    port map (
            O => \N__19216\,
            I => \N__19194\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__19215\,
            I => \N__19190\
        );

    \I__3403\ : CascadeMux
    port map (
            O => \N__19214\,
            I => \N__19187\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__19213\,
            I => \N__19184\
        );

    \I__3401\ : CascadeMux
    port map (
            O => \N__19212\,
            I => \N__19178\
        );

    \I__3400\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19175\
        );

    \I__3399\ : InMux
    port map (
            O => \N__19206\,
            I => \N__19172\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__19203\,
            I => \N__19169\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__19200\,
            I => \N__19166\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__19197\,
            I => \N__19162\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__19194\,
            I => \N__19159\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__19193\,
            I => \N__19156\
        );

    \I__3393\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19153\
        );

    \I__3392\ : InMux
    port map (
            O => \N__19187\,
            I => \N__19150\
        );

    \I__3391\ : InMux
    port map (
            O => \N__19184\,
            I => \N__19147\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__19183\,
            I => \N__19143\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__19182\,
            I => \N__19140\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__19181\,
            I => \N__19137\
        );

    \I__3387\ : InMux
    port map (
            O => \N__19178\,
            I => \N__19134\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__19175\,
            I => \N__19127\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__19172\,
            I => \N__19127\
        );

    \I__3384\ : Span4Mux_v
    port map (
            O => \N__19169\,
            I => \N__19127\
        );

    \I__3383\ : Span4Mux_h
    port map (
            O => \N__19166\,
            I => \N__19124\
        );

    \I__3382\ : CascadeMux
    port map (
            O => \N__19165\,
            I => \N__19121\
        );

    \I__3381\ : Span4Mux_h
    port map (
            O => \N__19162\,
            I => \N__19118\
        );

    \I__3380\ : Span4Mux_h
    port map (
            O => \N__19159\,
            I => \N__19115\
        );

    \I__3379\ : InMux
    port map (
            O => \N__19156\,
            I => \N__19112\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__19153\,
            I => \N__19109\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__19150\,
            I => \N__19106\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__19147\,
            I => \N__19103\
        );

    \I__3375\ : CascadeMux
    port map (
            O => \N__19146\,
            I => \N__19100\
        );

    \I__3374\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19097\
        );

    \I__3373\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19094\
        );

    \I__3372\ : InMux
    port map (
            O => \N__19137\,
            I => \N__19091\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__19134\,
            I => \N__19088\
        );

    \I__3370\ : Span4Mux_v
    port map (
            O => \N__19127\,
            I => \N__19085\
        );

    \I__3369\ : Span4Mux_v
    port map (
            O => \N__19124\,
            I => \N__19082\
        );

    \I__3368\ : InMux
    port map (
            O => \N__19121\,
            I => \N__19079\
        );

    \I__3367\ : Span4Mux_h
    port map (
            O => \N__19118\,
            I => \N__19076\
        );

    \I__3366\ : Span4Mux_h
    port map (
            O => \N__19115\,
            I => \N__19073\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__19112\,
            I => \N__19070\
        );

    \I__3364\ : Span4Mux_h
    port map (
            O => \N__19109\,
            I => \N__19067\
        );

    \I__3363\ : Span4Mux_h
    port map (
            O => \N__19106\,
            I => \N__19064\
        );

    \I__3362\ : Span4Mux_h
    port map (
            O => \N__19103\,
            I => \N__19061\
        );

    \I__3361\ : InMux
    port map (
            O => \N__19100\,
            I => \N__19058\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__19097\,
            I => \N__19055\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__19094\,
            I => \N__19052\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__19091\,
            I => \N__19049\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__19088\,
            I => \N__19046\
        );

    \I__3356\ : Span4Mux_h
    port map (
            O => \N__19085\,
            I => \N__19041\
        );

    \I__3355\ : Span4Mux_v
    port map (
            O => \N__19082\,
            I => \N__19041\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__19079\,
            I => \N__19038\
        );

    \I__3353\ : Sp12to4
    port map (
            O => \N__19076\,
            I => \N__19031\
        );

    \I__3352\ : Sp12to4
    port map (
            O => \N__19073\,
            I => \N__19031\
        );

    \I__3351\ : Span12Mux_h
    port map (
            O => \N__19070\,
            I => \N__19031\
        );

    \I__3350\ : Span4Mux_v
    port map (
            O => \N__19067\,
            I => \N__19028\
        );

    \I__3349\ : Sp12to4
    port map (
            O => \N__19064\,
            I => \N__19023\
        );

    \I__3348\ : Sp12to4
    port map (
            O => \N__19061\,
            I => \N__19023\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__19058\,
            I => \N__19020\
        );

    \I__3346\ : Span12Mux_h
    port map (
            O => \N__19055\,
            I => \N__19013\
        );

    \I__3345\ : Span12Mux_h
    port map (
            O => \N__19052\,
            I => \N__19013\
        );

    \I__3344\ : Span12Mux_h
    port map (
            O => \N__19049\,
            I => \N__19013\
        );

    \I__3343\ : Span4Mux_h
    port map (
            O => \N__19046\,
            I => \N__19008\
        );

    \I__3342\ : Span4Mux_h
    port map (
            O => \N__19041\,
            I => \N__19008\
        );

    \I__3341\ : Sp12to4
    port map (
            O => \N__19038\,
            I => \N__18999\
        );

    \I__3340\ : Span12Mux_v
    port map (
            O => \N__19031\,
            I => \N__18999\
        );

    \I__3339\ : Sp12to4
    port map (
            O => \N__19028\,
            I => \N__18999\
        );

    \I__3338\ : Span12Mux_v
    port map (
            O => \N__19023\,
            I => \N__18999\
        );

    \I__3337\ : Odrv12
    port map (
            O => \N__19020\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__3336\ : Odrv12
    port map (
            O => \N__19013\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__3335\ : Odrv4
    port map (
            O => \N__19008\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__3334\ : Odrv12
    port map (
            O => \N__18999\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__3333\ : InMux
    port map (
            O => \N__18990\,
            I => \N__18987\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__18987\,
            I => \N__18984\
        );

    \I__3331\ : Span4Mux_v
    port map (
            O => \N__18984\,
            I => \N__18981\
        );

    \I__3330\ : Span4Mux_h
    port map (
            O => \N__18981\,
            I => \N__18978\
        );

    \I__3329\ : Odrv4
    port map (
            O => \N__18978\,
            I => \this_sprites_ram.mem_out_bus7_2\
        );

    \I__3328\ : InMux
    port map (
            O => \N__18975\,
            I => \N__18972\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__18972\,
            I => \N__18969\
        );

    \I__3326\ : Span4Mux_v
    port map (
            O => \N__18969\,
            I => \N__18966\
        );

    \I__3325\ : Span4Mux_h
    port map (
            O => \N__18966\,
            I => \N__18963\
        );

    \I__3324\ : Span4Mux_h
    port map (
            O => \N__18963\,
            I => \N__18960\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__18960\,
            I => \this_sprites_ram.mem_out_bus3_2\
        );

    \I__3322\ : InMux
    port map (
            O => \N__18957\,
            I => \N__18954\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__18954\,
            I => \this_reset_cond.M_stage_qZ0Z_8\
        );

    \I__3320\ : InMux
    port map (
            O => \N__18951\,
            I => \N__18947\
        );

    \I__3319\ : InMux
    port map (
            O => \N__18950\,
            I => \N__18941\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__18947\,
            I => \N__18938\
        );

    \I__3317\ : InMux
    port map (
            O => \N__18946\,
            I => \N__18935\
        );

    \I__3316\ : InMux
    port map (
            O => \N__18945\,
            I => \N__18932\
        );

    \I__3315\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18929\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__18941\,
            I => \N__18922\
        );

    \I__3313\ : Span4Mux_h
    port map (
            O => \N__18938\,
            I => \N__18922\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__18935\,
            I => \N__18922\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__18932\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__18929\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__18922\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__3308\ : InMux
    port map (
            O => \N__18915\,
            I => \N__18912\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__18912\,
            I => \N__18909\
        );

    \I__3306\ : Odrv4
    port map (
            O => \N__18909\,
            I => \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_5\
        );

    \I__3305\ : InMux
    port map (
            O => \N__18906\,
            I => \N__18902\
        );

    \I__3304\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18899\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__18902\,
            I => \N__18896\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__18899\,
            I => \N__18893\
        );

    \I__3301\ : Span4Mux_v
    port map (
            O => \N__18896\,
            I => \N__18890\
        );

    \I__3300\ : Span4Mux_h
    port map (
            O => \N__18893\,
            I => \N__18887\
        );

    \I__3299\ : Odrv4
    port map (
            O => \N__18890\,
            I => \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_4\
        );

    \I__3298\ : Odrv4
    port map (
            O => \N__18887\,
            I => \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_4\
        );

    \I__3297\ : InMux
    port map (
            O => \N__18882\,
            I => \N__18878\
        );

    \I__3296\ : InMux
    port map (
            O => \N__18881\,
            I => \N__18875\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__18878\,
            I => \N__18872\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__18875\,
            I => \N__18869\
        );

    \I__3293\ : Odrv4
    port map (
            O => \N__18872\,
            I => \this_ppu.M_count_d_0_sqmuxa_1\
        );

    \I__3292\ : Odrv4
    port map (
            O => \N__18869\,
            I => \this_ppu.M_count_d_0_sqmuxa_1\
        );

    \I__3291\ : CascadeMux
    port map (
            O => \N__18864\,
            I => \this_ppu.M_count_d_0_sqmuxa_1_cascade_\
        );

    \I__3290\ : InMux
    port map (
            O => \N__18861\,
            I => \N__18858\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__18858\,
            I => \N__18853\
        );

    \I__3288\ : InMux
    port map (
            O => \N__18857\,
            I => \N__18850\
        );

    \I__3287\ : InMux
    port map (
            O => \N__18856\,
            I => \N__18846\
        );

    \I__3286\ : Span4Mux_h
    port map (
            O => \N__18853\,
            I => \N__18841\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__18850\,
            I => \N__18841\
        );

    \I__3284\ : InMux
    port map (
            O => \N__18849\,
            I => \N__18838\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__18846\,
            I => \this_ppu.M_line_clk_out_0\
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__18841\,
            I => \this_ppu.M_line_clk_out_0\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__18838\,
            I => \this_ppu.M_line_clk_out_0\
        );

    \I__3280\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18823\
        );

    \I__3279\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18816\
        );

    \I__3278\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18816\
        );

    \I__3277\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18816\
        );

    \I__3276\ : InMux
    port map (
            O => \N__18827\,
            I => \N__18811\
        );

    \I__3275\ : InMux
    port map (
            O => \N__18826\,
            I => \N__18811\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__18823\,
            I => \this_ppu.N_1417_0\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__18816\,
            I => \this_ppu.N_1417_0\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__18811\,
            I => \this_ppu.N_1417_0\
        );

    \I__3271\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18801\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__18801\,
            I => \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__18798\,
            I => \this_ppu.N_1417_0_cascade_\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__18795\,
            I => \N__18791\
        );

    \I__3267\ : CascadeMux
    port map (
            O => \N__18794\,
            I => \N__18788\
        );

    \I__3266\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18779\
        );

    \I__3265\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18779\
        );

    \I__3264\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18779\
        );

    \I__3263\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18774\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__18779\,
            I => \N__18771\
        );

    \I__3261\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18766\
        );

    \I__3260\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18766\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__18774\,
            I => \this_ppu.un13_0\
        );

    \I__3258\ : Odrv4
    port map (
            O => \N__18771\,
            I => \this_ppu.un13_0\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__18766\,
            I => \this_ppu.un13_0\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__18759\,
            I => \N__18755\
        );

    \I__3255\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18752\
        );

    \I__3254\ : InMux
    port map (
            O => \N__18755\,
            I => \N__18748\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__18752\,
            I => \N__18745\
        );

    \I__3252\ : InMux
    port map (
            O => \N__18751\,
            I => \N__18742\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__18748\,
            I => \N__18739\
        );

    \I__3250\ : Span4Mux_h
    port map (
            O => \N__18745\,
            I => \N__18736\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__18742\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__18739\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__18736\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__3246\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18726\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__18726\,
            I => \N__18723\
        );

    \I__3244\ : Span4Mux_h
    port map (
            O => \N__18723\,
            I => \N__18720\
        );

    \I__3243\ : Span4Mux_h
    port map (
            O => \N__18720\,
            I => \N__18717\
        );

    \I__3242\ : Odrv4
    port map (
            O => \N__18717\,
            I => \this_sprites_ram.mem_out_bus6_2\
        );

    \I__3241\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18711\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__18711\,
            I => \N__18708\
        );

    \I__3239\ : Span4Mux_h
    port map (
            O => \N__18708\,
            I => \N__18705\
        );

    \I__3238\ : Span4Mux_h
    port map (
            O => \N__18705\,
            I => \N__18702\
        );

    \I__3237\ : Span4Mux_h
    port map (
            O => \N__18702\,
            I => \N__18699\
        );

    \I__3236\ : Odrv4
    port map (
            O => \N__18699\,
            I => \this_sprites_ram.mem_out_bus2_2\
        );

    \I__3235\ : InMux
    port map (
            O => \N__18696\,
            I => \N__18693\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__18693\,
            I => \N__18690\
        );

    \I__3233\ : Odrv12
    port map (
            O => \N__18690\,
            I => \this_reset_cond.M_stage_qZ0Z_3\
        );

    \I__3232\ : InMux
    port map (
            O => \N__18687\,
            I => \N__18684\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__18684\,
            I => \this_reset_cond.M_stage_qZ0Z_6\
        );

    \I__3230\ : InMux
    port map (
            O => \N__18681\,
            I => \N__18678\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__18678\,
            I => \this_reset_cond.M_stage_qZ0Z_7\
        );

    \I__3228\ : InMux
    port map (
            O => \N__18675\,
            I => \N__18672\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__18672\,
            I => \N__18669\
        );

    \I__3226\ : Odrv4
    port map (
            O => \N__18669\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__18666\,
            I => \this_ppu.M_state_q_srsts_i_2_1_cascade_\
        );

    \I__3224\ : InMux
    port map (
            O => \N__18663\,
            I => \N__18658\
        );

    \I__3223\ : InMux
    port map (
            O => \N__18662\,
            I => \N__18655\
        );

    \I__3222\ : InMux
    port map (
            O => \N__18661\,
            I => \N__18652\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__18658\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__18655\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__18652\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__18645\,
            I => \N__18641\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__18644\,
            I => \N__18638\
        );

    \I__3216\ : InMux
    port map (
            O => \N__18641\,
            I => \N__18635\
        );

    \I__3215\ : InMux
    port map (
            O => \N__18638\,
            I => \N__18632\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__18635\,
            I => \N__18629\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__18632\,
            I => \N__18626\
        );

    \I__3212\ : Span4Mux_h
    port map (
            O => \N__18629\,
            I => \N__18623\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__18626\,
            I => \this_ppu.M_count_qZ0Z_7\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__18623\,
            I => \this_ppu.M_count_qZ0Z_7\
        );

    \I__3209\ : CascadeMux
    port map (
            O => \N__18618\,
            I => \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_5_cascade_\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__18615\,
            I => \N__18612\
        );

    \I__3207\ : InMux
    port map (
            O => \N__18612\,
            I => \N__18609\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__18609\,
            I => \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__18606\,
            I => \N__18601\
        );

    \I__3204\ : InMux
    port map (
            O => \N__18605\,
            I => \N__18598\
        );

    \I__3203\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18595\
        );

    \I__3202\ : InMux
    port map (
            O => \N__18601\,
            I => \N__18592\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__18598\,
            I => \N__18589\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__18595\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__18592\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__18589\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__3197\ : InMux
    port map (
            O => \N__18582\,
            I => \N__18577\
        );

    \I__3196\ : InMux
    port map (
            O => \N__18581\,
            I => \N__18574\
        );

    \I__3195\ : InMux
    port map (
            O => \N__18580\,
            I => \N__18571\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__18577\,
            I => \N__18568\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__18574\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__18571\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__18568\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__3190\ : InMux
    port map (
            O => \N__18561\,
            I => \N__18558\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__18558\,
            I => \M_this_sprites_address_qc_8_0\
        );

    \I__3188\ : InMux
    port map (
            O => \N__18555\,
            I => \N__18552\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__18552\,
            I => \N__18549\
        );

    \I__3186\ : Span12Mux_s10_h
    port map (
            O => \N__18549\,
            I => \N__18546\
        );

    \I__3185\ : Odrv12
    port map (
            O => \N__18546\,
            I => \M_this_map_ram_write_data_3\
        );

    \I__3184\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18540\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__18540\,
            I => \N__18537\
        );

    \I__3182\ : Span12Mux_h
    port map (
            O => \N__18537\,
            I => \N__18534\
        );

    \I__3181\ : Odrv12
    port map (
            O => \N__18534\,
            I => \M_this_oam_ram_read_data_2\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__18531\,
            I => \N__18528\
        );

    \I__3179\ : InMux
    port map (
            O => \N__18528\,
            I => \N__18525\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__18525\,
            I => \N__18522\
        );

    \I__3177\ : Span4Mux_v
    port map (
            O => \N__18522\,
            I => \N__18519\
        );

    \I__3176\ : Sp12to4
    port map (
            O => \N__18519\,
            I => \N__18516\
        );

    \I__3175\ : Span12Mux_v
    port map (
            O => \N__18516\,
            I => \N__18513\
        );

    \I__3174\ : Odrv12
    port map (
            O => \N__18513\,
            I => \M_this_map_ram_read_data_2\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__18510\,
            I => \N__18507\
        );

    \I__3172\ : InMux
    port map (
            O => \N__18507\,
            I => \N__18502\
        );

    \I__3171\ : CascadeMux
    port map (
            O => \N__18506\,
            I => \N__18499\
        );

    \I__3170\ : CascadeMux
    port map (
            O => \N__18505\,
            I => \N__18496\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__18502\,
            I => \N__18488\
        );

    \I__3168\ : InMux
    port map (
            O => \N__18499\,
            I => \N__18485\
        );

    \I__3167\ : InMux
    port map (
            O => \N__18496\,
            I => \N__18482\
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__18495\,
            I => \N__18477\
        );

    \I__3165\ : CascadeMux
    port map (
            O => \N__18494\,
            I => \N__18474\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__18493\,
            I => \N__18471\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__18492\,
            I => \N__18468\
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__18491\,
            I => \N__18461\
        );

    \I__3161\ : Span4Mux_v
    port map (
            O => \N__18488\,
            I => \N__18452\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__18485\,
            I => \N__18452\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__18482\,
            I => \N__18452\
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__18481\,
            I => \N__18449\
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__18480\,
            I => \N__18446\
        );

    \I__3156\ : InMux
    port map (
            O => \N__18477\,
            I => \N__18443\
        );

    \I__3155\ : InMux
    port map (
            O => \N__18474\,
            I => \N__18440\
        );

    \I__3154\ : InMux
    port map (
            O => \N__18471\,
            I => \N__18437\
        );

    \I__3153\ : InMux
    port map (
            O => \N__18468\,
            I => \N__18434\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__18467\,
            I => \N__18431\
        );

    \I__3151\ : CascadeMux
    port map (
            O => \N__18466\,
            I => \N__18428\
        );

    \I__3150\ : CascadeMux
    port map (
            O => \N__18465\,
            I => \N__18425\
        );

    \I__3149\ : CascadeMux
    port map (
            O => \N__18464\,
            I => \N__18422\
        );

    \I__3148\ : InMux
    port map (
            O => \N__18461\,
            I => \N__18419\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__18460\,
            I => \N__18416\
        );

    \I__3146\ : CascadeMux
    port map (
            O => \N__18459\,
            I => \N__18413\
        );

    \I__3145\ : Span4Mux_v
    port map (
            O => \N__18452\,
            I => \N__18410\
        );

    \I__3144\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18407\
        );

    \I__3143\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18404\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__18443\,
            I => \N__18395\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__18440\,
            I => \N__18395\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__18437\,
            I => \N__18395\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__18434\,
            I => \N__18395\
        );

    \I__3138\ : InMux
    port map (
            O => \N__18431\,
            I => \N__18392\
        );

    \I__3137\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18389\
        );

    \I__3136\ : InMux
    port map (
            O => \N__18425\,
            I => \N__18386\
        );

    \I__3135\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18383\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__18419\,
            I => \N__18380\
        );

    \I__3133\ : InMux
    port map (
            O => \N__18416\,
            I => \N__18377\
        );

    \I__3132\ : InMux
    port map (
            O => \N__18413\,
            I => \N__18374\
        );

    \I__3131\ : Sp12to4
    port map (
            O => \N__18410\,
            I => \N__18369\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__18407\,
            I => \N__18369\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__18404\,
            I => \N__18366\
        );

    \I__3128\ : Span12Mux_s9_v
    port map (
            O => \N__18395\,
            I => \N__18351\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__18392\,
            I => \N__18351\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__18389\,
            I => \N__18351\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__18386\,
            I => \N__18351\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__18383\,
            I => \N__18351\
        );

    \I__3123\ : Sp12to4
    port map (
            O => \N__18380\,
            I => \N__18351\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__18377\,
            I => \N__18351\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__18374\,
            I => \N__18348\
        );

    \I__3120\ : Span12Mux_h
    port map (
            O => \N__18369\,
            I => \N__18345\
        );

    \I__3119\ : Span12Mux_s10_v
    port map (
            O => \N__18366\,
            I => \N__18338\
        );

    \I__3118\ : Span12Mux_v
    port map (
            O => \N__18351\,
            I => \N__18338\
        );

    \I__3117\ : Span12Mux_s7_h
    port map (
            O => \N__18348\,
            I => \N__18338\
        );

    \I__3116\ : Odrv12
    port map (
            O => \N__18345\,
            I => \M_this_ppu_sprites_addr_8\
        );

    \I__3115\ : Odrv12
    port map (
            O => \N__18338\,
            I => \M_this_ppu_sprites_addr_8\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__18333\,
            I => \N__18330\
        );

    \I__3113\ : InMux
    port map (
            O => \N__18330\,
            I => \N__18323\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__18329\,
            I => \N__18320\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__18328\,
            I => \N__18317\
        );

    \I__3110\ : CascadeMux
    port map (
            O => \N__18327\,
            I => \N__18313\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__18326\,
            I => \N__18309\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__18323\,
            I => \N__18304\
        );

    \I__3107\ : InMux
    port map (
            O => \N__18320\,
            I => \N__18301\
        );

    \I__3106\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18298\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__18316\,
            I => \N__18295\
        );

    \I__3104\ : InMux
    port map (
            O => \N__18313\,
            I => \N__18292\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__18312\,
            I => \N__18289\
        );

    \I__3102\ : InMux
    port map (
            O => \N__18309\,
            I => \N__18285\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__18308\,
            I => \N__18282\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__18307\,
            I => \N__18276\
        );

    \I__3099\ : Span4Mux_v
    port map (
            O => \N__18304\,
            I => \N__18267\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__18301\,
            I => \N__18267\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__18298\,
            I => \N__18267\
        );

    \I__3096\ : InMux
    port map (
            O => \N__18295\,
            I => \N__18264\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__18292\,
            I => \N__18261\
        );

    \I__3094\ : InMux
    port map (
            O => \N__18289\,
            I => \N__18258\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__18288\,
            I => \N__18255\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__18285\,
            I => \N__18252\
        );

    \I__3091\ : InMux
    port map (
            O => \N__18282\,
            I => \N__18249\
        );

    \I__3090\ : CascadeMux
    port map (
            O => \N__18281\,
            I => \N__18246\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__18280\,
            I => \N__18243\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__18279\,
            I => \N__18240\
        );

    \I__3087\ : InMux
    port map (
            O => \N__18276\,
            I => \N__18237\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__18275\,
            I => \N__18234\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__18274\,
            I => \N__18231\
        );

    \I__3084\ : Span4Mux_v
    port map (
            O => \N__18267\,
            I => \N__18226\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__18264\,
            I => \N__18226\
        );

    \I__3082\ : Span4Mux_v
    port map (
            O => \N__18261\,
            I => \N__18221\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__18258\,
            I => \N__18221\
        );

    \I__3080\ : InMux
    port map (
            O => \N__18255\,
            I => \N__18218\
        );

    \I__3079\ : Span4Mux_v
    port map (
            O => \N__18252\,
            I => \N__18213\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__18249\,
            I => \N__18213\
        );

    \I__3077\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18210\
        );

    \I__3076\ : InMux
    port map (
            O => \N__18243\,
            I => \N__18207\
        );

    \I__3075\ : InMux
    port map (
            O => \N__18240\,
            I => \N__18204\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__18237\,
            I => \N__18201\
        );

    \I__3073\ : InMux
    port map (
            O => \N__18234\,
            I => \N__18198\
        );

    \I__3072\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18195\
        );

    \I__3071\ : Span4Mux_v
    port map (
            O => \N__18226\,
            I => \N__18191\
        );

    \I__3070\ : Span4Mux_v
    port map (
            O => \N__18221\,
            I => \N__18188\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__18218\,
            I => \N__18185\
        );

    \I__3068\ : Span4Mux_v
    port map (
            O => \N__18213\,
            I => \N__18178\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__18210\,
            I => \N__18178\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__18207\,
            I => \N__18178\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__18204\,
            I => \N__18175\
        );

    \I__3064\ : Span4Mux_v
    port map (
            O => \N__18201\,
            I => \N__18168\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__18198\,
            I => \N__18168\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__18195\,
            I => \N__18168\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__18194\,
            I => \N__18165\
        );

    \I__3060\ : Span4Mux_v
    port map (
            O => \N__18191\,
            I => \N__18162\
        );

    \I__3059\ : Sp12to4
    port map (
            O => \N__18188\,
            I => \N__18155\
        );

    \I__3058\ : Span12Mux_h
    port map (
            O => \N__18185\,
            I => \N__18155\
        );

    \I__3057\ : Sp12to4
    port map (
            O => \N__18178\,
            I => \N__18155\
        );

    \I__3056\ : Span4Mux_v
    port map (
            O => \N__18175\,
            I => \N__18150\
        );

    \I__3055\ : Span4Mux_v
    port map (
            O => \N__18168\,
            I => \N__18150\
        );

    \I__3054\ : InMux
    port map (
            O => \N__18165\,
            I => \N__18147\
        );

    \I__3053\ : Sp12to4
    port map (
            O => \N__18162\,
            I => \N__18144\
        );

    \I__3052\ : Span12Mux_v
    port map (
            O => \N__18155\,
            I => \N__18137\
        );

    \I__3051\ : Sp12to4
    port map (
            O => \N__18150\,
            I => \N__18137\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__18147\,
            I => \N__18137\
        );

    \I__3049\ : Odrv12
    port map (
            O => \N__18144\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__3048\ : Odrv12
    port map (
            O => \N__18137\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__3047\ : InMux
    port map (
            O => \N__18132\,
            I => \N__18129\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__18129\,
            I => \N__18126\
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__18126\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__3044\ : InMux
    port map (
            O => \N__18123\,
            I => \N__18120\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__18120\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__18117\,
            I => \N__18107\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__18116\,
            I => \N__18103\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__18115\,
            I => \N__18095\
        );

    \I__3039\ : CascadeMux
    port map (
            O => \N__18114\,
            I => \N__18091\
        );

    \I__3038\ : CascadeMux
    port map (
            O => \N__18113\,
            I => \N__18088\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__18112\,
            I => \N__18085\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__18111\,
            I => \N__18082\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__18110\,
            I => \N__18079\
        );

    \I__3034\ : InMux
    port map (
            O => \N__18107\,
            I => \N__18076\
        );

    \I__3033\ : CascadeMux
    port map (
            O => \N__18106\,
            I => \N__18073\
        );

    \I__3032\ : InMux
    port map (
            O => \N__18103\,
            I => \N__18070\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__18102\,
            I => \N__18067\
        );

    \I__3030\ : CascadeMux
    port map (
            O => \N__18101\,
            I => \N__18064\
        );

    \I__3029\ : CascadeMux
    port map (
            O => \N__18100\,
            I => \N__18061\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__18099\,
            I => \N__18058\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__18098\,
            I => \N__18055\
        );

    \I__3026\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18052\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__18094\,
            I => \N__18049\
        );

    \I__3024\ : InMux
    port map (
            O => \N__18091\,
            I => \N__18046\
        );

    \I__3023\ : InMux
    port map (
            O => \N__18088\,
            I => \N__18043\
        );

    \I__3022\ : InMux
    port map (
            O => \N__18085\,
            I => \N__18040\
        );

    \I__3021\ : InMux
    port map (
            O => \N__18082\,
            I => \N__18037\
        );

    \I__3020\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18034\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__18076\,
            I => \N__18031\
        );

    \I__3018\ : InMux
    port map (
            O => \N__18073\,
            I => \N__18028\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__18070\,
            I => \N__18025\
        );

    \I__3016\ : InMux
    port map (
            O => \N__18067\,
            I => \N__18021\
        );

    \I__3015\ : InMux
    port map (
            O => \N__18064\,
            I => \N__18018\
        );

    \I__3014\ : InMux
    port map (
            O => \N__18061\,
            I => \N__18015\
        );

    \I__3013\ : InMux
    port map (
            O => \N__18058\,
            I => \N__18012\
        );

    \I__3012\ : InMux
    port map (
            O => \N__18055\,
            I => \N__18009\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__18052\,
            I => \N__18006\
        );

    \I__3010\ : InMux
    port map (
            O => \N__18049\,
            I => \N__18003\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__18046\,
            I => \N__17998\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__18043\,
            I => \N__17998\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__18040\,
            I => \N__17995\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__18037\,
            I => \N__17992\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__18034\,
            I => \N__17985\
        );

    \I__3004\ : Span4Mux_v
    port map (
            O => \N__18031\,
            I => \N__17985\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__18028\,
            I => \N__17985\
        );

    \I__3002\ : Span4Mux_v
    port map (
            O => \N__18025\,
            I => \N__17982\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__18024\,
            I => \N__17979\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__18021\,
            I => \N__17976\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__18018\,
            I => \N__17973\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__18015\,
            I => \N__17970\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__18012\,
            I => \N__17967\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__18009\,
            I => \N__17960\
        );

    \I__2995\ : Span4Mux_v
    port map (
            O => \N__18006\,
            I => \N__17960\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__18003\,
            I => \N__17960\
        );

    \I__2993\ : Span4Mux_v
    port map (
            O => \N__17998\,
            I => \N__17957\
        );

    \I__2992\ : Span4Mux_v
    port map (
            O => \N__17995\,
            I => \N__17954\
        );

    \I__2991\ : Span4Mux_h
    port map (
            O => \N__17992\,
            I => \N__17949\
        );

    \I__2990\ : Span4Mux_v
    port map (
            O => \N__17985\,
            I => \N__17949\
        );

    \I__2989\ : Span4Mux_h
    port map (
            O => \N__17982\,
            I => \N__17946\
        );

    \I__2988\ : InMux
    port map (
            O => \N__17979\,
            I => \N__17943\
        );

    \I__2987\ : Span4Mux_v
    port map (
            O => \N__17976\,
            I => \N__17940\
        );

    \I__2986\ : Span4Mux_h
    port map (
            O => \N__17973\,
            I => \N__17935\
        );

    \I__2985\ : Span4Mux_v
    port map (
            O => \N__17970\,
            I => \N__17935\
        );

    \I__2984\ : Span4Mux_h
    port map (
            O => \N__17967\,
            I => \N__17930\
        );

    \I__2983\ : Span4Mux_v
    port map (
            O => \N__17960\,
            I => \N__17930\
        );

    \I__2982\ : Span4Mux_h
    port map (
            O => \N__17957\,
            I => \N__17927\
        );

    \I__2981\ : Span4Mux_h
    port map (
            O => \N__17954\,
            I => \N__17924\
        );

    \I__2980\ : Span4Mux_h
    port map (
            O => \N__17949\,
            I => \N__17921\
        );

    \I__2979\ : Span4Mux_h
    port map (
            O => \N__17946\,
            I => \N__17918\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__17943\,
            I => \N__17915\
        );

    \I__2977\ : Span4Mux_h
    port map (
            O => \N__17940\,
            I => \N__17912\
        );

    \I__2976\ : Span4Mux_h
    port map (
            O => \N__17935\,
            I => \N__17909\
        );

    \I__2975\ : Span4Mux_h
    port map (
            O => \N__17930\,
            I => \N__17906\
        );

    \I__2974\ : Span4Mux_h
    port map (
            O => \N__17927\,
            I => \N__17897\
        );

    \I__2973\ : Span4Mux_h
    port map (
            O => \N__17924\,
            I => \N__17897\
        );

    \I__2972\ : Span4Mux_h
    port map (
            O => \N__17921\,
            I => \N__17897\
        );

    \I__2971\ : Span4Mux_v
    port map (
            O => \N__17918\,
            I => \N__17897\
        );

    \I__2970\ : Span12Mux_s8_h
    port map (
            O => \N__17915\,
            I => \N__17894\
        );

    \I__2969\ : Span4Mux_h
    port map (
            O => \N__17912\,
            I => \N__17887\
        );

    \I__2968\ : Span4Mux_h
    port map (
            O => \N__17909\,
            I => \N__17887\
        );

    \I__2967\ : Span4Mux_h
    port map (
            O => \N__17906\,
            I => \N__17887\
        );

    \I__2966\ : Sp12to4
    port map (
            O => \N__17897\,
            I => \N__17884\
        );

    \I__2965\ : Odrv12
    port map (
            O => \N__17894\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__2964\ : Odrv4
    port map (
            O => \N__17887\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__2963\ : Odrv12
    port map (
            O => \N__17884\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__17877\,
            I => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_7_cascade_\
        );

    \I__2961\ : CascadeMux
    port map (
            O => \N__17874\,
            I => \N_597_cascade_\
        );

    \I__2960\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17868\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__17868\,
            I => \M_this_sprites_address_qc_7_0\
        );

    \I__2958\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17862\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__17862\,
            I => \N_1298_tz_0\
        );

    \I__2956\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17856\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__17856\,
            I => \N__17853\
        );

    \I__2954\ : Odrv4
    port map (
            O => \N__17853\,
            I => \N_1294_tz_0\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__17850\,
            I => \N_602_cascade_\
        );

    \I__2952\ : InMux
    port map (
            O => \N__17847\,
            I => \N__17844\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__17844\,
            I => \this_ppu.M_count_q_RNO_0Z0Z_7\
        );

    \I__2950\ : InMux
    port map (
            O => \N__17841\,
            I => \N__17838\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__17838\,
            I => \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\
        );

    \I__2948\ : InMux
    port map (
            O => \N__17835\,
            I => \N__17830\
        );

    \I__2947\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17827\
        );

    \I__2946\ : InMux
    port map (
            O => \N__17833\,
            I => \N__17824\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__17830\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__17827\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__17824\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__2942\ : InMux
    port map (
            O => \N__17817\,
            I => \N__17814\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__17814\,
            I => \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__17811\,
            I => \N__17806\
        );

    \I__2939\ : InMux
    port map (
            O => \N__17810\,
            I => \N__17803\
        );

    \I__2938\ : InMux
    port map (
            O => \N__17809\,
            I => \N__17800\
        );

    \I__2937\ : InMux
    port map (
            O => \N__17806\,
            I => \N__17797\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__17803\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__17800\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__17797\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__2933\ : CascadeMux
    port map (
            O => \N__17790\,
            I => \N__17787\
        );

    \I__2932\ : InMux
    port map (
            O => \N__17787\,
            I => \N__17784\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__17784\,
            I => \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__17781\,
            I => \N__17777\
        );

    \I__2929\ : InMux
    port map (
            O => \N__17780\,
            I => \N__17773\
        );

    \I__2928\ : InMux
    port map (
            O => \N__17777\,
            I => \N__17770\
        );

    \I__2927\ : InMux
    port map (
            O => \N__17776\,
            I => \N__17767\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__17773\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__17770\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__17767\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__17760\,
            I => \N__17753\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__17759\,
            I => \N__17750\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__17758\,
            I => \N__17745\
        );

    \I__2920\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17742\
        );

    \I__2919\ : InMux
    port map (
            O => \N__17756\,
            I => \N__17739\
        );

    \I__2918\ : InMux
    port map (
            O => \N__17753\,
            I => \N__17736\
        );

    \I__2917\ : InMux
    port map (
            O => \N__17750\,
            I => \N__17733\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__17749\,
            I => \N__17729\
        );

    \I__2915\ : InMux
    port map (
            O => \N__17748\,
            I => \N__17726\
        );

    \I__2914\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17723\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__17742\,
            I => \N__17716\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__17739\,
            I => \N__17716\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__17736\,
            I => \N__17716\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__17733\,
            I => \N__17713\
        );

    \I__2909\ : InMux
    port map (
            O => \N__17732\,
            I => \N__17710\
        );

    \I__2908\ : InMux
    port map (
            O => \N__17729\,
            I => \N__17707\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__17726\,
            I => \N__17704\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__17723\,
            I => \N__17697\
        );

    \I__2905\ : Span4Mux_v
    port map (
            O => \N__17716\,
            I => \N__17697\
        );

    \I__2904\ : Span4Mux_v
    port map (
            O => \N__17713\,
            I => \N__17697\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__17710\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__17707\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2901\ : Odrv12
    port map (
            O => \N__17704\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__17697\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2899\ : CEMux
    port map (
            O => \N__17688\,
            I => \N__17678\
        );

    \I__2898\ : InMux
    port map (
            O => \N__17687\,
            I => \N__17664\
        );

    \I__2897\ : InMux
    port map (
            O => \N__17686\,
            I => \N__17664\
        );

    \I__2896\ : InMux
    port map (
            O => \N__17685\,
            I => \N__17659\
        );

    \I__2895\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17659\
        );

    \I__2894\ : InMux
    port map (
            O => \N__17683\,
            I => \N__17654\
        );

    \I__2893\ : InMux
    port map (
            O => \N__17682\,
            I => \N__17654\
        );

    \I__2892\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17651\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__17678\,
            I => \N__17648\
        );

    \I__2890\ : InMux
    port map (
            O => \N__17677\,
            I => \N__17639\
        );

    \I__2889\ : InMux
    port map (
            O => \N__17676\,
            I => \N__17639\
        );

    \I__2888\ : InMux
    port map (
            O => \N__17675\,
            I => \N__17639\
        );

    \I__2887\ : InMux
    port map (
            O => \N__17674\,
            I => \N__17639\
        );

    \I__2886\ : InMux
    port map (
            O => \N__17673\,
            I => \N__17632\
        );

    \I__2885\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17632\
        );

    \I__2884\ : InMux
    port map (
            O => \N__17671\,
            I => \N__17632\
        );

    \I__2883\ : InMux
    port map (
            O => \N__17670\,
            I => \N__17629\
        );

    \I__2882\ : CEMux
    port map (
            O => \N__17669\,
            I => \N__17624\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__17664\,
            I => \N__17621\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__17659\,
            I => \N__17616\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__17654\,
            I => \N__17616\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__17651\,
            I => \N__17611\
        );

    \I__2877\ : Span4Mux_v
    port map (
            O => \N__17648\,
            I => \N__17608\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__17639\,
            I => \N__17601\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__17632\,
            I => \N__17601\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__17629\,
            I => \N__17601\
        );

    \I__2873\ : InMux
    port map (
            O => \N__17628\,
            I => \N__17596\
        );

    \I__2872\ : InMux
    port map (
            O => \N__17627\,
            I => \N__17596\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__17624\,
            I => \N__17589\
        );

    \I__2870\ : Span4Mux_h
    port map (
            O => \N__17621\,
            I => \N__17589\
        );

    \I__2869\ : Span4Mux_v
    port map (
            O => \N__17616\,
            I => \N__17589\
        );

    \I__2868\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17586\
        );

    \I__2867\ : InMux
    port map (
            O => \N__17614\,
            I => \N__17583\
        );

    \I__2866\ : Span4Mux_v
    port map (
            O => \N__17611\,
            I => \N__17574\
        );

    \I__2865\ : Span4Mux_v
    port map (
            O => \N__17608\,
            I => \N__17574\
        );

    \I__2864\ : Span4Mux_v
    port map (
            O => \N__17601\,
            I => \N__17574\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__17596\,
            I => \N__17574\
        );

    \I__2862\ : Odrv4
    port map (
            O => \N__17589\,
            I => \this_vga_signals.GZ0Z_394\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__17586\,
            I => \this_vga_signals.GZ0Z_394\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__17583\,
            I => \this_vga_signals.GZ0Z_394\
        );

    \I__2859\ : Odrv4
    port map (
            O => \N__17574\,
            I => \this_vga_signals.GZ0Z_394\
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__17565\,
            I => \N__17562\
        );

    \I__2857\ : InMux
    port map (
            O => \N__17562\,
            I => \N__17557\
        );

    \I__2856\ : InMux
    port map (
            O => \N__17561\,
            I => \N__17552\
        );

    \I__2855\ : InMux
    port map (
            O => \N__17560\,
            I => \N__17549\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__17557\,
            I => \N__17545\
        );

    \I__2853\ : InMux
    port map (
            O => \N__17556\,
            I => \N__17540\
        );

    \I__2852\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17540\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__17552\,
            I => \N__17537\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__17549\,
            I => \N__17534\
        );

    \I__2849\ : InMux
    port map (
            O => \N__17548\,
            I => \N__17531\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__17545\,
            I => \N__17522\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__17540\,
            I => \N__17522\
        );

    \I__2846\ : Span4Mux_h
    port map (
            O => \N__17537\,
            I => \N__17522\
        );

    \I__2845\ : Span4Mux_v
    port map (
            O => \N__17534\,
            I => \N__17522\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__17531\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2843\ : Odrv4
    port map (
            O => \N__17522\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2842\ : SRMux
    port map (
            O => \N__17517\,
            I => \N__17512\
        );

    \I__2841\ : SRMux
    port map (
            O => \N__17516\,
            I => \N__17509\
        );

    \I__2840\ : SRMux
    port map (
            O => \N__17515\,
            I => \N__17506\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__17512\,
            I => \N__17501\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__17509\,
            I => \N__17501\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__17506\,
            I => \N__17498\
        );

    \I__2836\ : Span4Mux_v
    port map (
            O => \N__17501\,
            I => \N__17494\
        );

    \I__2835\ : Span4Mux_h
    port map (
            O => \N__17498\,
            I => \N__17491\
        );

    \I__2834\ : InMux
    port map (
            O => \N__17497\,
            I => \N__17488\
        );

    \I__2833\ : Span4Mux_h
    port map (
            O => \N__17494\,
            I => \N__17484\
        );

    \I__2832\ : Span4Mux_h
    port map (
            O => \N__17491\,
            I => \N__17481\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__17488\,
            I => \N__17478\
        );

    \I__2830\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17475\
        );

    \I__2829\ : Odrv4
    port map (
            O => \N__17484\,
            I => \this_vga_signals.M_vcounter_q_501_0\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__17481\,
            I => \this_vga_signals.M_vcounter_q_501_0\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__17478\,
            I => \this_vga_signals.M_vcounter_q_501_0\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__17475\,
            I => \this_vga_signals.M_vcounter_q_501_0\
        );

    \I__2825\ : InMux
    port map (
            O => \N__17466\,
            I => \N__17463\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__17463\,
            I => \N__17460\
        );

    \I__2823\ : Odrv12
    port map (
            O => \N__17460\,
            I => \this_delay_clk.M_pipe_qZ0Z_1\
        );

    \I__2822\ : InMux
    port map (
            O => \N__17457\,
            I => \N__17454\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__17454\,
            I => \this_delay_clk.M_pipe_qZ0Z_2\
        );

    \I__2820\ : CEMux
    port map (
            O => \N__17451\,
            I => \N__17447\
        );

    \I__2819\ : CEMux
    port map (
            O => \N__17450\,
            I => \N__17444\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__17447\,
            I => \N__17439\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__17444\,
            I => \N__17439\
        );

    \I__2816\ : Span4Mux_v
    port map (
            O => \N__17439\,
            I => \N__17436\
        );

    \I__2815\ : Span4Mux_h
    port map (
            O => \N__17436\,
            I => \N__17433\
        );

    \I__2814\ : Span4Mux_h
    port map (
            O => \N__17433\,
            I => \N__17430\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__17430\,
            I => \this_sprites_ram.mem_WE_10\
        );

    \I__2812\ : InMux
    port map (
            O => \N__17427\,
            I => \N__17424\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__17424\,
            I => \N__17418\
        );

    \I__2810\ : InMux
    port map (
            O => \N__17423\,
            I => \N__17413\
        );

    \I__2809\ : InMux
    port map (
            O => \N__17422\,
            I => \N__17413\
        );

    \I__2808\ : InMux
    port map (
            O => \N__17421\,
            I => \N__17408\
        );

    \I__2807\ : Span4Mux_v
    port map (
            O => \N__17418\,
            I => \N__17401\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__17413\,
            I => \N__17401\
        );

    \I__2805\ : InMux
    port map (
            O => \N__17412\,
            I => \N__17396\
        );

    \I__2804\ : InMux
    port map (
            O => \N__17411\,
            I => \N__17396\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__17408\,
            I => \N__17392\
        );

    \I__2802\ : InMux
    port map (
            O => \N__17407\,
            I => \N__17389\
        );

    \I__2801\ : InMux
    port map (
            O => \N__17406\,
            I => \N__17386\
        );

    \I__2800\ : Span4Mux_h
    port map (
            O => \N__17401\,
            I => \N__17383\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__17396\,
            I => \N__17380\
        );

    \I__2798\ : InMux
    port map (
            O => \N__17395\,
            I => \N__17377\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__17392\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__17389\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__17386\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__17383\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2793\ : Odrv4
    port map (
            O => \N__17380\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__17377\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__17364\,
            I => \M_this_vga_signals_line_clk_0_cascade_\
        );

    \I__2790\ : InMux
    port map (
            O => \N__17361\,
            I => \this_ppu.un1_M_count_q_1_cry_0_s1\
        );

    \I__2789\ : InMux
    port map (
            O => \N__17358\,
            I => \this_ppu.un1_M_count_q_1_cry_1_s1\
        );

    \I__2788\ : InMux
    port map (
            O => \N__17355\,
            I => \this_ppu.un1_M_count_q_1_cry_2_s1\
        );

    \I__2787\ : InMux
    port map (
            O => \N__17352\,
            I => \this_ppu.un1_M_count_q_1_cry_3_s1\
        );

    \I__2786\ : InMux
    port map (
            O => \N__17349\,
            I => \this_ppu.un1_M_count_q_1_cry_4_s1\
        );

    \I__2785\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17343\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__17343\,
            I => \N__17340\
        );

    \I__2783\ : Odrv12
    port map (
            O => \N__17340\,
            I => \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\
        );

    \I__2782\ : InMux
    port map (
            O => \N__17337\,
            I => \this_ppu.un1_M_count_q_1_cry_5_s1\
        );

    \I__2781\ : InMux
    port map (
            O => \N__17334\,
            I => \this_ppu.un1_M_count_q_1_cry_6_s1\
        );

    \I__2780\ : InMux
    port map (
            O => \N__17331\,
            I => \N__17328\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__17328\,
            I => \N__17319\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__17327\,
            I => \N__17316\
        );

    \I__2777\ : InMux
    port map (
            O => \N__17326\,
            I => \N__17299\
        );

    \I__2776\ : InMux
    port map (
            O => \N__17325\,
            I => \N__17294\
        );

    \I__2775\ : InMux
    port map (
            O => \N__17324\,
            I => \N__17294\
        );

    \I__2774\ : InMux
    port map (
            O => \N__17323\,
            I => \N__17289\
        );

    \I__2773\ : InMux
    port map (
            O => \N__17322\,
            I => \N__17289\
        );

    \I__2772\ : Span4Mux_v
    port map (
            O => \N__17319\,
            I => \N__17286\
        );

    \I__2771\ : InMux
    port map (
            O => \N__17316\,
            I => \N__17283\
        );

    \I__2770\ : InMux
    port map (
            O => \N__17315\,
            I => \N__17277\
        );

    \I__2769\ : InMux
    port map (
            O => \N__17314\,
            I => \N__17272\
        );

    \I__2768\ : InMux
    port map (
            O => \N__17313\,
            I => \N__17272\
        );

    \I__2767\ : InMux
    port map (
            O => \N__17312\,
            I => \N__17265\
        );

    \I__2766\ : InMux
    port map (
            O => \N__17311\,
            I => \N__17265\
        );

    \I__2765\ : InMux
    port map (
            O => \N__17310\,
            I => \N__17265\
        );

    \I__2764\ : InMux
    port map (
            O => \N__17309\,
            I => \N__17260\
        );

    \I__2763\ : InMux
    port map (
            O => \N__17308\,
            I => \N__17260\
        );

    \I__2762\ : InMux
    port map (
            O => \N__17307\,
            I => \N__17250\
        );

    \I__2761\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17250\
        );

    \I__2760\ : InMux
    port map (
            O => \N__17305\,
            I => \N__17250\
        );

    \I__2759\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17250\
        );

    \I__2758\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17245\
        );

    \I__2757\ : InMux
    port map (
            O => \N__17302\,
            I => \N__17245\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__17299\,
            I => \N__17229\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__17294\,
            I => \N__17229\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__17289\,
            I => \N__17229\
        );

    \I__2753\ : Span4Mux_h
    port map (
            O => \N__17286\,
            I => \N__17229\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__17283\,
            I => \N__17229\
        );

    \I__2751\ : InMux
    port map (
            O => \N__17282\,
            I => \N__17222\
        );

    \I__2750\ : InMux
    port map (
            O => \N__17281\,
            I => \N__17222\
        );

    \I__2749\ : InMux
    port map (
            O => \N__17280\,
            I => \N__17222\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__17277\,
            I => \N__17219\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__17272\,
            I => \N__17212\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__17265\,
            I => \N__17212\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__17260\,
            I => \N__17212\
        );

    \I__2744\ : InMux
    port map (
            O => \N__17259\,
            I => \N__17209\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__17250\,
            I => \N__17206\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__17245\,
            I => \N__17203\
        );

    \I__2741\ : InMux
    port map (
            O => \N__17244\,
            I => \N__17192\
        );

    \I__2740\ : InMux
    port map (
            O => \N__17243\,
            I => \N__17192\
        );

    \I__2739\ : InMux
    port map (
            O => \N__17242\,
            I => \N__17192\
        );

    \I__2738\ : InMux
    port map (
            O => \N__17241\,
            I => \N__17192\
        );

    \I__2737\ : InMux
    port map (
            O => \N__17240\,
            I => \N__17192\
        );

    \I__2736\ : Span4Mux_v
    port map (
            O => \N__17229\,
            I => \N__17189\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__17222\,
            I => \N__17186\
        );

    \I__2734\ : Span4Mux_v
    port map (
            O => \N__17219\,
            I => \N__17181\
        );

    \I__2733\ : Span4Mux_v
    port map (
            O => \N__17212\,
            I => \N__17181\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__17209\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2731\ : Odrv4
    port map (
            O => \N__17206\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2730\ : Odrv4
    port map (
            O => \N__17203\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__17192\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__17189\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__17186\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__17181\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2725\ : InMux
    port map (
            O => \N__17166\,
            I => \N__17157\
        );

    \I__2724\ : InMux
    port map (
            O => \N__17165\,
            I => \N__17154\
        );

    \I__2723\ : InMux
    port map (
            O => \N__17164\,
            I => \N__17144\
        );

    \I__2722\ : InMux
    port map (
            O => \N__17163\,
            I => \N__17144\
        );

    \I__2721\ : InMux
    port map (
            O => \N__17162\,
            I => \N__17144\
        );

    \I__2720\ : InMux
    port map (
            O => \N__17161\,
            I => \N__17144\
        );

    \I__2719\ : InMux
    port map (
            O => \N__17160\,
            I => \N__17135\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__17157\,
            I => \N__17130\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__17154\,
            I => \N__17130\
        );

    \I__2716\ : InMux
    port map (
            O => \N__17153\,
            I => \N__17127\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__17144\,
            I => \N__17124\
        );

    \I__2714\ : InMux
    port map (
            O => \N__17143\,
            I => \N__17119\
        );

    \I__2713\ : InMux
    port map (
            O => \N__17142\,
            I => \N__17119\
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__17141\,
            I => \N__17115\
        );

    \I__2711\ : InMux
    port map (
            O => \N__17140\,
            I => \N__17109\
        );

    \I__2710\ : InMux
    port map (
            O => \N__17139\,
            I => \N__17109\
        );

    \I__2709\ : InMux
    port map (
            O => \N__17138\,
            I => \N__17106\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__17135\,
            I => \N__17101\
        );

    \I__2707\ : Span4Mux_v
    port map (
            O => \N__17130\,
            I => \N__17101\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__17127\,
            I => \N__17094\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__17124\,
            I => \N__17094\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__17119\,
            I => \N__17094\
        );

    \I__2703\ : InMux
    port map (
            O => \N__17118\,
            I => \N__17091\
        );

    \I__2702\ : InMux
    port map (
            O => \N__17115\,
            I => \N__17086\
        );

    \I__2701\ : InMux
    port map (
            O => \N__17114\,
            I => \N__17086\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__17109\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__17106\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__17101\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__17094\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__17091\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__17086\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__17073\,
            I => \N__17070\
        );

    \I__2693\ : InMux
    port map (
            O => \N__17070\,
            I => \N__17067\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__17067\,
            I => \this_vga_signals.vaddress_0_0_6\
        );

    \I__2691\ : InMux
    port map (
            O => \N__17064\,
            I => \N__17059\
        );

    \I__2690\ : InMux
    port map (
            O => \N__17063\,
            I => \N__17053\
        );

    \I__2689\ : InMux
    port map (
            O => \N__17062\,
            I => \N__17053\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__17059\,
            I => \N__17050\
        );

    \I__2687\ : InMux
    port map (
            O => \N__17058\,
            I => \N__17046\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__17053\,
            I => \N__17042\
        );

    \I__2685\ : Span4Mux_h
    port map (
            O => \N__17050\,
            I => \N__17039\
        );

    \I__2684\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17036\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__17046\,
            I => \N__17033\
        );

    \I__2682\ : InMux
    port map (
            O => \N__17045\,
            I => \N__17030\
        );

    \I__2681\ : Span4Mux_v
    port map (
            O => \N__17042\,
            I => \N__17023\
        );

    \I__2680\ : Span4Mux_h
    port map (
            O => \N__17039\,
            I => \N__17020\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__17036\,
            I => \N__17017\
        );

    \I__2678\ : Span4Mux_v
    port map (
            O => \N__17033\,
            I => \N__17012\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__17030\,
            I => \N__17012\
        );

    \I__2676\ : InMux
    port map (
            O => \N__17029\,
            I => \N__17009\
        );

    \I__2675\ : InMux
    port map (
            O => \N__17028\,
            I => \N__17004\
        );

    \I__2674\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17004\
        );

    \I__2673\ : InMux
    port map (
            O => \N__17026\,
            I => \N__17001\
        );

    \I__2672\ : Odrv4
    port map (
            O => \N__17023\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__17020\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__2670\ : Odrv4
    port map (
            O => \N__17017\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__2669\ : Odrv4
    port map (
            O => \N__17012\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__17009\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__17004\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__17001\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__2665\ : InMux
    port map (
            O => \N__16986\,
            I => \N__16977\
        );

    \I__2664\ : InMux
    port map (
            O => \N__16985\,
            I => \N__16974\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__16984\,
            I => \N__16966\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__16983\,
            I => \N__16963\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__16982\,
            I => \N__16958\
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__16981\,
            I => \N__16954\
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__16980\,
            I => \N__16949\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__16977\,
            I => \N__16942\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__16974\,
            I => \N__16942\
        );

    \I__2656\ : InMux
    port map (
            O => \N__16973\,
            I => \N__16939\
        );

    \I__2655\ : InMux
    port map (
            O => \N__16972\,
            I => \N__16936\
        );

    \I__2654\ : InMux
    port map (
            O => \N__16971\,
            I => \N__16933\
        );

    \I__2653\ : InMux
    port map (
            O => \N__16970\,
            I => \N__16924\
        );

    \I__2652\ : InMux
    port map (
            O => \N__16969\,
            I => \N__16924\
        );

    \I__2651\ : InMux
    port map (
            O => \N__16966\,
            I => \N__16924\
        );

    \I__2650\ : InMux
    port map (
            O => \N__16963\,
            I => \N__16919\
        );

    \I__2649\ : InMux
    port map (
            O => \N__16962\,
            I => \N__16919\
        );

    \I__2648\ : InMux
    port map (
            O => \N__16961\,
            I => \N__16914\
        );

    \I__2647\ : InMux
    port map (
            O => \N__16958\,
            I => \N__16914\
        );

    \I__2646\ : InMux
    port map (
            O => \N__16957\,
            I => \N__16911\
        );

    \I__2645\ : InMux
    port map (
            O => \N__16954\,
            I => \N__16903\
        );

    \I__2644\ : InMux
    port map (
            O => \N__16953\,
            I => \N__16903\
        );

    \I__2643\ : InMux
    port map (
            O => \N__16952\,
            I => \N__16898\
        );

    \I__2642\ : InMux
    port map (
            O => \N__16949\,
            I => \N__16898\
        );

    \I__2641\ : InMux
    port map (
            O => \N__16948\,
            I => \N__16895\
        );

    \I__2640\ : InMux
    port map (
            O => \N__16947\,
            I => \N__16892\
        );

    \I__2639\ : Span4Mux_v
    port map (
            O => \N__16942\,
            I => \N__16889\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__16939\,
            I => \N__16882\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__16936\,
            I => \N__16882\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__16933\,
            I => \N__16882\
        );

    \I__2635\ : InMux
    port map (
            O => \N__16932\,
            I => \N__16879\
        );

    \I__2634\ : InMux
    port map (
            O => \N__16931\,
            I => \N__16876\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__16924\,
            I => \N__16871\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__16919\,
            I => \N__16871\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__16914\,
            I => \N__16866\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__16911\,
            I => \N__16866\
        );

    \I__2629\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16863\
        );

    \I__2628\ : InMux
    port map (
            O => \N__16909\,
            I => \N__16860\
        );

    \I__2627\ : InMux
    port map (
            O => \N__16908\,
            I => \N__16857\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__16903\,
            I => \N__16848\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__16898\,
            I => \N__16848\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__16895\,
            I => \N__16848\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__16892\,
            I => \N__16848\
        );

    \I__2622\ : Span4Mux_h
    port map (
            O => \N__16889\,
            I => \N__16843\
        );

    \I__2621\ : Span4Mux_v
    port map (
            O => \N__16882\,
            I => \N__16843\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__16879\,
            I => \N__16832\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__16876\,
            I => \N__16832\
        );

    \I__2618\ : Span4Mux_v
    port map (
            O => \N__16871\,
            I => \N__16832\
        );

    \I__2617\ : Span4Mux_h
    port map (
            O => \N__16866\,
            I => \N__16832\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__16863\,
            I => \N__16832\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__16860\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__16857\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2613\ : Odrv12
    port map (
            O => \N__16848\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2612\ : Odrv4
    port map (
            O => \N__16843\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__16832\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__16821\,
            I => \N__16815\
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__16820\,
            I => \N__16812\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__16819\,
            I => \N__16806\
        );

    \I__2607\ : InMux
    port map (
            O => \N__16818\,
            I => \N__16799\
        );

    \I__2606\ : InMux
    port map (
            O => \N__16815\,
            I => \N__16799\
        );

    \I__2605\ : InMux
    port map (
            O => \N__16812\,
            I => \N__16799\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__16811\,
            I => \N__16796\
        );

    \I__2603\ : CascadeMux
    port map (
            O => \N__16810\,
            I => \N__16785\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__16809\,
            I => \N__16780\
        );

    \I__2601\ : InMux
    port map (
            O => \N__16806\,
            I => \N__16775\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__16799\,
            I => \N__16772\
        );

    \I__2599\ : InMux
    port map (
            O => \N__16796\,
            I => \N__16767\
        );

    \I__2598\ : InMux
    port map (
            O => \N__16795\,
            I => \N__16767\
        );

    \I__2597\ : InMux
    port map (
            O => \N__16794\,
            I => \N__16761\
        );

    \I__2596\ : CascadeMux
    port map (
            O => \N__16793\,
            I => \N__16758\
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__16792\,
            I => \N__16751\
        );

    \I__2594\ : InMux
    port map (
            O => \N__16791\,
            I => \N__16747\
        );

    \I__2593\ : InMux
    port map (
            O => \N__16790\,
            I => \N__16744\
        );

    \I__2592\ : InMux
    port map (
            O => \N__16789\,
            I => \N__16741\
        );

    \I__2591\ : InMux
    port map (
            O => \N__16788\,
            I => \N__16738\
        );

    \I__2590\ : InMux
    port map (
            O => \N__16785\,
            I => \N__16733\
        );

    \I__2589\ : InMux
    port map (
            O => \N__16784\,
            I => \N__16733\
        );

    \I__2588\ : InMux
    port map (
            O => \N__16783\,
            I => \N__16729\
        );

    \I__2587\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16722\
        );

    \I__2586\ : InMux
    port map (
            O => \N__16779\,
            I => \N__16722\
        );

    \I__2585\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16722\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__16775\,
            I => \N__16711\
        );

    \I__2583\ : Span4Mux_h
    port map (
            O => \N__16772\,
            I => \N__16711\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__16767\,
            I => \N__16711\
        );

    \I__2581\ : InMux
    port map (
            O => \N__16766\,
            I => \N__16708\
        );

    \I__2580\ : InMux
    port map (
            O => \N__16765\,
            I => \N__16703\
        );

    \I__2579\ : InMux
    port map (
            O => \N__16764\,
            I => \N__16703\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__16761\,
            I => \N__16700\
        );

    \I__2577\ : InMux
    port map (
            O => \N__16758\,
            I => \N__16697\
        );

    \I__2576\ : InMux
    port map (
            O => \N__16757\,
            I => \N__16690\
        );

    \I__2575\ : InMux
    port map (
            O => \N__16756\,
            I => \N__16690\
        );

    \I__2574\ : InMux
    port map (
            O => \N__16755\,
            I => \N__16690\
        );

    \I__2573\ : InMux
    port map (
            O => \N__16754\,
            I => \N__16683\
        );

    \I__2572\ : InMux
    port map (
            O => \N__16751\,
            I => \N__16683\
        );

    \I__2571\ : InMux
    port map (
            O => \N__16750\,
            I => \N__16683\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__16747\,
            I => \N__16676\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__16744\,
            I => \N__16676\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__16741\,
            I => \N__16676\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__16738\,
            I => \N__16671\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__16733\,
            I => \N__16671\
        );

    \I__2565\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16668\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__16729\,
            I => \N__16665\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__16722\,
            I => \N__16662\
        );

    \I__2562\ : InMux
    port map (
            O => \N__16721\,
            I => \N__16655\
        );

    \I__2561\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16655\
        );

    \I__2560\ : InMux
    port map (
            O => \N__16719\,
            I => \N__16655\
        );

    \I__2559\ : InMux
    port map (
            O => \N__16718\,
            I => \N__16652\
        );

    \I__2558\ : Span4Mux_v
    port map (
            O => \N__16711\,
            I => \N__16649\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__16708\,
            I => \N__16640\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__16703\,
            I => \N__16640\
        );

    \I__2555\ : Span4Mux_v
    port map (
            O => \N__16700\,
            I => \N__16640\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__16697\,
            I => \N__16640\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__16690\,
            I => \N__16635\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__16683\,
            I => \N__16635\
        );

    \I__2551\ : Span4Mux_v
    port map (
            O => \N__16676\,
            I => \N__16632\
        );

    \I__2550\ : Span4Mux_v
    port map (
            O => \N__16671\,
            I => \N__16629\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__16668\,
            I => \N__16626\
        );

    \I__2548\ : Span4Mux_h
    port map (
            O => \N__16665\,
            I => \N__16619\
        );

    \I__2547\ : Span4Mux_h
    port map (
            O => \N__16662\,
            I => \N__16619\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__16655\,
            I => \N__16619\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__16652\,
            I => \N__16608\
        );

    \I__2544\ : Span4Mux_h
    port map (
            O => \N__16649\,
            I => \N__16608\
        );

    \I__2543\ : Span4Mux_v
    port map (
            O => \N__16640\,
            I => \N__16608\
        );

    \I__2542\ : Span4Mux_v
    port map (
            O => \N__16635\,
            I => \N__16608\
        );

    \I__2541\ : Span4Mux_h
    port map (
            O => \N__16632\,
            I => \N__16608\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__16629\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2539\ : Odrv12
    port map (
            O => \N__16626\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__16619\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__16608\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__16599\,
            I => \this_vga_signals.mult1_un54_sum_axb1_0_1_cascade_\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__16596\,
            I => \N__16593\
        );

    \I__2534\ : InMux
    port map (
            O => \N__16593\,
            I => \N__16586\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__16592\,
            I => \N__16583\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__16591\,
            I => \N__16579\
        );

    \I__2531\ : InMux
    port map (
            O => \N__16590\,
            I => \N__16576\
        );

    \I__2530\ : InMux
    port map (
            O => \N__16589\,
            I => \N__16573\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__16586\,
            I => \N__16570\
        );

    \I__2528\ : InMux
    port map (
            O => \N__16583\,
            I => \N__16563\
        );

    \I__2527\ : InMux
    port map (
            O => \N__16582\,
            I => \N__16563\
        );

    \I__2526\ : InMux
    port map (
            O => \N__16579\,
            I => \N__16563\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__16576\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__16573\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__16570\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__16563\,
            I => \this_vga_signals.mult1_un54_sum_c3_1\
        );

    \I__2521\ : InMux
    port map (
            O => \N__16554\,
            I => \N__16551\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__16551\,
            I => \N__16548\
        );

    \I__2519\ : Span4Mux_h
    port map (
            O => \N__16548\,
            I => \N__16545\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__16545\,
            I => \this_vga_signals.g0_0_0\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__16542\,
            I => \this_ppu.un13_0_cascade_\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__16539\,
            I => \this_ppu.M_line_clk_out_0_cascade_\
        );

    \I__2515\ : InMux
    port map (
            O => \N__16536\,
            I => \N__16532\
        );

    \I__2514\ : InMux
    port map (
            O => \N__16535\,
            I => \N__16529\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__16532\,
            I => \N__16525\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__16529\,
            I => \N__16522\
        );

    \I__2511\ : InMux
    port map (
            O => \N__16528\,
            I => \N__16519\
        );

    \I__2510\ : Span4Mux_v
    port map (
            O => \N__16525\,
            I => \N__16516\
        );

    \I__2509\ : Span4Mux_h
    port map (
            O => \N__16522\,
            I => \N__16513\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__16519\,
            I => \this_vga_signals.M_vcounter_d7lt9_1\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__16516\,
            I => \this_vga_signals.M_vcounter_d7lt9_1\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__16513\,
            I => \this_vga_signals.M_vcounter_d7lt9_1\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__16506\,
            I => \N__16502\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__16505\,
            I => \N__16496\
        );

    \I__2503\ : InMux
    port map (
            O => \N__16502\,
            I => \N__16491\
        );

    \I__2502\ : InMux
    port map (
            O => \N__16501\,
            I => \N__16488\
        );

    \I__2501\ : InMux
    port map (
            O => \N__16500\,
            I => \N__16485\
        );

    \I__2500\ : InMux
    port map (
            O => \N__16499\,
            I => \N__16482\
        );

    \I__2499\ : InMux
    port map (
            O => \N__16496\,
            I => \N__16479\
        );

    \I__2498\ : InMux
    port map (
            O => \N__16495\,
            I => \N__16473\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__16494\,
            I => \N__16469\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__16491\,
            I => \N__16461\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__16488\,
            I => \N__16461\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__16485\,
            I => \N__16456\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__16482\,
            I => \N__16456\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__16479\,
            I => \N__16453\
        );

    \I__2491\ : InMux
    port map (
            O => \N__16478\,
            I => \N__16448\
        );

    \I__2490\ : InMux
    port map (
            O => \N__16477\,
            I => \N__16448\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__16476\,
            I => \N__16443\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__16473\,
            I => \N__16440\
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__16472\,
            I => \N__16437\
        );

    \I__2486\ : InMux
    port map (
            O => \N__16469\,
            I => \N__16432\
        );

    \I__2485\ : InMux
    port map (
            O => \N__16468\,
            I => \N__16432\
        );

    \I__2484\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16427\
        );

    \I__2483\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16427\
        );

    \I__2482\ : Span4Mux_v
    port map (
            O => \N__16461\,
            I => \N__16418\
        );

    \I__2481\ : Span4Mux_v
    port map (
            O => \N__16456\,
            I => \N__16418\
        );

    \I__2480\ : Span4Mux_h
    port map (
            O => \N__16453\,
            I => \N__16418\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__16448\,
            I => \N__16418\
        );

    \I__2478\ : InMux
    port map (
            O => \N__16447\,
            I => \N__16411\
        );

    \I__2477\ : InMux
    port map (
            O => \N__16446\,
            I => \N__16411\
        );

    \I__2476\ : InMux
    port map (
            O => \N__16443\,
            I => \N__16411\
        );

    \I__2475\ : Span4Mux_v
    port map (
            O => \N__16440\,
            I => \N__16407\
        );

    \I__2474\ : InMux
    port map (
            O => \N__16437\,
            I => \N__16404\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__16432\,
            I => \N__16401\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__16427\,
            I => \N__16396\
        );

    \I__2471\ : Span4Mux_h
    port map (
            O => \N__16418\,
            I => \N__16396\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__16411\,
            I => \N__16393\
        );

    \I__2469\ : InMux
    port map (
            O => \N__16410\,
            I => \N__16390\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__16407\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__16404\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__16401\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__16396\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2464\ : Odrv12
    port map (
            O => \N__16393\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__16390\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__16377\,
            I => \N__16372\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__16376\,
            I => \N__16369\
        );

    \I__2460\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16357\
        );

    \I__2459\ : InMux
    port map (
            O => \N__16372\,
            I => \N__16354\
        );

    \I__2458\ : InMux
    port map (
            O => \N__16369\,
            I => \N__16351\
        );

    \I__2457\ : InMux
    port map (
            O => \N__16368\,
            I => \N__16347\
        );

    \I__2456\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16344\
        );

    \I__2455\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16339\
        );

    \I__2454\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16339\
        );

    \I__2453\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16336\
        );

    \I__2452\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16332\
        );

    \I__2451\ : InMux
    port map (
            O => \N__16362\,
            I => \N__16327\
        );

    \I__2450\ : InMux
    port map (
            O => \N__16361\,
            I => \N__16327\
        );

    \I__2449\ : InMux
    port map (
            O => \N__16360\,
            I => \N__16324\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__16357\,
            I => \N__16321\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__16354\,
            I => \N__16318\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__16351\,
            I => \N__16315\
        );

    \I__2445\ : InMux
    port map (
            O => \N__16350\,
            I => \N__16312\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__16347\,
            I => \N__16303\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__16344\,
            I => \N__16303\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__16339\,
            I => \N__16303\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__16336\,
            I => \N__16303\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__16335\,
            I => \N__16298\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__16332\,
            I => \N__16291\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__16327\,
            I => \N__16291\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__16324\,
            I => \N__16291\
        );

    \I__2436\ : Span4Mux_v
    port map (
            O => \N__16321\,
            I => \N__16284\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__16318\,
            I => \N__16284\
        );

    \I__2434\ : Span4Mux_v
    port map (
            O => \N__16315\,
            I => \N__16284\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__16312\,
            I => \N__16279\
        );

    \I__2432\ : Span4Mux_v
    port map (
            O => \N__16303\,
            I => \N__16279\
        );

    \I__2431\ : InMux
    port map (
            O => \N__16302\,
            I => \N__16274\
        );

    \I__2430\ : InMux
    port map (
            O => \N__16301\,
            I => \N__16274\
        );

    \I__2429\ : InMux
    port map (
            O => \N__16298\,
            I => \N__16271\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__16291\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2427\ : Odrv4
    port map (
            O => \N__16284\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__16279\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__16274\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__16271\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__16260\,
            I => \N__16257\
        );

    \I__2422\ : InMux
    port map (
            O => \N__16257\,
            I => \N__16254\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__16254\,
            I => \this_vga_signals.un4_lvisibility_1\
        );

    \I__2420\ : InMux
    port map (
            O => \N__16251\,
            I => \N__16245\
        );

    \I__2419\ : InMux
    port map (
            O => \N__16250\,
            I => \N__16245\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__16245\,
            I => \N__16242\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__16242\,
            I => \N__16239\
        );

    \I__2416\ : Odrv4
    port map (
            O => \N__16239\,
            I => \this_vga_signals.line_clk_1\
        );

    \I__2415\ : InMux
    port map (
            O => \N__16236\,
            I => \N__16230\
        );

    \I__2414\ : InMux
    port map (
            O => \N__16235\,
            I => \N__16225\
        );

    \I__2413\ : InMux
    port map (
            O => \N__16234\,
            I => \N__16225\
        );

    \I__2412\ : InMux
    port map (
            O => \N__16233\,
            I => \N__16219\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__16230\,
            I => \N__16214\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__16225\,
            I => \N__16211\
        );

    \I__2409\ : InMux
    port map (
            O => \N__16224\,
            I => \N__16206\
        );

    \I__2408\ : InMux
    port map (
            O => \N__16223\,
            I => \N__16206\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__16222\,
            I => \N__16203\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__16219\,
            I => \N__16200\
        );

    \I__2405\ : InMux
    port map (
            O => \N__16218\,
            I => \N__16197\
        );

    \I__2404\ : InMux
    port map (
            O => \N__16217\,
            I => \N__16194\
        );

    \I__2403\ : Span4Mux_v
    port map (
            O => \N__16214\,
            I => \N__16189\
        );

    \I__2402\ : Span4Mux_v
    port map (
            O => \N__16211\,
            I => \N__16189\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__16206\,
            I => \N__16186\
        );

    \I__2400\ : InMux
    port map (
            O => \N__16203\,
            I => \N__16183\
        );

    \I__2399\ : Odrv4
    port map (
            O => \N__16200\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__16197\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__16194\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2396\ : Odrv4
    port map (
            O => \N__16189\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__16186\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__16183\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2393\ : CascadeMux
    port map (
            O => \N__16170\,
            I => \this_vga_signals.un4_lvisibility_1_cascade_\
        );

    \I__2392\ : InMux
    port map (
            O => \N__16167\,
            I => \N__16162\
        );

    \I__2391\ : InMux
    port map (
            O => \N__16166\,
            I => \N__16158\
        );

    \I__2390\ : InMux
    port map (
            O => \N__16165\,
            I => \N__16155\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__16162\,
            I => \N__16152\
        );

    \I__2388\ : InMux
    port map (
            O => \N__16161\,
            I => \N__16149\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__16158\,
            I => \N__16143\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__16155\,
            I => \N__16143\
        );

    \I__2385\ : Span4Mux_v
    port map (
            O => \N__16152\,
            I => \N__16138\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__16149\,
            I => \N__16138\
        );

    \I__2383\ : InMux
    port map (
            O => \N__16148\,
            I => \N__16135\
        );

    \I__2382\ : Span4Mux_h
    port map (
            O => \N__16143\,
            I => \N__16132\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__16138\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__16135\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__16132\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__2378\ : InMux
    port map (
            O => \N__16125\,
            I => \N__16116\
        );

    \I__2377\ : InMux
    port map (
            O => \N__16124\,
            I => \N__16116\
        );

    \I__2376\ : InMux
    port map (
            O => \N__16123\,
            I => \N__16111\
        );

    \I__2375\ : InMux
    port map (
            O => \N__16122\,
            I => \N__16104\
        );

    \I__2374\ : InMux
    port map (
            O => \N__16121\,
            I => \N__16101\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__16116\,
            I => \N__16098\
        );

    \I__2372\ : InMux
    port map (
            O => \N__16115\,
            I => \N__16095\
        );

    \I__2371\ : InMux
    port map (
            O => \N__16114\,
            I => \N__16088\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__16111\,
            I => \N__16085\
        );

    \I__2369\ : InMux
    port map (
            O => \N__16110\,
            I => \N__16080\
        );

    \I__2368\ : InMux
    port map (
            O => \N__16109\,
            I => \N__16080\
        );

    \I__2367\ : InMux
    port map (
            O => \N__16108\,
            I => \N__16075\
        );

    \I__2366\ : InMux
    port map (
            O => \N__16107\,
            I => \N__16075\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__16104\,
            I => \N__16068\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__16101\,
            I => \N__16068\
        );

    \I__2363\ : Span4Mux_h
    port map (
            O => \N__16098\,
            I => \N__16068\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__16095\,
            I => \N__16065\
        );

    \I__2361\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16060\
        );

    \I__2360\ : InMux
    port map (
            O => \N__16093\,
            I => \N__16060\
        );

    \I__2359\ : InMux
    port map (
            O => \N__16092\,
            I => \N__16055\
        );

    \I__2358\ : InMux
    port map (
            O => \N__16091\,
            I => \N__16055\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__16088\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__16085\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__16080\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__16075\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__2353\ : Odrv4
    port map (
            O => \N__16068\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__2352\ : Odrv4
    port map (
            O => \N__16065\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__16060\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__16055\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__16038\,
            I => \this_vga_signals.mult1_un54_sum_c3_1_cascade_\
        );

    \I__2348\ : InMux
    port map (
            O => \N__16035\,
            I => \N__16032\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__16032\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0\
        );

    \I__2346\ : InMux
    port map (
            O => \N__16029\,
            I => \N__16023\
        );

    \I__2345\ : InMux
    port map (
            O => \N__16028\,
            I => \N__16018\
        );

    \I__2344\ : InMux
    port map (
            O => \N__16027\,
            I => \N__16018\
        );

    \I__2343\ : InMux
    port map (
            O => \N__16026\,
            I => \N__16015\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__16023\,
            I => \N__16012\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__16018\,
            I => \N__16009\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__16015\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__16012\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__2338\ : Odrv12
    port map (
            O => \N__16009\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__16002\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_cascade_\
        );

    \I__2336\ : InMux
    port map (
            O => \N__15999\,
            I => \N__15996\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__15996\,
            I => \N__15989\
        );

    \I__2334\ : InMux
    port map (
            O => \N__15995\,
            I => \N__15978\
        );

    \I__2333\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15978\
        );

    \I__2332\ : InMux
    port map (
            O => \N__15993\,
            I => \N__15978\
        );

    \I__2331\ : InMux
    port map (
            O => \N__15992\,
            I => \N__15975\
        );

    \I__2330\ : Span4Mux_h
    port map (
            O => \N__15989\,
            I => \N__15972\
        );

    \I__2329\ : InMux
    port map (
            O => \N__15988\,
            I => \N__15969\
        );

    \I__2328\ : InMux
    port map (
            O => \N__15987\,
            I => \N__15962\
        );

    \I__2327\ : InMux
    port map (
            O => \N__15986\,
            I => \N__15962\
        );

    \I__2326\ : InMux
    port map (
            O => \N__15985\,
            I => \N__15962\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__15978\,
            I => \this_vga_signals.mult1_un68_sum_axb1_654_ns\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__15975\,
            I => \this_vga_signals.mult1_un68_sum_axb1_654_ns\
        );

    \I__2323\ : Odrv4
    port map (
            O => \N__15972\,
            I => \this_vga_signals.mult1_un68_sum_axb1_654_ns\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__15969\,
            I => \this_vga_signals.mult1_un68_sum_axb1_654_ns\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__15962\,
            I => \this_vga_signals.mult1_un68_sum_axb1_654_ns\
        );

    \I__2320\ : InMux
    port map (
            O => \N__15951\,
            I => \N__15948\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__15948\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_x1\
        );

    \I__2318\ : CascadeMux
    port map (
            O => \N__15945\,
            I => \N__15942\
        );

    \I__2317\ : InMux
    port map (
            O => \N__15942\,
            I => \N__15939\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__15939\,
            I => \N__15936\
        );

    \I__2315\ : Odrv4
    port map (
            O => \N__15936\,
            I => \this_vga_signals.g0_i_i_a5_1_0_0_0\
        );

    \I__2314\ : InMux
    port map (
            O => \N__15933\,
            I => \N__15930\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__15930\,
            I => \this_vga_signals.g0_i_i_0_0_0\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__15927\,
            I => \this_vga_signals.vaddress_2_6_cascade_\
        );

    \I__2311\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15921\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__15921\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i_0\
        );

    \I__2309\ : CascadeMux
    port map (
            O => \N__15918\,
            I => \N__15915\
        );

    \I__2308\ : InMux
    port map (
            O => \N__15915\,
            I => \N__15912\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__15912\,
            I => \this_vga_signals.mult1_un54_sum_axb1_0_0\
        );

    \I__2306\ : InMux
    port map (
            O => \N__15909\,
            I => \N__15903\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__15908\,
            I => \N__15900\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__15907\,
            I => \N__15896\
        );

    \I__2303\ : InMux
    port map (
            O => \N__15906\,
            I => \N__15893\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__15903\,
            I => \N__15890\
        );

    \I__2301\ : InMux
    port map (
            O => \N__15900\,
            I => \N__15887\
        );

    \I__2300\ : InMux
    port map (
            O => \N__15899\,
            I => \N__15882\
        );

    \I__2299\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15882\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__15893\,
            I => \N__15877\
        );

    \I__2297\ : Span4Mux_v
    port map (
            O => \N__15890\,
            I => \N__15877\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__15887\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__15882\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__15877\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__2293\ : InMux
    port map (
            O => \N__15870\,
            I => \N__15867\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__15867\,
            I => \this_vga_signals.mult1_un47_sum_c3_0\
        );

    \I__2291\ : InMux
    port map (
            O => \N__15864\,
            I => \N__15861\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__15861\,
            I => \N__15856\
        );

    \I__2289\ : InMux
    port map (
            O => \N__15860\,
            I => \N__15851\
        );

    \I__2288\ : InMux
    port map (
            O => \N__15859\,
            I => \N__15851\
        );

    \I__2287\ : Odrv12
    port map (
            O => \N__15856\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i_0_0\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__15851\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i_0_0\
        );

    \I__2285\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15843\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__15843\,
            I => \N__15840\
        );

    \I__2283\ : Span4Mux_v
    port map (
            O => \N__15840\,
            I => \N__15837\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__15837\,
            I => \this_vga_signals.N_7_1_0\
        );

    \I__2281\ : InMux
    port map (
            O => \N__15834\,
            I => \bfn_15_21_0_\
        );

    \I__2280\ : InMux
    port map (
            O => \N__15831\,
            I => \N__15828\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__15828\,
            I => \N__15822\
        );

    \I__2278\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15819\
        );

    \I__2277\ : InMux
    port map (
            O => \N__15826\,
            I => \N__15815\
        );

    \I__2276\ : InMux
    port map (
            O => \N__15825\,
            I => \N__15811\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__15822\,
            I => \N__15805\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__15819\,
            I => \N__15805\
        );

    \I__2273\ : InMux
    port map (
            O => \N__15818\,
            I => \N__15802\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__15815\,
            I => \N__15799\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__15814\,
            I => \N__15795\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__15811\,
            I => \N__15791\
        );

    \I__2269\ : InMux
    port map (
            O => \N__15810\,
            I => \N__15788\
        );

    \I__2268\ : Span4Mux_h
    port map (
            O => \N__15805\,
            I => \N__15785\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__15802\,
            I => \N__15780\
        );

    \I__2266\ : Span4Mux_h
    port map (
            O => \N__15799\,
            I => \N__15780\
        );

    \I__2265\ : InMux
    port map (
            O => \N__15798\,
            I => \N__15775\
        );

    \I__2264\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15775\
        );

    \I__2263\ : InMux
    port map (
            O => \N__15794\,
            I => \N__15772\
        );

    \I__2262\ : Odrv12
    port map (
            O => \N__15791\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__15788\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__15785\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2259\ : Odrv4
    port map (
            O => \N__15780\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__15775\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__15772\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2256\ : CEMux
    port map (
            O => \N__15759\,
            I => \N__15756\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__15756\,
            I => \this_vga_signals.N_966_1\
        );

    \I__2254\ : CEMux
    port map (
            O => \N__15753\,
            I => \N__15749\
        );

    \I__2253\ : CEMux
    port map (
            O => \N__15752\,
            I => \N__15746\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__15749\,
            I => \N__15743\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__15746\,
            I => \N__15740\
        );

    \I__2250\ : Span4Mux_h
    port map (
            O => \N__15743\,
            I => \N__15737\
        );

    \I__2249\ : Span4Mux_v
    port map (
            O => \N__15740\,
            I => \N__15734\
        );

    \I__2248\ : Span4Mux_h
    port map (
            O => \N__15737\,
            I => \N__15731\
        );

    \I__2247\ : Span4Mux_h
    port map (
            O => \N__15734\,
            I => \N__15728\
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__15731\,
            I => \this_sprites_ram.mem_WE_8\
        );

    \I__2245\ : Odrv4
    port map (
            O => \N__15728\,
            I => \this_sprites_ram.mem_WE_8\
        );

    \I__2244\ : InMux
    port map (
            O => \N__15723\,
            I => \N__15720\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__15720\,
            I => \N__15717\
        );

    \I__2242\ : Odrv12
    port map (
            O => \N__15717\,
            I => \M_this_map_ram_write_data_2\
        );

    \I__2241\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15711\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__15711\,
            I => \N__15707\
        );

    \I__2239\ : InMux
    port map (
            O => \N__15710\,
            I => \N__15704\
        );

    \I__2238\ : Span4Mux_h
    port map (
            O => \N__15707\,
            I => \N__15698\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__15704\,
            I => \N__15698\
        );

    \I__2236\ : InMux
    port map (
            O => \N__15703\,
            I => \N__15695\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__15698\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__15695\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__2233\ : InMux
    port map (
            O => \N__15690\,
            I => \N__15687\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__15687\,
            I => \N__15684\
        );

    \I__2231\ : Span4Mux_h
    port map (
            O => \N__15684\,
            I => \N__15681\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__15681\,
            I => \this_vga_signals.g0_0_0_0\
        );

    \I__2229\ : InMux
    port map (
            O => \N__15678\,
            I => \N__15674\
        );

    \I__2228\ : InMux
    port map (
            O => \N__15677\,
            I => \N__15669\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__15674\,
            I => \N__15666\
        );

    \I__2226\ : InMux
    port map (
            O => \N__15673\,
            I => \N__15663\
        );

    \I__2225\ : InMux
    port map (
            O => \N__15672\,
            I => \N__15660\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__15669\,
            I => \N__15657\
        );

    \I__2223\ : Span4Mux_v
    port map (
            O => \N__15666\,
            I => \N__15649\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__15663\,
            I => \N__15649\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__15660\,
            I => \N__15646\
        );

    \I__2220\ : Span4Mux_h
    port map (
            O => \N__15657\,
            I => \N__15643\
        );

    \I__2219\ : InMux
    port map (
            O => \N__15656\,
            I => \N__15640\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__15655\,
            I => \N__15637\
        );

    \I__2217\ : InMux
    port map (
            O => \N__15654\,
            I => \N__15632\
        );

    \I__2216\ : Span4Mux_h
    port map (
            O => \N__15649\,
            I => \N__15629\
        );

    \I__2215\ : Span4Mux_h
    port map (
            O => \N__15646\,
            I => \N__15622\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__15643\,
            I => \N__15622\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__15640\,
            I => \N__15622\
        );

    \I__2212\ : InMux
    port map (
            O => \N__15637\,
            I => \N__15617\
        );

    \I__2211\ : InMux
    port map (
            O => \N__15636\,
            I => \N__15617\
        );

    \I__2210\ : InMux
    port map (
            O => \N__15635\,
            I => \N__15614\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__15632\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2208\ : Odrv4
    port map (
            O => \N__15629\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__15622\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__15617\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__15614\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__15603\,
            I => \this_vga_signals.g2_0_0_cascade_\
        );

    \I__2203\ : InMux
    port map (
            O => \N__15600\,
            I => \N__15594\
        );

    \I__2202\ : InMux
    port map (
            O => \N__15599\,
            I => \N__15591\
        );

    \I__2201\ : InMux
    port map (
            O => \N__15598\,
            I => \N__15588\
        );

    \I__2200\ : InMux
    port map (
            O => \N__15597\,
            I => \N__15585\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__15594\,
            I => \N__15582\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__15591\,
            I => \N__15575\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__15588\,
            I => \N__15575\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__15585\,
            I => \N__15572\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__15582\,
            I => \N__15569\
        );

    \I__2194\ : InMux
    port map (
            O => \N__15581\,
            I => \N__15563\
        );

    \I__2193\ : InMux
    port map (
            O => \N__15580\,
            I => \N__15560\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__15575\,
            I => \N__15557\
        );

    \I__2191\ : Span4Mux_h
    port map (
            O => \N__15572\,
            I => \N__15552\
        );

    \I__2190\ : Span4Mux_v
    port map (
            O => \N__15569\,
            I => \N__15552\
        );

    \I__2189\ : InMux
    port map (
            O => \N__15568\,
            I => \N__15549\
        );

    \I__2188\ : InMux
    port map (
            O => \N__15567\,
            I => \N__15544\
        );

    \I__2187\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15544\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__15563\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__15560\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__15557\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__15552\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__15549\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__15544\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2180\ : InMux
    port map (
            O => \N__15531\,
            I => \N__15528\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__15528\,
            I => \N__15525\
        );

    \I__2178\ : Span12Mux_h
    port map (
            O => \N__15525\,
            I => \N__15522\
        );

    \I__2177\ : Odrv12
    port map (
            O => \N__15522\,
            I => \this_vga_signals.g0_2_0\
        );

    \I__2176\ : InMux
    port map (
            O => \N__15519\,
            I => \N__15513\
        );

    \I__2175\ : InMux
    port map (
            O => \N__15518\,
            I => \N__15508\
        );

    \I__2174\ : InMux
    port map (
            O => \N__15517\,
            I => \N__15508\
        );

    \I__2173\ : InMux
    port map (
            O => \N__15516\,
            I => \N__15505\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__15513\,
            I => \this_vga_signals.mult1_un40_sum_axb1_0\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__15508\,
            I => \this_vga_signals.mult1_un40_sum_axb1_0\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__15505\,
            I => \this_vga_signals.mult1_un40_sum_axb1_0\
        );

    \I__2169\ : InMux
    port map (
            O => \N__15498\,
            I => \N__15495\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__15495\,
            I => \N__15491\
        );

    \I__2167\ : InMux
    port map (
            O => \N__15494\,
            I => \N__15486\
        );

    \I__2166\ : Span4Mux_v
    port map (
            O => \N__15491\,
            I => \N__15483\
        );

    \I__2165\ : InMux
    port map (
            O => \N__15490\,
            I => \N__15480\
        );

    \I__2164\ : InMux
    port map (
            O => \N__15489\,
            I => \N__15477\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__15486\,
            I => \this_vga_signals.SUM_2_i_1_0_3\
        );

    \I__2162\ : Odrv4
    port map (
            O => \N__15483\,
            I => \this_vga_signals.SUM_2_i_1_0_3\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__15480\,
            I => \this_vga_signals.SUM_2_i_1_0_3\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__15477\,
            I => \this_vga_signals.SUM_2_i_1_0_3\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__15468\,
            I => \N__15465\
        );

    \I__2158\ : InMux
    port map (
            O => \N__15465\,
            I => \N__15461\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__15464\,
            I => \N__15457\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__15461\,
            I => \N__15454\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__15460\,
            I => \N__15451\
        );

    \I__2154\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15448\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__15454\,
            I => \N__15445\
        );

    \I__2152\ : InMux
    port map (
            O => \N__15451\,
            I => \N__15442\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__15448\,
            I => \this_vga_signals.SUM_2_i_1_2_3\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__15445\,
            I => \this_vga_signals.SUM_2_i_1_2_3\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__15442\,
            I => \this_vga_signals.SUM_2_i_1_2_3\
        );

    \I__2148\ : InMux
    port map (
            O => \N__15435\,
            I => \N__15432\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__15432\,
            I => \N__15429\
        );

    \I__2146\ : Span4Mux_h
    port map (
            O => \N__15429\,
            I => \N__15423\
        );

    \I__2145\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15418\
        );

    \I__2144\ : InMux
    port map (
            O => \N__15427\,
            I => \N__15418\
        );

    \I__2143\ : InMux
    port map (
            O => \N__15426\,
            I => \N__15415\
        );

    \I__2142\ : Odrv4
    port map (
            O => \N__15423\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__15418\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__15415\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4\
        );

    \I__2139\ : InMux
    port map (
            O => \N__15408\,
            I => \N__15398\
        );

    \I__2138\ : InMux
    port map (
            O => \N__15407\,
            I => \N__15398\
        );

    \I__2137\ : InMux
    port map (
            O => \N__15406\,
            I => \N__15398\
        );

    \I__2136\ : InMux
    port map (
            O => \N__15405\,
            I => \N__15395\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__15398\,
            I => \N__15390\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__15395\,
            I => \N__15387\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__15394\,
            I => \N__15381\
        );

    \I__2132\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15378\
        );

    \I__2131\ : Span4Mux_v
    port map (
            O => \N__15390\,
            I => \N__15375\
        );

    \I__2130\ : Span4Mux_h
    port map (
            O => \N__15387\,
            I => \N__15372\
        );

    \I__2129\ : InMux
    port map (
            O => \N__15386\,
            I => \N__15369\
        );

    \I__2128\ : InMux
    port map (
            O => \N__15385\,
            I => \N__15362\
        );

    \I__2127\ : InMux
    port map (
            O => \N__15384\,
            I => \N__15362\
        );

    \I__2126\ : InMux
    port map (
            O => \N__15381\,
            I => \N__15362\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__15378\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__15375\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__15372\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__15369\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__15362\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__15351\,
            I => \this_vga_signals.vaddress_0_0_6_cascade_\
        );

    \I__2119\ : InMux
    port map (
            O => \N__15348\,
            I => \N__15345\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__15345\,
            I => \N__15342\
        );

    \I__2117\ : Span4Mux_v
    port map (
            O => \N__15342\,
            I => \N__15339\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__15339\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i_0_0\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__15336\,
            I => \N__15333\
        );

    \I__2114\ : InMux
    port map (
            O => \N__15333\,
            I => \N__15328\
        );

    \I__2113\ : InMux
    port map (
            O => \N__15332\,
            I => \N__15322\
        );

    \I__2112\ : InMux
    port map (
            O => \N__15331\,
            I => \N__15319\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__15328\,
            I => \N__15313\
        );

    \I__2110\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15310\
        );

    \I__2109\ : InMux
    port map (
            O => \N__15326\,
            I => \N__15307\
        );

    \I__2108\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15304\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__15322\,
            I => \N__15299\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__15319\,
            I => \N__15299\
        );

    \I__2105\ : InMux
    port map (
            O => \N__15318\,
            I => \N__15294\
        );

    \I__2104\ : InMux
    port map (
            O => \N__15317\,
            I => \N__15294\
        );

    \I__2103\ : InMux
    port map (
            O => \N__15316\,
            I => \N__15291\
        );

    \I__2102\ : Odrv4
    port map (
            O => \N__15313\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__15310\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__15307\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__15304\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2098\ : Odrv4
    port map (
            O => \N__15299\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__15294\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__15291\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2095\ : InMux
    port map (
            O => \N__15276\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__2094\ : InMux
    port map (
            O => \N__15273\,
            I => \N__15269\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__15272\,
            I => \N__15266\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__15269\,
            I => \N__15260\
        );

    \I__2091\ : InMux
    port map (
            O => \N__15266\,
            I => \N__15257\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__15265\,
            I => \N__15250\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__15264\,
            I => \N__15247\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__15263\,
            I => \N__15244\
        );

    \I__2087\ : Span4Mux_v
    port map (
            O => \N__15260\,
            I => \N__15239\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__15257\,
            I => \N__15239\
        );

    \I__2085\ : InMux
    port map (
            O => \N__15256\,
            I => \N__15236\
        );

    \I__2084\ : InMux
    port map (
            O => \N__15255\,
            I => \N__15232\
        );

    \I__2083\ : InMux
    port map (
            O => \N__15254\,
            I => \N__15229\
        );

    \I__2082\ : InMux
    port map (
            O => \N__15253\,
            I => \N__15220\
        );

    \I__2081\ : InMux
    port map (
            O => \N__15250\,
            I => \N__15220\
        );

    \I__2080\ : InMux
    port map (
            O => \N__15247\,
            I => \N__15220\
        );

    \I__2079\ : InMux
    port map (
            O => \N__15244\,
            I => \N__15220\
        );

    \I__2078\ : Span4Mux_h
    port map (
            O => \N__15239\,
            I => \N__15215\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__15236\,
            I => \N__15215\
        );

    \I__2076\ : InMux
    port map (
            O => \N__15235\,
            I => \N__15212\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__15232\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__15229\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__15220\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__15215\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__15212\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2070\ : InMux
    port map (
            O => \N__15201\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__2069\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15192\
        );

    \I__2068\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15187\
        );

    \I__2067\ : InMux
    port map (
            O => \N__15196\,
            I => \N__15182\
        );

    \I__2066\ : InMux
    port map (
            O => \N__15195\,
            I => \N__15182\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__15192\,
            I => \N__15174\
        );

    \I__2064\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15171\
        );

    \I__2063\ : InMux
    port map (
            O => \N__15190\,
            I => \N__15168\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__15187\,
            I => \N__15165\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__15182\,
            I => \N__15162\
        );

    \I__2060\ : InMux
    port map (
            O => \N__15181\,
            I => \N__15157\
        );

    \I__2059\ : InMux
    port map (
            O => \N__15180\,
            I => \N__15157\
        );

    \I__2058\ : InMux
    port map (
            O => \N__15179\,
            I => \N__15154\
        );

    \I__2057\ : InMux
    port map (
            O => \N__15178\,
            I => \N__15151\
        );

    \I__2056\ : InMux
    port map (
            O => \N__15177\,
            I => \N__15148\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__15174\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__15171\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__15168\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__15165\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__15162\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__15157\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__15154\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__15151\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__15148\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2046\ : InMux
    port map (
            O => \N__15129\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__2045\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15121\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__15125\,
            I => \N__15116\
        );

    \I__2043\ : InMux
    port map (
            O => \N__15124\,
            I => \N__15107\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__15121\,
            I => \N__15104\
        );

    \I__2041\ : InMux
    port map (
            O => \N__15120\,
            I => \N__15097\
        );

    \I__2040\ : InMux
    port map (
            O => \N__15119\,
            I => \N__15097\
        );

    \I__2039\ : InMux
    port map (
            O => \N__15116\,
            I => \N__15097\
        );

    \I__2038\ : InMux
    port map (
            O => \N__15115\,
            I => \N__15092\
        );

    \I__2037\ : InMux
    port map (
            O => \N__15114\,
            I => \N__15092\
        );

    \I__2036\ : InMux
    port map (
            O => \N__15113\,
            I => \N__15083\
        );

    \I__2035\ : InMux
    port map (
            O => \N__15112\,
            I => \N__15083\
        );

    \I__2034\ : InMux
    port map (
            O => \N__15111\,
            I => \N__15083\
        );

    \I__2033\ : InMux
    port map (
            O => \N__15110\,
            I => \N__15083\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__15107\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__15104\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__15097\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__15092\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__15083\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2027\ : InMux
    port map (
            O => \N__15072\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__2026\ : InMux
    port map (
            O => \N__15069\,
            I => \N__15066\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__15066\,
            I => \N__15060\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__15065\,
            I => \N__15051\
        );

    \I__2023\ : CascadeMux
    port map (
            O => \N__15064\,
            I => \N__15048\
        );

    \I__2022\ : InMux
    port map (
            O => \N__15063\,
            I => \N__15045\
        );

    \I__2021\ : Span4Mux_h
    port map (
            O => \N__15060\,
            I => \N__15042\
        );

    \I__2020\ : InMux
    port map (
            O => \N__15059\,
            I => \N__15037\
        );

    \I__2019\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15037\
        );

    \I__2018\ : InMux
    port map (
            O => \N__15057\,
            I => \N__15028\
        );

    \I__2017\ : InMux
    port map (
            O => \N__15056\,
            I => \N__15028\
        );

    \I__2016\ : InMux
    port map (
            O => \N__15055\,
            I => \N__15028\
        );

    \I__2015\ : InMux
    port map (
            O => \N__15054\,
            I => \N__15028\
        );

    \I__2014\ : InMux
    port map (
            O => \N__15051\,
            I => \N__15023\
        );

    \I__2013\ : InMux
    port map (
            O => \N__15048\,
            I => \N__15023\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__15045\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__15042\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__15037\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__15028\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__15023\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2007\ : InMux
    port map (
            O => \N__15012\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__2006\ : InMux
    port map (
            O => \N__15009\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__2005\ : InMux
    port map (
            O => \N__15006\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__2004\ : InMux
    port map (
            O => \N__15003\,
            I => \N__15000\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__15000\,
            I => \this_vga_signals.mult1_un54_sum_c3_1_0\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__14997\,
            I => \this_vga_signals.mult1_un54_sum_c3_1_0_cascade_\
        );

    \I__2001\ : InMux
    port map (
            O => \N__14994\,
            I => \N__14991\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__14991\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_1\
        );

    \I__1999\ : InMux
    port map (
            O => \N__14988\,
            I => \N__14982\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__14987\,
            I => \N__14977\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__14986\,
            I => \N__14974\
        );

    \I__1996\ : InMux
    port map (
            O => \N__14985\,
            I => \N__14969\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__14982\,
            I => \N__14966\
        );

    \I__1994\ : InMux
    port map (
            O => \N__14981\,
            I => \N__14963\
        );

    \I__1993\ : InMux
    port map (
            O => \N__14980\,
            I => \N__14960\
        );

    \I__1992\ : InMux
    port map (
            O => \N__14977\,
            I => \N__14955\
        );

    \I__1991\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14955\
        );

    \I__1990\ : CascadeMux
    port map (
            O => \N__14973\,
            I => \N__14952\
        );

    \I__1989\ : InMux
    port map (
            O => \N__14972\,
            I => \N__14949\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__14969\,
            I => \N__14939\
        );

    \I__1987\ : Span4Mux_h
    port map (
            O => \N__14966\,
            I => \N__14939\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__14963\,
            I => \N__14932\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__14960\,
            I => \N__14932\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__14955\,
            I => \N__14932\
        );

    \I__1983\ : InMux
    port map (
            O => \N__14952\,
            I => \N__14929\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__14949\,
            I => \N__14926\
        );

    \I__1981\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14923\
        );

    \I__1980\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14920\
        );

    \I__1979\ : InMux
    port map (
            O => \N__14946\,
            I => \N__14915\
        );

    \I__1978\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14915\
        );

    \I__1977\ : InMux
    port map (
            O => \N__14944\,
            I => \N__14912\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__14939\,
            I => \N__14909\
        );

    \I__1975\ : Span4Mux_v
    port map (
            O => \N__14932\,
            I => \N__14906\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__14929\,
            I => \N__14901\
        );

    \I__1973\ : Span4Mux_h
    port map (
            O => \N__14926\,
            I => \N__14901\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__14923\,
            I => \N__14896\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__14920\,
            I => \N__14896\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__14915\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__14912\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__14909\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__14906\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__14901\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1965\ : Odrv12
    port map (
            O => \N__14896\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1964\ : InMux
    port map (
            O => \N__14883\,
            I => \N__14880\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__14880\,
            I => \N__14877\
        );

    \I__1962\ : Span4Mux_h
    port map (
            O => \N__14877\,
            I => \N__14869\
        );

    \I__1961\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14864\
        );

    \I__1960\ : InMux
    port map (
            O => \N__14875\,
            I => \N__14864\
        );

    \I__1959\ : InMux
    port map (
            O => \N__14874\,
            I => \N__14861\
        );

    \I__1958\ : InMux
    port map (
            O => \N__14873\,
            I => \N__14858\
        );

    \I__1957\ : InMux
    port map (
            O => \N__14872\,
            I => \N__14855\
        );

    \I__1956\ : Span4Mux_v
    port map (
            O => \N__14869\,
            I => \N__14852\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__14864\,
            I => \N__14847\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__14861\,
            I => \N__14847\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__14858\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__14855\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__14852\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__1950\ : Odrv12
    port map (
            O => \N__14847\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__1949\ : InMux
    port map (
            O => \N__14838\,
            I => \N__14835\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__14835\,
            I => \this_vga_signals.mult1_un68_sum_axb1\
        );

    \I__1947\ : InMux
    port map (
            O => \N__14832\,
            I => \N__14829\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__14829\,
            I => \this_vga_signals.if_m5_s\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__14826\,
            I => \N__14822\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__14825\,
            I => \N__14819\
        );

    \I__1943\ : InMux
    port map (
            O => \N__14822\,
            I => \N__14816\
        );

    \I__1942\ : InMux
    port map (
            O => \N__14819\,
            I => \N__14813\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__14816\,
            I => \N__14810\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__14813\,
            I => \N__14805\
        );

    \I__1939\ : Span4Mux_v
    port map (
            O => \N__14810\,
            I => \N__14805\
        );

    \I__1938\ : Span4Mux_h
    port map (
            O => \N__14805\,
            I => \N__14802\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__14802\,
            I => \this_vga_signals.M_vcounter_d7lto8_1\
        );

    \I__1936\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14794\
        );

    \I__1935\ : InMux
    port map (
            O => \N__14798\,
            I => \N__14787\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__14797\,
            I => \N__14784\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__14794\,
            I => \N__14780\
        );

    \I__1932\ : InMux
    port map (
            O => \N__14793\,
            I => \N__14777\
        );

    \I__1931\ : InMux
    port map (
            O => \N__14792\,
            I => \N__14772\
        );

    \I__1930\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14772\
        );

    \I__1929\ : InMux
    port map (
            O => \N__14790\,
            I => \N__14767\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__14787\,
            I => \N__14764\
        );

    \I__1927\ : InMux
    port map (
            O => \N__14784\,
            I => \N__14759\
        );

    \I__1926\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14759\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__14780\,
            I => \N__14754\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__14777\,
            I => \N__14754\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__14772\,
            I => \N__14749\
        );

    \I__1922\ : InMux
    port map (
            O => \N__14771\,
            I => \N__14746\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__14770\,
            I => \N__14743\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__14767\,
            I => \N__14732\
        );

    \I__1919\ : Span4Mux_v
    port map (
            O => \N__14764\,
            I => \N__14732\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__14759\,
            I => \N__14732\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__14754\,
            I => \N__14732\
        );

    \I__1916\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14729\
        );

    \I__1915\ : InMux
    port map (
            O => \N__14752\,
            I => \N__14726\
        );

    \I__1914\ : Span4Mux_v
    port map (
            O => \N__14749\,
            I => \N__14721\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__14746\,
            I => \N__14721\
        );

    \I__1912\ : InMux
    port map (
            O => \N__14743\,
            I => \N__14718\
        );

    \I__1911\ : InMux
    port map (
            O => \N__14742\,
            I => \N__14713\
        );

    \I__1910\ : InMux
    port map (
            O => \N__14741\,
            I => \N__14713\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__14732\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__14729\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__14726\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__14721\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__14718\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__14713\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1903\ : IoInMux
    port map (
            O => \N__14700\,
            I => \N__14697\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__14697\,
            I => \N__14694\
        );

    \I__1901\ : IoSpan4Mux
    port map (
            O => \N__14694\,
            I => \N__14691\
        );

    \I__1900\ : Span4Mux_s3_v
    port map (
            O => \N__14691\,
            I => \N__14688\
        );

    \I__1899\ : Sp12to4
    port map (
            O => \N__14688\,
            I => \N__14684\
        );

    \I__1898\ : InMux
    port map (
            O => \N__14687\,
            I => \N__14681\
        );

    \I__1897\ : Span12Mux_v
    port map (
            O => \N__14684\,
            I => \N__14678\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__14681\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\
        );

    \I__1895\ : Odrv12
    port map (
            O => \N__14678\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\
        );

    \I__1894\ : InMux
    port map (
            O => \N__14673\,
            I => \N__14670\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__14670\,
            I => \this_vga_signals.M_hcounter_d7lto4_0\
        );

    \I__1892\ : InMux
    port map (
            O => \N__14667\,
            I => \N__14664\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__14664\,
            I => \N__14661\
        );

    \I__1890\ : Span4Mux_v
    port map (
            O => \N__14661\,
            I => \N__14658\
        );

    \I__1889\ : Sp12to4
    port map (
            O => \N__14658\,
            I => \N__14655\
        );

    \I__1888\ : Odrv12
    port map (
            O => \N__14655\,
            I => \this_sprites_ram.mem_out_bus7_0\
        );

    \I__1887\ : InMux
    port map (
            O => \N__14652\,
            I => \N__14649\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__14649\,
            I => \N__14646\
        );

    \I__1885\ : Span4Mux_h
    port map (
            O => \N__14646\,
            I => \N__14643\
        );

    \I__1884\ : Span4Mux_v
    port map (
            O => \N__14643\,
            I => \N__14640\
        );

    \I__1883\ : Span4Mux_h
    port map (
            O => \N__14640\,
            I => \N__14637\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__14637\,
            I => \this_sprites_ram.mem_out_bus3_0\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__14634\,
            I => \N__14631\
        );

    \I__1880\ : InMux
    port map (
            O => \N__14631\,
            I => \N__14627\
        );

    \I__1879\ : InMux
    port map (
            O => \N__14630\,
            I => \N__14621\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__14627\,
            I => \N__14618\
        );

    \I__1877\ : InMux
    port map (
            O => \N__14626\,
            I => \N__14615\
        );

    \I__1876\ : InMux
    port map (
            O => \N__14625\,
            I => \N__14610\
        );

    \I__1875\ : InMux
    port map (
            O => \N__14624\,
            I => \N__14610\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__14621\,
            I => \N__14605\
        );

    \I__1873\ : Span4Mux_h
    port map (
            O => \N__14618\,
            I => \N__14605\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__14615\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__14610\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__14605\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__14598\,
            I => \N__14595\
        );

    \I__1868\ : InMux
    port map (
            O => \N__14595\,
            I => \N__14592\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__14592\,
            I => \this_vga_signals.mult1_un68_sum_axb1_654_x0\
        );

    \I__1866\ : InMux
    port map (
            O => \N__14589\,
            I => \N__14586\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__14586\,
            I => \this_vga_signals.mult1_un68_sum_axb1_654_x1\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__14583\,
            I => \this_vga_signals.mult1_un68_sum_axb1_654_ns_cascade_\
        );

    \I__1863\ : InMux
    port map (
            O => \N__14580\,
            I => \N__14577\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__14577\,
            I => \this_vga_signals.if_m1_3\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__14574\,
            I => \this_vga_signals.if_m1_3_cascade_\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__14571\,
            I => \N__14568\
        );

    \I__1859\ : InMux
    port map (
            O => \N__14568\,
            I => \N__14565\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__14565\,
            I => \N__14562\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__14562\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x1\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__14559\,
            I => \N__14556\
        );

    \I__1855\ : InMux
    port map (
            O => \N__14556\,
            I => \N__14553\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__14553\,
            I => \N__14550\
        );

    \I__1853\ : Span4Mux_h
    port map (
            O => \N__14550\,
            I => \N__14547\
        );

    \I__1852\ : Odrv4
    port map (
            O => \N__14547\,
            I => \this_vga_signals.vaddress_0_6\
        );

    \I__1851\ : InMux
    port map (
            O => \N__14544\,
            I => \N__14541\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__14541\,
            I => \this_vga_signals.mult1_un47_sum_c3_1_0\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__14538\,
            I => \N__14533\
        );

    \I__1848\ : InMux
    port map (
            O => \N__14537\,
            I => \N__14529\
        );

    \I__1847\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14526\
        );

    \I__1846\ : InMux
    port map (
            O => \N__14533\,
            I => \N__14523\
        );

    \I__1845\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14520\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__14529\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__14526\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__14523\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__14520\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3\
        );

    \I__1840\ : InMux
    port map (
            O => \N__14511\,
            I => \N__14508\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__14508\,
            I => \this_vga_signals.g1\
        );

    \I__1838\ : InMux
    port map (
            O => \N__14505\,
            I => \N__14502\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__14502\,
            I => \N__14489\
        );

    \I__1836\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14484\
        );

    \I__1835\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14481\
        );

    \I__1834\ : InMux
    port map (
            O => \N__14499\,
            I => \N__14474\
        );

    \I__1833\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14474\
        );

    \I__1832\ : InMux
    port map (
            O => \N__14497\,
            I => \N__14474\
        );

    \I__1831\ : InMux
    port map (
            O => \N__14496\,
            I => \N__14467\
        );

    \I__1830\ : InMux
    port map (
            O => \N__14495\,
            I => \N__14467\
        );

    \I__1829\ : InMux
    port map (
            O => \N__14494\,
            I => \N__14467\
        );

    \I__1828\ : InMux
    port map (
            O => \N__14493\,
            I => \N__14462\
        );

    \I__1827\ : InMux
    port map (
            O => \N__14492\,
            I => \N__14462\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__14489\,
            I => \N__14459\
        );

    \I__1825\ : InMux
    port map (
            O => \N__14488\,
            I => \N__14454\
        );

    \I__1824\ : InMux
    port map (
            O => \N__14487\,
            I => \N__14454\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__14484\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__14481\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__14474\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__14467\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__14462\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__14459\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__14454\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__14439\,
            I => \this_vga_signals.g0_2_cascade_\
        );

    \I__1815\ : InMux
    port map (
            O => \N__14436\,
            I => \N__14433\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__14433\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0_0_1\
        );

    \I__1813\ : InMux
    port map (
            O => \N__14430\,
            I => \N__14427\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__14427\,
            I => \this_vga_signals.N_3_1_0\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__14424\,
            I => \this_vga_signals.N_11_0_0_cascade_\
        );

    \I__1810\ : InMux
    port map (
            O => \N__14421\,
            I => \N__14418\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__14418\,
            I => \this_vga_signals.N_4_1_0_0\
        );

    \I__1808\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14412\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__14412\,
            I => \N__14409\
        );

    \I__1806\ : Odrv4
    port map (
            O => \N__14409\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i_2\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__14406\,
            I => \N__14403\
        );

    \I__1804\ : InMux
    port map (
            O => \N__14403\,
            I => \N__14400\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__14400\,
            I => \N__14397\
        );

    \I__1802\ : Span4Mux_h
    port map (
            O => \N__14397\,
            I => \N__14393\
        );

    \I__1801\ : InMux
    port map (
            O => \N__14396\,
            I => \N__14390\
        );

    \I__1800\ : Odrv4
    port map (
            O => \N__14393\,
            I => \this_vga_signals.vaddress_3_6\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__14390\,
            I => \this_vga_signals.vaddress_3_6\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__14385\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i_2_cascade_\
        );

    \I__1797\ : InMux
    port map (
            O => \N__14382\,
            I => \N__14379\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__14379\,
            I => \this_vga_signals.mult1_un47_sum_c3_2\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__14376\,
            I => \this_vga_signals.mult1_un47_sum_c3_2_cascade_\
        );

    \I__1794\ : InMux
    port map (
            O => \N__14373\,
            I => \N__14370\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__14370\,
            I => \this_vga_signals.g0_1\
        );

    \I__1792\ : InMux
    port map (
            O => \N__14367\,
            I => \N__14361\
        );

    \I__1791\ : InMux
    port map (
            O => \N__14366\,
            I => \N__14356\
        );

    \I__1790\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14356\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__14364\,
            I => \N__14350\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__14361\,
            I => \N__14345\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__14356\,
            I => \N__14345\
        );

    \I__1786\ : InMux
    port map (
            O => \N__14355\,
            I => \N__14342\
        );

    \I__1785\ : InMux
    port map (
            O => \N__14354\,
            I => \N__14339\
        );

    \I__1784\ : InMux
    port map (
            O => \N__14353\,
            I => \N__14334\
        );

    \I__1783\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14334\
        );

    \I__1782\ : Span4Mux_h
    port map (
            O => \N__14345\,
            I => \N__14331\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__14342\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__14339\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__14334\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__14331\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__14322\,
            I => \this_vga_signals.vaddress_6_cascade_\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__14319\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_\
        );

    \I__1775\ : InMux
    port map (
            O => \N__14316\,
            I => \N__14313\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__14313\,
            I => \N__14310\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__14310\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_i\
        );

    \I__1772\ : InMux
    port map (
            O => \N__14307\,
            I => \N__14304\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__14304\,
            I => \N__14301\
        );

    \I__1770\ : Span4Mux_h
    port map (
            O => \N__14301\,
            I => \N__14296\
        );

    \I__1769\ : InMux
    port map (
            O => \N__14300\,
            I => \N__14293\
        );

    \I__1768\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14290\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__14296\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__14293\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__14290\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3\
        );

    \I__1764\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14280\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__14280\,
            I => \N__14277\
        );

    \I__1762\ : Span4Mux_v
    port map (
            O => \N__14277\,
            I => \N__14274\
        );

    \I__1761\ : Span4Mux_h
    port map (
            O => \N__14274\,
            I => \N__14270\
        );

    \I__1760\ : InMux
    port map (
            O => \N__14273\,
            I => \N__14267\
        );

    \I__1759\ : Odrv4
    port map (
            O => \N__14270\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__14267\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__1757\ : InMux
    port map (
            O => \N__14262\,
            I => \N__14259\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__14259\,
            I => \N__14256\
        );

    \I__1755\ : Span4Mux_v
    port map (
            O => \N__14256\,
            I => \N__14251\
        );

    \I__1754\ : InMux
    port map (
            O => \N__14255\,
            I => \N__14246\
        );

    \I__1753\ : InMux
    port map (
            O => \N__14254\,
            I => \N__14246\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__14251\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__14246\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__14241\,
            I => \N__14234\
        );

    \I__1749\ : InMux
    port map (
            O => \N__14240\,
            I => \N__14229\
        );

    \I__1748\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14229\
        );

    \I__1747\ : InMux
    port map (
            O => \N__14238\,
            I => \N__14226\
        );

    \I__1746\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14221\
        );

    \I__1745\ : InMux
    port map (
            O => \N__14234\,
            I => \N__14221\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__14229\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__14226\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__14221\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__14214\,
            I => \N__14210\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__14213\,
            I => \N__14207\
        );

    \I__1739\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14200\
        );

    \I__1738\ : InMux
    port map (
            O => \N__14207\,
            I => \N__14200\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__14206\,
            I => \N__14197\
        );

    \I__1736\ : InMux
    port map (
            O => \N__14205\,
            I => \N__14193\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__14200\,
            I => \N__14190\
        );

    \I__1734\ : InMux
    port map (
            O => \N__14197\,
            I => \N__14185\
        );

    \I__1733\ : InMux
    port map (
            O => \N__14196\,
            I => \N__14185\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__14193\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__14190\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__14185\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1729\ : InMux
    port map (
            O => \N__14178\,
            I => \N__14172\
        );

    \I__1728\ : InMux
    port map (
            O => \N__14177\,
            I => \N__14172\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__14172\,
            I => \N__14169\
        );

    \I__1726\ : Span4Mux_h
    port map (
            O => \N__14169\,
            I => \N__14165\
        );

    \I__1725\ : InMux
    port map (
            O => \N__14168\,
            I => \N__14162\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__14165\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__14162\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1722\ : CEMux
    port map (
            O => \N__14157\,
            I => \N__14151\
        );

    \I__1721\ : CEMux
    port map (
            O => \N__14156\,
            I => \N__14147\
        );

    \I__1720\ : CEMux
    port map (
            O => \N__14155\,
            I => \N__14144\
        );

    \I__1719\ : CEMux
    port map (
            O => \N__14154\,
            I => \N__14141\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__14151\,
            I => \N__14138\
        );

    \I__1717\ : CEMux
    port map (
            O => \N__14150\,
            I => \N__14135\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__14147\,
            I => \N__14132\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__14144\,
            I => \N__14129\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__14141\,
            I => \N__14122\
        );

    \I__1713\ : Span4Mux_h
    port map (
            O => \N__14138\,
            I => \N__14122\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__14135\,
            I => \N__14122\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__14132\,
            I => \N__14119\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__14129\,
            I => \N__14114\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__14122\,
            I => \N__14114\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__14119\,
            I => \this_vga_signals.N_966_0\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__14114\,
            I => \this_vga_signals.N_966_0\
        );

    \I__1706\ : SRMux
    port map (
            O => \N__14109\,
            I => \N__14091\
        );

    \I__1705\ : SRMux
    port map (
            O => \N__14108\,
            I => \N__14091\
        );

    \I__1704\ : SRMux
    port map (
            O => \N__14107\,
            I => \N__14091\
        );

    \I__1703\ : SRMux
    port map (
            O => \N__14106\,
            I => \N__14091\
        );

    \I__1702\ : SRMux
    port map (
            O => \N__14105\,
            I => \N__14091\
        );

    \I__1701\ : SRMux
    port map (
            O => \N__14104\,
            I => \N__14091\
        );

    \I__1700\ : GlobalMux
    port map (
            O => \N__14091\,
            I => \N__14088\
        );

    \I__1699\ : gio2CtrlBuf
    port map (
            O => \N__14088\,
            I => \this_vga_signals.N_1332_g\
        );

    \I__1698\ : InMux
    port map (
            O => \N__14085\,
            I => \N__14082\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__14082\,
            I => \N__14079\
        );

    \I__1696\ : Span4Mux_h
    port map (
            O => \N__14079\,
            I => \N__14076\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__14076\,
            I => \this_vga_signals.g1_0_0_0_0\
        );

    \I__1694\ : InMux
    port map (
            O => \N__14073\,
            I => \N__14070\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__14070\,
            I => \N__14067\
        );

    \I__1692\ : Span4Mux_h
    port map (
            O => \N__14067\,
            I => \N__14064\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__14064\,
            I => \this_vga_signals.g0_2_2_1\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__14061\,
            I => \this_vga_signals.N_473_0_cascade_\
        );

    \I__1689\ : InMux
    port map (
            O => \N__14058\,
            I => \N__14055\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__14055\,
            I => \this_vga_signals.N_554\
        );

    \I__1687\ : InMux
    port map (
            O => \N__14052\,
            I => \N__14048\
        );

    \I__1686\ : InMux
    port map (
            O => \N__14051\,
            I => \N__14045\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__14048\,
            I => \this_vga_signals.SUM_3_i_1_0\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__14045\,
            I => \this_vga_signals.SUM_3_i_1_0\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__14040\,
            I => \this_vga_signals.N_735_0_cascade_\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__14037\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_2_cascade_\
        );

    \I__1681\ : InMux
    port map (
            O => \N__14034\,
            I => \N__14027\
        );

    \I__1680\ : InMux
    port map (
            O => \N__14033\,
            I => \N__14027\
        );

    \I__1679\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14024\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__14027\,
            I => \this_vga_signals.N_735_0\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__14024\,
            I => \this_vga_signals.N_735_0\
        );

    \I__1676\ : InMux
    port map (
            O => \N__14019\,
            I => \N__14016\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__14016\,
            I => \N__14012\
        );

    \I__1674\ : InMux
    port map (
            O => \N__14015\,
            I => \N__14009\
        );

    \I__1673\ : Span4Mux_h
    port map (
            O => \N__14012\,
            I => \N__14003\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__14009\,
            I => \N__14000\
        );

    \I__1671\ : InMux
    port map (
            O => \N__14008\,
            I => \N__13997\
        );

    \I__1670\ : InMux
    port map (
            O => \N__14007\,
            I => \N__13992\
        );

    \I__1669\ : InMux
    port map (
            O => \N__14006\,
            I => \N__13992\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__14003\,
            I => \this_vga_signals.mult1_un61_sum_0_3\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__14000\,
            I => \this_vga_signals.mult1_un61_sum_0_3\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__13997\,
            I => \this_vga_signals.mult1_un61_sum_0_3\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__13992\,
            I => \this_vga_signals.mult1_un61_sum_0_3\
        );

    \I__1664\ : InMux
    port map (
            O => \N__13983\,
            I => \N__13980\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__13980\,
            I => \this_vga_signals.hsync_1_i_0_1\
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__13977\,
            I => \N__13974\
        );

    \I__1661\ : InMux
    port map (
            O => \N__13974\,
            I => \N__13971\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__13971\,
            I => \this_vga_signals.N_507_0\
        );

    \I__1659\ : InMux
    port map (
            O => \N__13968\,
            I => \N__13965\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__13965\,
            I => \N__13962\
        );

    \I__1657\ : Odrv12
    port map (
            O => \N__13962\,
            I => \M_this_map_ram_write_data_6\
        );

    \I__1656\ : InMux
    port map (
            O => \N__13959\,
            I => \N__13956\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__13956\,
            I => \N__13953\
        );

    \I__1654\ : Span4Mux_v
    port map (
            O => \N__13953\,
            I => \N__13948\
        );

    \I__1653\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13943\
        );

    \I__1652\ : InMux
    port map (
            O => \N__13951\,
            I => \N__13943\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__13948\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__13943\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__13938\,
            I => \N__13935\
        );

    \I__1648\ : InMux
    port map (
            O => \N__13935\,
            I => \N__13932\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__13932\,
            I => \N__13929\
        );

    \I__1646\ : Span4Mux_v
    port map (
            O => \N__13929\,
            I => \N__13926\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__13926\,
            I => \this_vga_signals.M_lcounter_d_0_sqmuxa\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__13923\,
            I => \N__13918\
        );

    \I__1643\ : InMux
    port map (
            O => \N__13922\,
            I => \N__13915\
        );

    \I__1642\ : InMux
    port map (
            O => \N__13921\,
            I => \N__13912\
        );

    \I__1641\ : InMux
    port map (
            O => \N__13918\,
            I => \N__13909\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__13915\,
            I => \N__13905\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__13912\,
            I => \N__13900\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__13909\,
            I => \N__13900\
        );

    \I__1637\ : InMux
    port map (
            O => \N__13908\,
            I => \N__13893\
        );

    \I__1636\ : Span4Mux_v
    port map (
            O => \N__13905\,
            I => \N__13890\
        );

    \I__1635\ : Span4Mux_v
    port map (
            O => \N__13900\,
            I => \N__13887\
        );

    \I__1634\ : InMux
    port map (
            O => \N__13899\,
            I => \N__13880\
        );

    \I__1633\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13880\
        );

    \I__1632\ : InMux
    port map (
            O => \N__13897\,
            I => \N__13880\
        );

    \I__1631\ : InMux
    port map (
            O => \N__13896\,
            I => \N__13877\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__13893\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__13890\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__13887\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__13880\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__13877\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__1625\ : InMux
    port map (
            O => \N__13866\,
            I => \N__13860\
        );

    \I__1624\ : InMux
    port map (
            O => \N__13865\,
            I => \N__13860\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__13860\,
            I => \N__13856\
        );

    \I__1622\ : InMux
    port map (
            O => \N__13859\,
            I => \N__13853\
        );

    \I__1621\ : Span4Mux_v
    port map (
            O => \N__13856\,
            I => \N__13850\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__13853\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__13850\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__13845\,
            I => \this_vga_signals.SUM_3_i_1_0_cascade_\
        );

    \I__1617\ : InMux
    port map (
            O => \N__13842\,
            I => \N__13839\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__13839\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_1\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__13836\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_1_cascade_\
        );

    \I__1614\ : InMux
    port map (
            O => \N__13833\,
            I => \N__13830\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__13830\,
            I => \this_vga_signals.if_N_8_i_0\
        );

    \I__1612\ : InMux
    port map (
            O => \N__13827\,
            I => \N__13824\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__13824\,
            I => \N__13821\
        );

    \I__1610\ : Odrv4
    port map (
            O => \N__13821\,
            I => \this_vga_signals.M_hcounter_d7lto7_0\
        );

    \I__1609\ : InMux
    port map (
            O => \N__13818\,
            I => \N__13815\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__13815\,
            I => \N__13812\
        );

    \I__1607\ : Span4Mux_h
    port map (
            O => \N__13812\,
            I => \N__13807\
        );

    \I__1606\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13804\
        );

    \I__1605\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13801\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__13807\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__13804\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__13801\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__13794\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\
        );

    \I__1600\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13788\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__13788\,
            I => \this_vga_signals.mult1_un61_sum_axbxc1\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__13785\,
            I => \this_vga_signals.mult1_un61_sum_axbxc1_cascade_\
        );

    \I__1597\ : InMux
    port map (
            O => \N__13782\,
            I => \N__13779\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__13779\,
            I => \N__13775\
        );

    \I__1595\ : InMux
    port map (
            O => \N__13778\,
            I => \N__13772\
        );

    \I__1594\ : Span4Mux_h
    port map (
            O => \N__13775\,
            I => \N__13765\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__13772\,
            I => \N__13762\
        );

    \I__1592\ : InMux
    port map (
            O => \N__13771\,
            I => \N__13757\
        );

    \I__1591\ : InMux
    port map (
            O => \N__13770\,
            I => \N__13757\
        );

    \I__1590\ : InMux
    port map (
            O => \N__13769\,
            I => \N__13752\
        );

    \I__1589\ : InMux
    port map (
            O => \N__13768\,
            I => \N__13752\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__13765\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__13762\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__13757\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__13752\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__1584\ : IoInMux
    port map (
            O => \N__13743\,
            I => \N__13740\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__13740\,
            I => \N__13737\
        );

    \I__1582\ : Span12Mux_s11_v
    port map (
            O => \N__13737\,
            I => \N__13734\
        );

    \I__1581\ : Span12Mux_h
    port map (
            O => \N__13734\,
            I => \N__13731\
        );

    \I__1580\ : Odrv12
    port map (
            O => \N__13731\,
            I => \M_hcounter_q_esr_RNIR18F4_9\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__13728\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0_1_1_cascade_\
        );

    \I__1578\ : InMux
    port map (
            O => \N__13725\,
            I => \N__13719\
        );

    \I__1577\ : InMux
    port map (
            O => \N__13724\,
            I => \N__13719\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__13719\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_1\
        );

    \I__1575\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13713\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__13713\,
            I => \this_vga_signals.mult1_un89_sum_c3\
        );

    \I__1573\ : InMux
    port map (
            O => \N__13710\,
            I => \N__13707\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__13707\,
            I => \this_vga_signals.mult1_un75_sum_c2_0\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__13704\,
            I => \this_vga_signals.mult1_un75_sum_c2_0_cascade_\
        );

    \I__1570\ : InMux
    port map (
            O => \N__13701\,
            I => \N__13698\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__13698\,
            I => \this_vga_signals.if_N_9_1\
        );

    \I__1568\ : InMux
    port map (
            O => \N__13695\,
            I => \N__13690\
        );

    \I__1567\ : InMux
    port map (
            O => \N__13694\,
            I => \N__13685\
        );

    \I__1566\ : InMux
    port map (
            O => \N__13693\,
            I => \N__13685\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__13690\,
            I => \this_vga_signals.if_m7_0_x4_0\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__13685\,
            I => \this_vga_signals.if_m7_0_x4_0\
        );

    \I__1563\ : InMux
    port map (
            O => \N__13680\,
            I => \N__13676\
        );

    \I__1562\ : InMux
    port map (
            O => \N__13679\,
            I => \N__13673\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__13676\,
            I => \this_vga_signals.mult1_un75_sum_c3\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__13673\,
            I => \this_vga_signals.mult1_un75_sum_c3\
        );

    \I__1559\ : InMux
    port map (
            O => \N__13668\,
            I => \N__13661\
        );

    \I__1558\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13658\
        );

    \I__1557\ : InMux
    port map (
            O => \N__13666\,
            I => \N__13651\
        );

    \I__1556\ : InMux
    port map (
            O => \N__13665\,
            I => \N__13651\
        );

    \I__1555\ : InMux
    port map (
            O => \N__13664\,
            I => \N__13651\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__13661\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_2\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__13658\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_2\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__13651\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_2\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__13644\,
            I => \this_vga_signals.mult1_un75_sum_c3_cascade_\
        );

    \I__1550\ : InMux
    port map (
            O => \N__13641\,
            I => \N__13637\
        );

    \I__1549\ : InMux
    port map (
            O => \N__13640\,
            I => \N__13634\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__13637\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_0\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__13634\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_0\
        );

    \I__1546\ : InMux
    port map (
            O => \N__13629\,
            I => \N__13623\
        );

    \I__1545\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13620\
        );

    \I__1544\ : InMux
    port map (
            O => \N__13627\,
            I => \N__13615\
        );

    \I__1543\ : InMux
    port map (
            O => \N__13626\,
            I => \N__13615\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__13623\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__13620\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__13615\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1539\ : InMux
    port map (
            O => \N__13608\,
            I => \N__13603\
        );

    \I__1538\ : InMux
    port map (
            O => \N__13607\,
            I => \N__13600\
        );

    \I__1537\ : InMux
    port map (
            O => \N__13606\,
            I => \N__13597\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__13603\,
            I => \this_vga_signals.N_3_0\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__13600\,
            I => \this_vga_signals.N_3_0\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__13597\,
            I => \this_vga_signals.N_3_0\
        );

    \I__1533\ : InMux
    port map (
            O => \N__13590\,
            I => \N__13580\
        );

    \I__1532\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13580\
        );

    \I__1531\ : InMux
    port map (
            O => \N__13588\,
            I => \N__13580\
        );

    \I__1530\ : InMux
    port map (
            O => \N__13587\,
            I => \N__13577\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__13580\,
            I => \this_vga_signals.M_pcounter_q_i_3_1\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__13577\,
            I => \this_vga_signals.M_pcounter_q_i_3_1\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__13572\,
            I => \this_vga_signals.M_lcounter_d_0_sqmuxa_cascade_\
        );

    \I__1526\ : InMux
    port map (
            O => \N__13569\,
            I => \N__13565\
        );

    \I__1525\ : InMux
    port map (
            O => \N__13568\,
            I => \N__13562\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__13565\,
            I => \this_vga_signals.N_2_0\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__13562\,
            I => \this_vga_signals.N_2_0\
        );

    \I__1522\ : InMux
    port map (
            O => \N__13557\,
            I => \N__13553\
        );

    \I__1521\ : InMux
    port map (
            O => \N__13556\,
            I => \N__13550\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__13553\,
            I => \this_vga_signals.M_pcounter_q_i_3_0\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__13550\,
            I => \this_vga_signals.M_pcounter_q_i_3_0\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__13545\,
            I => \this_vga_signals.M_hcounter_d7lt7_0_cascade_\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__13542\,
            I => \this_vga_signals.M_hcounter_d7_0_cascade_\
        );

    \I__1516\ : InMux
    port map (
            O => \N__13539\,
            I => \N__13536\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__13536\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__13533\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0_x0_cascade_\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__13530\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0_cascade_\
        );

    \I__1512\ : InMux
    port map (
            O => \N__13527\,
            I => \N__13524\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__13524\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__13521\,
            I => \this_vga_signals.g1_5_cascade_\
        );

    \I__1509\ : InMux
    port map (
            O => \N__13518\,
            I => \N__13515\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__13515\,
            I => \this_vga_signals.g1_0_0\
        );

    \I__1507\ : InMux
    port map (
            O => \N__13512\,
            I => \N__13509\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__13509\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0_x1\
        );

    \I__1505\ : InMux
    port map (
            O => \N__13506\,
            I => \N__13503\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__13503\,
            I => \this_vga_signals.g1_2\
        );

    \I__1503\ : InMux
    port map (
            O => \N__13500\,
            I => \N__13489\
        );

    \I__1502\ : InMux
    port map (
            O => \N__13499\,
            I => \N__13489\
        );

    \I__1501\ : InMux
    port map (
            O => \N__13498\,
            I => \N__13486\
        );

    \I__1500\ : InMux
    port map (
            O => \N__13497\,
            I => \N__13483\
        );

    \I__1499\ : InMux
    port map (
            O => \N__13496\,
            I => \N__13478\
        );

    \I__1498\ : InMux
    port map (
            O => \N__13495\,
            I => \N__13478\
        );

    \I__1497\ : InMux
    port map (
            O => \N__13494\,
            I => \N__13475\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__13489\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_ns\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__13486\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_ns\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__13483\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_ns\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__13478\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_ns\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__13475\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_ns\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__13464\,
            I => \this_vga_signals.mult1_un68_sum_axb1_cascade_\
        );

    \I__1490\ : InMux
    port map (
            O => \N__13461\,
            I => \N__13458\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__13458\,
            I => \this_vga_signals.mult1_un68_sum_c2_0\
        );

    \I__1488\ : CascadeMux
    port map (
            O => \N__13455\,
            I => \this_vga_signals.mult1_un54_sum_axb1_cascade_\
        );

    \I__1487\ : InMux
    port map (
            O => \N__13452\,
            I => \N__13449\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__13449\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x0\
        );

    \I__1485\ : InMux
    port map (
            O => \N__13446\,
            I => \N__13442\
        );

    \I__1484\ : InMux
    port map (
            O => \N__13445\,
            I => \N__13439\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__13442\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_0_0\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__13439\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_0_0\
        );

    \I__1481\ : InMux
    port map (
            O => \N__13434\,
            I => \N__13430\
        );

    \I__1480\ : InMux
    port map (
            O => \N__13433\,
            I => \N__13427\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__13430\,
            I => \this_vga_signals.if_i2_mux\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__13427\,
            I => \this_vga_signals.if_i2_mux\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__13422\,
            I => \this_vga_signals.g0_1_1_x0_cascade_\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__13419\,
            I => \this_vga_signals.g0_1_1_cascade_\
        );

    \I__1475\ : InMux
    port map (
            O => \N__13416\,
            I => \N__13413\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__13413\,
            I => \this_vga_signals.N_4_0_0_0\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__13410\,
            I => \this_vga_signals.g0_0_0_0_0_cascade_\
        );

    \I__1472\ : InMux
    port map (
            O => \N__13407\,
            I => \N__13398\
        );

    \I__1471\ : InMux
    port map (
            O => \N__13406\,
            I => \N__13398\
        );

    \I__1470\ : InMux
    port map (
            O => \N__13405\,
            I => \N__13393\
        );

    \I__1469\ : InMux
    port map (
            O => \N__13404\,
            I => \N__13393\
        );

    \I__1468\ : InMux
    port map (
            O => \N__13403\,
            I => \N__13390\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__13398\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__13393\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__13390\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1464\ : InMux
    port map (
            O => \N__13383\,
            I => \N__13375\
        );

    \I__1463\ : InMux
    port map (
            O => \N__13382\,
            I => \N__13375\
        );

    \I__1462\ : InMux
    port map (
            O => \N__13381\,
            I => \N__13370\
        );

    \I__1461\ : InMux
    port map (
            O => \N__13380\,
            I => \N__13370\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__13375\,
            I => \N__13367\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__13370\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1458\ : Odrv4
    port map (
            O => \N__13367\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__13362\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_\
        );

    \I__1456\ : InMux
    port map (
            O => \N__13359\,
            I => \N__13356\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__13356\,
            I => \N__13351\
        );

    \I__1454\ : InMux
    port map (
            O => \N__13355\,
            I => \N__13346\
        );

    \I__1453\ : InMux
    port map (
            O => \N__13354\,
            I => \N__13346\
        );

    \I__1452\ : Span4Mux_v
    port map (
            O => \N__13351\,
            I => \N__13343\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__13346\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__13343\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__13338\,
            I => \N__13335\
        );

    \I__1448\ : InMux
    port map (
            O => \N__13335\,
            I => \N__13332\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__13332\,
            I => \N__13329\
        );

    \I__1446\ : Odrv4
    port map (
            O => \N__13329\,
            I => \this_vga_signals.g0_0_0_1\
        );

    \I__1445\ : InMux
    port map (
            O => \N__13326\,
            I => \N__13323\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__13323\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i_0\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__13320\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_cascade_\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__13317\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_cascade_\
        );

    \I__1441\ : InMux
    port map (
            O => \N__13314\,
            I => \N__13311\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__13311\,
            I => \N__13308\
        );

    \I__1439\ : Odrv12
    port map (
            O => \N__13308\,
            I => \M_this_map_ram_write_data_0\
        );

    \I__1438\ : InMux
    port map (
            O => \N__13305\,
            I => \N__13302\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__13302\,
            I => \N__13299\
        );

    \I__1436\ : Span4Mux_h
    port map (
            O => \N__13299\,
            I => \N__13296\
        );

    \I__1435\ : Span4Mux_h
    port map (
            O => \N__13296\,
            I => \N__13293\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__13293\,
            I => \M_this_map_ram_write_data_7\
        );

    \I__1433\ : InMux
    port map (
            O => \N__13290\,
            I => \N__13287\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__13287\,
            I => \N__13284\
        );

    \I__1431\ : Span4Mux_v
    port map (
            O => \N__13284\,
            I => \N__13281\
        );

    \I__1430\ : Odrv4
    port map (
            O => \N__13281\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__1429\ : InMux
    port map (
            O => \N__13278\,
            I => \N__13275\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__13275\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__13272\,
            I => \this_vga_signals.N_1_4_1_cascade_\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__13269\,
            I => \this_vga_signals.SUM_2_i_1_2_3_cascade_\
        );

    \I__1425\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13263\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__13263\,
            I => \N__13255\
        );

    \I__1423\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13250\
        );

    \I__1422\ : InMux
    port map (
            O => \N__13261\,
            I => \N__13250\
        );

    \I__1421\ : InMux
    port map (
            O => \N__13260\,
            I => \N__13243\
        );

    \I__1420\ : InMux
    port map (
            O => \N__13259\,
            I => \N__13243\
        );

    \I__1419\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13243\
        );

    \I__1418\ : Odrv4
    port map (
            O => \N__13255\,
            I => \N_880_0\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__13250\,
            I => \N_880_0\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__13243\,
            I => \N_880_0\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__13236\,
            I => \N__13233\
        );

    \I__1414\ : InMux
    port map (
            O => \N__13233\,
            I => \N__13230\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__13230\,
            I => \N__13227\
        );

    \I__1412\ : Span4Mux_h
    port map (
            O => \N__13227\,
            I => \N__13224\
        );

    \I__1411\ : Span4Mux_h
    port map (
            O => \N__13224\,
            I => \N__13221\
        );

    \I__1410\ : Odrv4
    port map (
            O => \N__13221\,
            I => \M_this_vga_signals_address_2\
        );

    \I__1409\ : InMux
    port map (
            O => \N__13218\,
            I => \N__13215\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__13215\,
            I => \this_vga_signals.mult1_un82_sum_c2_0\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__13212\,
            I => \this_vga_signals.mult1_un82_sum_c2_0_cascade_\
        );

    \I__1406\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13203\
        );

    \I__1405\ : InMux
    port map (
            O => \N__13208\,
            I => \N__13203\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__13203\,
            I => \this_vga_signals.mult1_un82_sum_c3_0\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__13200\,
            I => \N__13197\
        );

    \I__1402\ : InMux
    port map (
            O => \N__13197\,
            I => \N__13193\
        );

    \I__1401\ : InMux
    port map (
            O => \N__13196\,
            I => \N__13190\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__13193\,
            I => \this_vga_signals.mult1_un75_sum_axbxc1\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__13190\,
            I => \this_vga_signals.mult1_un75_sum_axbxc1\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__13185\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_2_0_cascade_\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__13182\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_2_cascade_\
        );

    \I__1396\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13175\
        );

    \I__1395\ : InMux
    port map (
            O => \N__13178\,
            I => \N__13172\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__13175\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__13172\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1\
        );

    \I__1392\ : InMux
    port map (
            O => \N__13167\,
            I => \N__13164\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__13164\,
            I => \N__13161\
        );

    \I__1390\ : Span12Mux_v
    port map (
            O => \N__13161\,
            I => \N__13158\
        );

    \I__1389\ : Span12Mux_v
    port map (
            O => \N__13158\,
            I => \N__13155\
        );

    \I__1388\ : Span12Mux_h
    port map (
            O => \N__13155\,
            I => \N__13152\
        );

    \I__1387\ : Odrv12
    port map (
            O => \N__13152\,
            I => \M_this_oam_ram_read_data_4\
        );

    \I__1386\ : InMux
    port map (
            O => \N__13149\,
            I => \N__13146\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__13146\,
            I => \N__13143\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__13143\,
            I => \N__13140\
        );

    \I__1383\ : Span4Mux_v
    port map (
            O => \N__13140\,
            I => \N__13137\
        );

    \I__1382\ : Span4Mux_h
    port map (
            O => \N__13137\,
            I => \N__13134\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__13134\,
            I => \M_this_map_ram_read_data_4\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__13131\,
            I => \N__13128\
        );

    \I__1379\ : InMux
    port map (
            O => \N__13128\,
            I => \N__13122\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__13127\,
            I => \N__13119\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__13126\,
            I => \N__13114\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__13125\,
            I => \N__13108\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__13122\,
            I => \N__13102\
        );

    \I__1374\ : InMux
    port map (
            O => \N__13119\,
            I => \N__13099\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__13118\,
            I => \N__13096\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__13117\,
            I => \N__13093\
        );

    \I__1371\ : InMux
    port map (
            O => \N__13114\,
            I => \N__13090\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__13113\,
            I => \N__13087\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__13112\,
            I => \N__13083\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__13111\,
            I => \N__13078\
        );

    \I__1367\ : InMux
    port map (
            O => \N__13108\,
            I => \N__13075\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__13107\,
            I => \N__13072\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__13106\,
            I => \N__13069\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__13105\,
            I => \N__13066\
        );

    \I__1363\ : Span4Mux_s3_v
    port map (
            O => \N__13102\,
            I => \N__13061\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__13099\,
            I => \N__13061\
        );

    \I__1361\ : InMux
    port map (
            O => \N__13096\,
            I => \N__13058\
        );

    \I__1360\ : InMux
    port map (
            O => \N__13093\,
            I => \N__13055\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__13090\,
            I => \N__13052\
        );

    \I__1358\ : InMux
    port map (
            O => \N__13087\,
            I => \N__13049\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__13086\,
            I => \N__13046\
        );

    \I__1356\ : InMux
    port map (
            O => \N__13083\,
            I => \N__13043\
        );

    \I__1355\ : CascadeMux
    port map (
            O => \N__13082\,
            I => \N__13040\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__13081\,
            I => \N__13037\
        );

    \I__1353\ : InMux
    port map (
            O => \N__13078\,
            I => \N__13033\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__13075\,
            I => \N__13030\
        );

    \I__1351\ : InMux
    port map (
            O => \N__13072\,
            I => \N__13027\
        );

    \I__1350\ : InMux
    port map (
            O => \N__13069\,
            I => \N__13024\
        );

    \I__1349\ : InMux
    port map (
            O => \N__13066\,
            I => \N__13021\
        );

    \I__1348\ : Span4Mux_v
    port map (
            O => \N__13061\,
            I => \N__13014\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__13058\,
            I => \N__13014\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__13055\,
            I => \N__13014\
        );

    \I__1345\ : Span4Mux_h
    port map (
            O => \N__13052\,
            I => \N__13009\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__13049\,
            I => \N__13009\
        );

    \I__1343\ : InMux
    port map (
            O => \N__13046\,
            I => \N__13006\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__13043\,
            I => \N__13003\
        );

    \I__1341\ : InMux
    port map (
            O => \N__13040\,
            I => \N__13000\
        );

    \I__1340\ : InMux
    port map (
            O => \N__13037\,
            I => \N__12997\
        );

    \I__1339\ : CascadeMux
    port map (
            O => \N__13036\,
            I => \N__12994\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__13033\,
            I => \N__12991\
        );

    \I__1337\ : Span4Mux_v
    port map (
            O => \N__13030\,
            I => \N__12988\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__13027\,
            I => \N__12985\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__13024\,
            I => \N__12982\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__13021\,
            I => \N__12979\
        );

    \I__1333\ : Span4Mux_v
    port map (
            O => \N__13014\,
            I => \N__12972\
        );

    \I__1332\ : Span4Mux_v
    port map (
            O => \N__13009\,
            I => \N__12972\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__13006\,
            I => \N__12972\
        );

    \I__1330\ : Span4Mux_v
    port map (
            O => \N__13003\,
            I => \N__12967\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__13000\,
            I => \N__12967\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__12997\,
            I => \N__12964\
        );

    \I__1327\ : InMux
    port map (
            O => \N__12994\,
            I => \N__12961\
        );

    \I__1326\ : Span12Mux_h
    port map (
            O => \N__12991\,
            I => \N__12958\
        );

    \I__1325\ : Sp12to4
    port map (
            O => \N__12988\,
            I => \N__12953\
        );

    \I__1324\ : Span12Mux_v
    port map (
            O => \N__12985\,
            I => \N__12953\
        );

    \I__1323\ : Span12Mux_s6_v
    port map (
            O => \N__12982\,
            I => \N__12948\
        );

    \I__1322\ : Span12Mux_v
    port map (
            O => \N__12979\,
            I => \N__12948\
        );

    \I__1321\ : Span4Mux_h
    port map (
            O => \N__12972\,
            I => \N__12945\
        );

    \I__1320\ : Span4Mux_v
    port map (
            O => \N__12967\,
            I => \N__12940\
        );

    \I__1319\ : Span4Mux_h
    port map (
            O => \N__12964\,
            I => \N__12940\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__12961\,
            I => \N__12937\
        );

    \I__1317\ : Span12Mux_v
    port map (
            O => \N__12958\,
            I => \N__12934\
        );

    \I__1316\ : Span12Mux_h
    port map (
            O => \N__12953\,
            I => \N__12929\
        );

    \I__1315\ : Span12Mux_h
    port map (
            O => \N__12948\,
            I => \N__12929\
        );

    \I__1314\ : Sp12to4
    port map (
            O => \N__12945\,
            I => \N__12926\
        );

    \I__1313\ : Span4Mux_h
    port map (
            O => \N__12940\,
            I => \N__12923\
        );

    \I__1312\ : Span4Mux_h
    port map (
            O => \N__12937\,
            I => \N__12920\
        );

    \I__1311\ : Odrv12
    port map (
            O => \N__12934\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__1310\ : Odrv12
    port map (
            O => \N__12929\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__1309\ : Odrv12
    port map (
            O => \N__12926\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__12923\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__1307\ : Odrv4
    port map (
            O => \N__12920\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__12909\,
            I => \this_vga_signals.M_vcounter_d7lt3_cascade_\
        );

    \I__1305\ : InMux
    port map (
            O => \N__12906\,
            I => \N__12903\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__12903\,
            I => \this_vga_ramdac.N_24_mux\
        );

    \I__1303\ : InMux
    port map (
            O => \N__12900\,
            I => \N__12897\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__12897\,
            I => \N__12888\
        );

    \I__1301\ : InMux
    port map (
            O => \N__12896\,
            I => \N__12885\
        );

    \I__1300\ : InMux
    port map (
            O => \N__12895\,
            I => \N__12880\
        );

    \I__1299\ : InMux
    port map (
            O => \N__12894\,
            I => \N__12880\
        );

    \I__1298\ : InMux
    port map (
            O => \N__12893\,
            I => \N__12877\
        );

    \I__1297\ : InMux
    port map (
            O => \N__12892\,
            I => \N__12872\
        );

    \I__1296\ : InMux
    port map (
            O => \N__12891\,
            I => \N__12872\
        );

    \I__1295\ : Odrv4
    port map (
            O => \N__12888\,
            I => \M_pcounter_q_ret_2_RNIH7PG8\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__12885\,
            I => \M_pcounter_q_ret_2_RNIH7PG8\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__12880\,
            I => \M_pcounter_q_ret_2_RNIH7PG8\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__12877\,
            I => \M_pcounter_q_ret_2_RNIH7PG8\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__12872\,
            I => \M_pcounter_q_ret_2_RNIH7PG8\
        );

    \I__1290\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12857\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__12860\,
            I => \N__12854\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__12857\,
            I => \N__12851\
        );

    \I__1287\ : InMux
    port map (
            O => \N__12854\,
            I => \N__12848\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__12851\,
            I => \this_vga_ramdac.N_3298_reto\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__12848\,
            I => \this_vga_ramdac.N_3298_reto\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__12843\,
            I => \this_vga_signals.M_pcounter_q_3_1_cascade_\
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__12840\,
            I => \N__12836\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__12839\,
            I => \N__12832\
        );

    \I__1281\ : InMux
    port map (
            O => \N__12836\,
            I => \N__12825\
        );

    \I__1280\ : InMux
    port map (
            O => \N__12835\,
            I => \N__12825\
        );

    \I__1279\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12825\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__12825\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__1277\ : InMux
    port map (
            O => \N__12822\,
            I => \N__12817\
        );

    \I__1276\ : InMux
    port map (
            O => \N__12821\,
            I => \N__12812\
        );

    \I__1275\ : InMux
    port map (
            O => \N__12820\,
            I => \N__12812\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__12817\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__12812\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__12807\,
            I => \N__12804\
        );

    \I__1271\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12801\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__12801\,
            I => \N__12798\
        );

    \I__1269\ : Span4Mux_h
    port map (
            O => \N__12798\,
            I => \N__12795\
        );

    \I__1268\ : Span4Mux_h
    port map (
            O => \N__12795\,
            I => \N__12792\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__12792\,
            I => \M_this_vga_signals_address_1\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__12789\,
            I => \this_vga_signals.mult1_un89_sum_axbxc3_1_cascade_\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__12786\,
            I => \N__12783\
        );

    \I__1264\ : InMux
    port map (
            O => \N__12783\,
            I => \N__12780\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__12780\,
            I => \N__12777\
        );

    \I__1262\ : Span12Mux_h
    port map (
            O => \N__12777\,
            I => \N__12774\
        );

    \I__1261\ : Odrv12
    port map (
            O => \N__12774\,
            I => \M_this_vga_signals_address_0\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__12771\,
            I => \this_vga_signals.g0_2_1_cascade_\
        );

    \I__1259\ : InMux
    port map (
            O => \N__12768\,
            I => \N__12765\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__12765\,
            I => \this_vga_signals.N_5_0_0\
        );

    \I__1257\ : InMux
    port map (
            O => \N__12762\,
            I => \N__12759\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__12759\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_x1\
        );

    \I__1255\ : InMux
    port map (
            O => \N__12756\,
            I => \N__12753\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__12753\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_x0\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__12750\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_ns_cascade_\
        );

    \I__1252\ : InMux
    port map (
            O => \N__12747\,
            I => \N__12744\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__12744\,
            I => \this_vga_signals.g0_31_N_4L6\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__12741\,
            I => \this_vga_signals.g0_31_N_2L1_cascade_\
        );

    \I__1249\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12735\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__12735\,
            I => \this_vga_signals.g0_31_N_5L8\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__12732\,
            I => \this_vga_signals.M_pcounter_q_3_0_cascade_\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__12729\,
            I => \this_vga_signals.N_2_0_cascade_\
        );

    \I__1245\ : InMux
    port map (
            O => \N__12726\,
            I => \N__12723\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__12723\,
            I => \this_vga_signals.M_this_vga_signals_pixel_clk_0_0\
        );

    \I__1243\ : InMux
    port map (
            O => \N__12720\,
            I => \N__12715\
        );

    \I__1242\ : InMux
    port map (
            O => \N__12719\,
            I => \N__12712\
        );

    \I__1241\ : InMux
    port map (
            O => \N__12718\,
            I => \N__12709\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__12715\,
            I => \N__12704\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__12712\,
            I => \N__12704\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__12709\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1237\ : Odrv12
    port map (
            O => \N__12704\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__12699\,
            I => \this_vga_signals.if_i1_mux_0_cascade_\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__12696\,
            I => \N__12693\
        );

    \I__1234\ : InMux
    port map (
            O => \N__12693\,
            I => \N__12690\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__12690\,
            I => \N__12687\
        );

    \I__1232\ : Span4Mux_h
    port map (
            O => \N__12687\,
            I => \N__12684\
        );

    \I__1231\ : Span4Mux_h
    port map (
            O => \N__12684\,
            I => \N__12681\
        );

    \I__1230\ : Odrv4
    port map (
            O => \N__12681\,
            I => \M_this_vga_signals_address_7\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__12678\,
            I => \this_vga_signals.N_5_i_0_cascade_\
        );

    \I__1228\ : InMux
    port map (
            O => \N__12675\,
            I => \N__12672\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__12672\,
            I => \this_vga_signals.mult1_un82_sum_c3\
        );

    \I__1226\ : InMux
    port map (
            O => \N__12669\,
            I => \N__12666\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__12666\,
            I => \this_vga_signals.N_3_2_0_1\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__12663\,
            I => \this_vga_signals.g0_i_x4_0_0_cascade_\
        );

    \I__1223\ : InMux
    port map (
            O => \N__12660\,
            I => \N__12657\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__12657\,
            I => \this_vga_signals.N_3_3_0_0\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__12654\,
            I => \this_vga_signals.g0_0_2_0_0_cascade_\
        );

    \I__1220\ : InMux
    port map (
            O => \N__12651\,
            I => \N__12648\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__12648\,
            I => \this_vga_signals.g0_6_2\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__12645\,
            I => \this_vga_signals.g1_1_0_0_0_cascade_\
        );

    \I__1217\ : InMux
    port map (
            O => \N__12642\,
            I => \N__12639\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__12639\,
            I => \this_vga_signals.N_5_i_1_0_0\
        );

    \I__1215\ : InMux
    port map (
            O => \N__12636\,
            I => \N__12633\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__12633\,
            I => \N__12628\
        );

    \I__1213\ : InMux
    port map (
            O => \N__12632\,
            I => \N__12623\
        );

    \I__1212\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12623\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__12628\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__12623\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__1209\ : InMux
    port map (
            O => \N__12618\,
            I => \N__12615\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__12615\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__12612\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__12609\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__12606\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\
        );

    \I__1204\ : InMux
    port map (
            O => \N__12603\,
            I => \N__12600\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__12600\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_0\
        );

    \I__1202\ : InMux
    port map (
            O => \N__12597\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_1\
        );

    \I__1201\ : InMux
    port map (
            O => \N__12594\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_2\
        );

    \I__1200\ : InMux
    port map (
            O => \N__12591\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3\
        );

    \I__1199\ : InMux
    port map (
            O => \N__12588\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4\
        );

    \I__1198\ : InMux
    port map (
            O => \N__12585\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5\
        );

    \I__1197\ : InMux
    port map (
            O => \N__12582\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6\
        );

    \I__1196\ : InMux
    port map (
            O => \N__12579\,
            I => \bfn_13_13_0_\
        );

    \I__1195\ : InMux
    port map (
            O => \N__12576\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__12573\,
            I => \N_880_0_cascade_\
        );

    \I__1193\ : CascadeMux
    port map (
            O => \N__12570\,
            I => \N__12567\
        );

    \I__1192\ : InMux
    port map (
            O => \N__12567\,
            I => \N__12564\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__12564\,
            I => \N__12561\
        );

    \I__1190\ : Span4Mux_v
    port map (
            O => \N__12561\,
            I => \N__12558\
        );

    \I__1189\ : Odrv4
    port map (
            O => \N__12558\,
            I => \M_this_vga_signals_address_5\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__12555\,
            I => \N__12552\
        );

    \I__1187\ : InMux
    port map (
            O => \N__12552\,
            I => \N__12549\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__12549\,
            I => \N__12546\
        );

    \I__1185\ : Span4Mux_h
    port map (
            O => \N__12546\,
            I => \N__12543\
        );

    \I__1184\ : Odrv4
    port map (
            O => \N__12543\,
            I => \M_this_vga_signals_address_3\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__12540\,
            I => \N__12537\
        );

    \I__1182\ : InMux
    port map (
            O => \N__12537\,
            I => \N__12534\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__12534\,
            I => \N__12531\
        );

    \I__1180\ : Span4Mux_h
    port map (
            O => \N__12531\,
            I => \N__12528\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__12528\,
            I => \M_this_vga_signals_address_4\
        );

    \I__1178\ : InMux
    port map (
            O => \N__12525\,
            I => \N__12522\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__12522\,
            I => \N__12519\
        );

    \I__1176\ : Span12Mux_h
    port map (
            O => \N__12519\,
            I => \N__12516\
        );

    \I__1175\ : Odrv12
    port map (
            O => \N__12516\,
            I => port_clk_c
        );

    \I__1174\ : InMux
    port map (
            O => \N__12513\,
            I => \N__12510\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__12510\,
            I => \this_delay_clk.M_pipe_qZ0Z_0\
        );

    \I__1172\ : InMux
    port map (
            O => \N__12507\,
            I => \N__12504\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__12504\,
            I => \N__12501\
        );

    \I__1170\ : Span4Mux_h
    port map (
            O => \N__12501\,
            I => \N__12498\
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__12498\,
            I => \M_this_map_ram_write_data_1\
        );

    \I__1168\ : InMux
    port map (
            O => \N__12495\,
            I => \N__12492\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__12492\,
            I => \N__12489\
        );

    \I__1166\ : Span4Mux_h
    port map (
            O => \N__12489\,
            I => \N__12486\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__12486\,
            I => \M_this_map_ram_write_data_5\
        );

    \I__1164\ : InMux
    port map (
            O => \N__12483\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_0\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__12480\,
            I => \this_vga_ramdac.m19_cascade_\
        );

    \I__1162\ : InMux
    port map (
            O => \N__12477\,
            I => \N__12474\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__12474\,
            I => \N__12471\
        );

    \I__1160\ : Span4Mux_h
    port map (
            O => \N__12471\,
            I => \N__12468\
        );

    \I__1159\ : Sp12to4
    port map (
            O => \N__12468\,
            I => \N__12464\
        );

    \I__1158\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12461\
        );

    \I__1157\ : Odrv12
    port map (
            O => \N__12464\,
            I => \this_vga_ramdac.N_3302_reto\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__12461\,
            I => \this_vga_ramdac.N_3302_reto\
        );

    \I__1155\ : InMux
    port map (
            O => \N__12456\,
            I => \N__12453\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__12453\,
            I => \N__12449\
        );

    \I__1153\ : InMux
    port map (
            O => \N__12452\,
            I => \N__12446\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__12449\,
            I => \this_vga_ramdac.N_3303_reto\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__12446\,
            I => \this_vga_ramdac.N_3303_reto\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__12441\,
            I => \N__12437\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__12440\,
            I => \N__12434\
        );

    \I__1148\ : InMux
    port map (
            O => \N__12437\,
            I => \N__12425\
        );

    \I__1147\ : InMux
    port map (
            O => \N__12434\,
            I => \N__12425\
        );

    \I__1146\ : InMux
    port map (
            O => \N__12433\,
            I => \N__12416\
        );

    \I__1145\ : InMux
    port map (
            O => \N__12432\,
            I => \N__12416\
        );

    \I__1144\ : InMux
    port map (
            O => \N__12431\,
            I => \N__12416\
        );

    \I__1143\ : InMux
    port map (
            O => \N__12430\,
            I => \N__12416\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__12425\,
            I => \N__12411\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__12416\,
            I => \N__12411\
        );

    \I__1140\ : Span4Mux_h
    port map (
            O => \N__12411\,
            I => \N__12408\
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__12408\,
            I => \M_this_vram_read_data_0\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__12405\,
            I => \N__12400\
        );

    \I__1137\ : InMux
    port map (
            O => \N__12404\,
            I => \N__12392\
        );

    \I__1136\ : InMux
    port map (
            O => \N__12403\,
            I => \N__12392\
        );

    \I__1135\ : InMux
    port map (
            O => \N__12400\,
            I => \N__12383\
        );

    \I__1134\ : InMux
    port map (
            O => \N__12399\,
            I => \N__12383\
        );

    \I__1133\ : InMux
    port map (
            O => \N__12398\,
            I => \N__12383\
        );

    \I__1132\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12383\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__12392\,
            I => \N__12378\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__12383\,
            I => \N__12378\
        );

    \I__1129\ : Span4Mux_h
    port map (
            O => \N__12378\,
            I => \N__12375\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__12375\,
            I => \M_this_vram_read_data_3\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__12372\,
            I => \N__12365\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__12371\,
            I => \N__12362\
        );

    \I__1125\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12357\
        );

    \I__1124\ : InMux
    port map (
            O => \N__12369\,
            I => \N__12357\
        );

    \I__1123\ : InMux
    port map (
            O => \N__12368\,
            I => \N__12350\
        );

    \I__1122\ : InMux
    port map (
            O => \N__12365\,
            I => \N__12350\
        );

    \I__1121\ : InMux
    port map (
            O => \N__12362\,
            I => \N__12350\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__12357\,
            I => \N__12345\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__12350\,
            I => \N__12345\
        );

    \I__1118\ : Span4Mux_h
    port map (
            O => \N__12345\,
            I => \N__12342\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__12342\,
            I => \M_this_vram_read_data_2\
        );

    \I__1116\ : InMux
    port map (
            O => \N__12339\,
            I => \N__12329\
        );

    \I__1115\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12329\
        );

    \I__1114\ : InMux
    port map (
            O => \N__12337\,
            I => \N__12320\
        );

    \I__1113\ : InMux
    port map (
            O => \N__12336\,
            I => \N__12320\
        );

    \I__1112\ : InMux
    port map (
            O => \N__12335\,
            I => \N__12320\
        );

    \I__1111\ : InMux
    port map (
            O => \N__12334\,
            I => \N__12320\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__12329\,
            I => \N__12315\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__12320\,
            I => \N__12315\
        );

    \I__1108\ : Span4Mux_h
    port map (
            O => \N__12315\,
            I => \N__12312\
        );

    \I__1107\ : Odrv4
    port map (
            O => \N__12312\,
            I => \M_this_vram_read_data_1\
        );

    \I__1106\ : InMux
    port map (
            O => \N__12309\,
            I => \N__12306\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__12306\,
            I => \this_vga_ramdac.i2_mux_0\
        );

    \I__1104\ : InMux
    port map (
            O => \N__12303\,
            I => \N__12297\
        );

    \I__1103\ : InMux
    port map (
            O => \N__12302\,
            I => \N__12297\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__12297\,
            I => \this_pixel_clk_M_counter_q_i_1\
        );

    \I__1101\ : InMux
    port map (
            O => \N__12294\,
            I => \N__12289\
        );

    \I__1100\ : InMux
    port map (
            O => \N__12293\,
            I => \N__12286\
        );

    \I__1099\ : InMux
    port map (
            O => \N__12292\,
            I => \N__12283\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__12289\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__12286\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__12283\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__1095\ : InMux
    port map (
            O => \N__12276\,
            I => \N__12272\
        );

    \I__1094\ : InMux
    port map (
            O => \N__12275\,
            I => \N__12269\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__12272\,
            I => \N__12263\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__12269\,
            I => \N__12263\
        );

    \I__1091\ : InMux
    port map (
            O => \N__12268\,
            I => \N__12259\
        );

    \I__1090\ : Span4Mux_v
    port map (
            O => \N__12263\,
            I => \N__12254\
        );

    \I__1089\ : InMux
    port map (
            O => \N__12262\,
            I => \N__12251\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__12259\,
            I => \N__12248\
        );

    \I__1087\ : InMux
    port map (
            O => \N__12258\,
            I => \N__12245\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__12257\,
            I => \N__12241\
        );

    \I__1085\ : Span4Mux_h
    port map (
            O => \N__12254\,
            I => \N__12236\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__12251\,
            I => \N__12236\
        );

    \I__1083\ : Span4Mux_h
    port map (
            O => \N__12248\,
            I => \N__12231\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__12245\,
            I => \N__12231\
        );

    \I__1081\ : InMux
    port map (
            O => \N__12244\,
            I => \N__12228\
        );

    \I__1080\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12225\
        );

    \I__1079\ : Odrv4
    port map (
            O => \N__12236\,
            I => \this_vga_ramdac.N_880_i_reto\
        );

    \I__1078\ : Odrv4
    port map (
            O => \N__12231\,
            I => \this_vga_ramdac.N_880_i_reto\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__12228\,
            I => \this_vga_ramdac.N_880_i_reto\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__12225\,
            I => \this_vga_ramdac.N_880_i_reto\
        );

    \I__1075\ : InMux
    port map (
            O => \N__12216\,
            I => \N__12213\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__12213\,
            I => \this_vga_signals.if_m8_0_a3_1_1_1\
        );

    \I__1073\ : CascadeMux
    port map (
            O => \N__12210\,
            I => \this_vga_signals.if_N_5_cascade_\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__12207\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\
        );

    \I__1071\ : InMux
    port map (
            O => \N__12204\,
            I => \N__12201\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__12201\,
            I => \N__12198\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__12198\,
            I => \this_vga_signals.mult1_un47_sum_c3_1_1_0\
        );

    \I__1068\ : InMux
    port map (
            O => \N__12195\,
            I => \N__12192\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__12192\,
            I => \N__12188\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__12191\,
            I => \N__12185\
        );

    \I__1065\ : Span4Mux_v
    port map (
            O => \N__12188\,
            I => \N__12182\
        );

    \I__1064\ : InMux
    port map (
            O => \N__12185\,
            I => \N__12179\
        );

    \I__1063\ : Odrv4
    port map (
            O => \N__12182\,
            I => \this_vga_ramdac.N_3301_reto\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__12179\,
            I => \this_vga_ramdac.N_3301_reto\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__12174\,
            I => \this_vga_signals.vvisibility_1_cascade_\
        );

    \I__1060\ : InMux
    port map (
            O => \N__12171\,
            I => \N__12168\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__12168\,
            I => \this_vga_ramdac.m16\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__12165\,
            I => \N__12162\
        );

    \I__1057\ : InMux
    port map (
            O => \N__12162\,
            I => \N__12159\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__12159\,
            I => \this_vga_signals.vaddress_5_0_6\
        );

    \I__1055\ : InMux
    port map (
            O => \N__12156\,
            I => \N__12153\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__12153\,
            I => \this_vga_signals.N_5\
        );

    \I__1053\ : InMux
    port map (
            O => \N__12150\,
            I => \N__12147\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__12147\,
            I => \this_vga_signals.if_m8_0_a3_1_1_0\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__12144\,
            I => \N__12141\
        );

    \I__1050\ : InMux
    port map (
            O => \N__12141\,
            I => \N__12138\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__12138\,
            I => \this_vga_signals.g2_5\
        );

    \I__1048\ : InMux
    port map (
            O => \N__12135\,
            I => \N__12132\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__12132\,
            I => \this_vga_signals.N_18_0\
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__12129\,
            I => \this_vga_signals.g0_7_0_cascade_\
        );

    \I__1045\ : InMux
    port map (
            O => \N__12126\,
            I => \N__12123\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__12123\,
            I => \N__12120\
        );

    \I__1043\ : Odrv4
    port map (
            O => \N__12120\,
            I => \this_vga_signals.g1_0_0_0\
        );

    \I__1042\ : CascadeMux
    port map (
            O => \N__12117\,
            I => \this_vga_signals.N_4_0_0_cascade_\
        );

    \I__1041\ : IoInMux
    port map (
            O => \N__12114\,
            I => \N__12111\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__12111\,
            I => \N__12108\
        );

    \I__1039\ : IoSpan4Mux
    port map (
            O => \N__12108\,
            I => \N__12105\
        );

    \I__1038\ : Span4Mux_s3_v
    port map (
            O => \N__12105\,
            I => \N__12102\
        );

    \I__1037\ : Span4Mux_h
    port map (
            O => \N__12102\,
            I => \N__12099\
        );

    \I__1036\ : Sp12to4
    port map (
            O => \N__12099\,
            I => \N__12096\
        );

    \I__1035\ : Odrv12
    port map (
            O => \N__12096\,
            I => \N_495\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__12093\,
            I => \this_vga_signals.un2_vsynclt8_cascade_\
        );

    \I__1033\ : IoInMux
    port map (
            O => \N__12090\,
            I => \N__12087\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__12087\,
            I => \N__12084\
        );

    \I__1031\ : Span4Mux_s2_v
    port map (
            O => \N__12084\,
            I => \N__12081\
        );

    \I__1030\ : Span4Mux_h
    port map (
            O => \N__12081\,
            I => \N__12078\
        );

    \I__1029\ : Span4Mux_v
    port map (
            O => \N__12078\,
            I => \N__12075\
        );

    \I__1028\ : Sp12to4
    port map (
            O => \N__12075\,
            I => \N__12072\
        );

    \I__1027\ : Span12Mux_v
    port map (
            O => \N__12072\,
            I => \N__12069\
        );

    \I__1026\ : Odrv12
    port map (
            O => \N__12069\,
            I => this_vga_signals_vsync_1_i
        );

    \I__1025\ : InMux
    port map (
            O => \N__12066\,
            I => \N__12063\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__12063\,
            I => \this_vga_signals.vsync_1_2\
        );

    \I__1023\ : InMux
    port map (
            O => \N__12060\,
            I => \N__12057\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__12057\,
            I => \this_vga_signals.vsync_1_3\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__12054\,
            I => \this_vga_signals.mult1_un47_sum_c3_1_1_0_cascade_\
        );

    \I__1020\ : IoInMux
    port map (
            O => \N__12051\,
            I => \N__12048\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__12048\,
            I => \N__12045\
        );

    \I__1018\ : Span12Mux_s10_h
    port map (
            O => \N__12045\,
            I => \N__12042\
        );

    \I__1017\ : Odrv12
    port map (
            O => \N__12042\,
            I => rgb_c_0
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__12039\,
            I => \this_vga_ramdac.i2_mux_cascade_\
        );

    \I__1015\ : InMux
    port map (
            O => \N__12036\,
            I => \N__12033\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__12033\,
            I => \N__12029\
        );

    \I__1013\ : InMux
    port map (
            O => \N__12032\,
            I => \N__12026\
        );

    \I__1012\ : Odrv12
    port map (
            O => \N__12029\,
            I => \this_vga_ramdac.N_3300_reto\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__12026\,
            I => \this_vga_ramdac.N_3300_reto\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__12021\,
            I => \this_vga_ramdac.m6_cascade_\
        );

    \I__1009\ : InMux
    port map (
            O => \N__12018\,
            I => \N__12015\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__12015\,
            I => \N__12012\
        );

    \I__1007\ : Span4Mux_v
    port map (
            O => \N__12012\,
            I => \N__12008\
        );

    \I__1006\ : InMux
    port map (
            O => \N__12011\,
            I => \N__12005\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__12008\,
            I => \this_vga_ramdac.N_3299_reto\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__12005\,
            I => \this_vga_ramdac.N_3299_reto\
        );

    \I__1003\ : IoInMux
    port map (
            O => \N__12000\,
            I => \N__11997\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__11997\,
            I => \N__11994\
        );

    \I__1001\ : Span4Mux_s2_h
    port map (
            O => \N__11994\,
            I => \N__11991\
        );

    \I__1000\ : Span4Mux_h
    port map (
            O => \N__11991\,
            I => \N__11988\
        );

    \I__999\ : Span4Mux_h
    port map (
            O => \N__11988\,
            I => \N__11985\
        );

    \I__998\ : Sp12to4
    port map (
            O => \N__11985\,
            I => \N__11982\
        );

    \I__997\ : Odrv12
    port map (
            O => \N__11982\,
            I => rgb_c_5
        );

    \I__996\ : CascadeMux
    port map (
            O => \N__11979\,
            I => \N__11976\
        );

    \I__995\ : InMux
    port map (
            O => \N__11976\,
            I => \N__11973\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__11973\,
            I => \N__11970\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__11970\,
            I => \this_vga_signals.N_729\
        );

    \I__992\ : InMux
    port map (
            O => \N__11967\,
            I => \un1_M_this_map_address_q_cry_1\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__11964\,
            I => \N__11961\
        );

    \I__990\ : CascadeBuf
    port map (
            O => \N__11961\,
            I => \N__11958\
        );

    \I__989\ : CascadeMux
    port map (
            O => \N__11958\,
            I => \N__11955\
        );

    \I__988\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11952\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__11952\,
            I => \N__11948\
        );

    \I__986\ : InMux
    port map (
            O => \N__11951\,
            I => \N__11945\
        );

    \I__985\ : Span4Mux_h
    port map (
            O => \N__11948\,
            I => \N__11942\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__11945\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__983\ : Odrv4
    port map (
            O => \N__11942\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__982\ : InMux
    port map (
            O => \N__11937\,
            I => \un1_M_this_map_address_q_cry_2\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__11934\,
            I => \N__11931\
        );

    \I__980\ : CascadeBuf
    port map (
            O => \N__11931\,
            I => \N__11928\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__11928\,
            I => \N__11925\
        );

    \I__978\ : InMux
    port map (
            O => \N__11925\,
            I => \N__11922\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__11922\,
            I => \N__11918\
        );

    \I__976\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11915\
        );

    \I__975\ : Span4Mux_h
    port map (
            O => \N__11918\,
            I => \N__11912\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__11915\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__973\ : Odrv4
    port map (
            O => \N__11912\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__972\ : InMux
    port map (
            O => \N__11907\,
            I => \un1_M_this_map_address_q_cry_3\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__11904\,
            I => \N__11901\
        );

    \I__970\ : CascadeBuf
    port map (
            O => \N__11901\,
            I => \N__11898\
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__11898\,
            I => \N__11895\
        );

    \I__968\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11892\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__11892\,
            I => \N__11888\
        );

    \I__966\ : InMux
    port map (
            O => \N__11891\,
            I => \N__11885\
        );

    \I__965\ : Span4Mux_h
    port map (
            O => \N__11888\,
            I => \N__11882\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__11885\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__963\ : Odrv4
    port map (
            O => \N__11882\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__962\ : InMux
    port map (
            O => \N__11877\,
            I => \un1_M_this_map_address_q_cry_4\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__11874\,
            I => \N__11871\
        );

    \I__960\ : CascadeBuf
    port map (
            O => \N__11871\,
            I => \N__11868\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__11868\,
            I => \N__11865\
        );

    \I__958\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11862\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__11862\,
            I => \N__11858\
        );

    \I__956\ : InMux
    port map (
            O => \N__11861\,
            I => \N__11855\
        );

    \I__955\ : Span4Mux_h
    port map (
            O => \N__11858\,
            I => \N__11852\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__11855\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__11852\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__952\ : InMux
    port map (
            O => \N__11847\,
            I => \un1_M_this_map_address_q_cry_5\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__11844\,
            I => \N__11841\
        );

    \I__950\ : CascadeBuf
    port map (
            O => \N__11841\,
            I => \N__11838\
        );

    \I__949\ : CascadeMux
    port map (
            O => \N__11838\,
            I => \N__11835\
        );

    \I__948\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11832\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__11832\,
            I => \N__11828\
        );

    \I__946\ : InMux
    port map (
            O => \N__11831\,
            I => \N__11825\
        );

    \I__945\ : Span4Mux_h
    port map (
            O => \N__11828\,
            I => \N__11822\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__11825\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__943\ : Odrv4
    port map (
            O => \N__11822\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__942\ : InMux
    port map (
            O => \N__11817\,
            I => \un1_M_this_map_address_q_cry_6\
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__11814\,
            I => \N__11811\
        );

    \I__940\ : CascadeBuf
    port map (
            O => \N__11811\,
            I => \N__11808\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__11808\,
            I => \N__11805\
        );

    \I__938\ : InMux
    port map (
            O => \N__11805\,
            I => \N__11802\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__11802\,
            I => \N__11798\
        );

    \I__936\ : InMux
    port map (
            O => \N__11801\,
            I => \N__11795\
        );

    \I__935\ : Span4Mux_h
    port map (
            O => \N__11798\,
            I => \N__11792\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__11795\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__11792\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__932\ : InMux
    port map (
            O => \N__11787\,
            I => \bfn_10_28_0_\
        );

    \I__931\ : InMux
    port map (
            O => \N__11784\,
            I => \un1_M_this_map_address_q_cry_8\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__11781\,
            I => \N__11778\
        );

    \I__929\ : CascadeBuf
    port map (
            O => \N__11778\,
            I => \N__11775\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__11775\,
            I => \N__11772\
        );

    \I__927\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11769\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__11769\,
            I => \N__11765\
        );

    \I__925\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11762\
        );

    \I__924\ : Span4Mux_h
    port map (
            O => \N__11765\,
            I => \N__11759\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__11762\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__11759\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__921\ : IoInMux
    port map (
            O => \N__11754\,
            I => \N__11751\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__11751\,
            I => \N__11748\
        );

    \I__919\ : Span12Mux_s1_h
    port map (
            O => \N__11748\,
            I => \N__11745\
        );

    \I__918\ : Odrv12
    port map (
            O => \N__11745\,
            I => rgb_c_2
        );

    \I__917\ : IoInMux
    port map (
            O => \N__11742\,
            I => \N__11739\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__11739\,
            I => \N__11736\
        );

    \I__915\ : Odrv12
    port map (
            O => \N__11736\,
            I => rgb_c_1
        );

    \I__914\ : IoInMux
    port map (
            O => \N__11733\,
            I => \N__11730\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__11730\,
            I => \N__11727\
        );

    \I__912\ : IoSpan4Mux
    port map (
            O => \N__11727\,
            I => \N__11724\
        );

    \I__911\ : Span4Mux_s2_h
    port map (
            O => \N__11724\,
            I => \N__11721\
        );

    \I__910\ : Span4Mux_h
    port map (
            O => \N__11721\,
            I => \N__11718\
        );

    \I__909\ : Span4Mux_v
    port map (
            O => \N__11718\,
            I => \N__11715\
        );

    \I__908\ : Span4Mux_v
    port map (
            O => \N__11715\,
            I => \N__11712\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__11712\,
            I => rgb_c_4
        );

    \I__906\ : InMux
    port map (
            O => \N__11709\,
            I => \N__11706\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__11706\,
            I => \N__11703\
        );

    \I__904\ : Odrv4
    port map (
            O => \N__11703\,
            I => \M_this_map_ram_write_data_4\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__11700\,
            I => \N__11697\
        );

    \I__902\ : InMux
    port map (
            O => \N__11697\,
            I => \N__11694\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__11694\,
            I => \N__11691\
        );

    \I__900\ : Odrv4
    port map (
            O => \N__11691\,
            I => \N_393_0\
        );

    \I__899\ : IoInMux
    port map (
            O => \N__11688\,
            I => \N__11685\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__11685\,
            I => \N__11682\
        );

    \I__897\ : IoSpan4Mux
    port map (
            O => \N__11682\,
            I => \N__11679\
        );

    \I__896\ : Span4Mux_s1_h
    port map (
            O => \N__11679\,
            I => \N__11676\
        );

    \I__895\ : Span4Mux_h
    port map (
            O => \N__11676\,
            I => \N__11673\
        );

    \I__894\ : Span4Mux_h
    port map (
            O => \N__11673\,
            I => \N__11670\
        );

    \I__893\ : Odrv4
    port map (
            O => \N__11670\,
            I => rgb_c_3
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__11667\,
            I => \N__11664\
        );

    \I__891\ : CascadeBuf
    port map (
            O => \N__11664\,
            I => \N__11661\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__11661\,
            I => \N__11658\
        );

    \I__889\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11654\
        );

    \I__888\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11651\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__11654\,
            I => \N__11648\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__11651\,
            I => \N__11643\
        );

    \I__885\ : Span4Mux_v
    port map (
            O => \N__11648\,
            I => \N__11643\
        );

    \I__884\ : Odrv4
    port map (
            O => \N__11643\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__11640\,
            I => \N__11637\
        );

    \I__882\ : CascadeBuf
    port map (
            O => \N__11637\,
            I => \N__11634\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__11634\,
            I => \N__11631\
        );

    \I__880\ : InMux
    port map (
            O => \N__11631\,
            I => \N__11628\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__11628\,
            I => \N__11624\
        );

    \I__878\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11621\
        );

    \I__877\ : Span4Mux_v
    port map (
            O => \N__11624\,
            I => \N__11618\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__11621\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__875\ : Odrv4
    port map (
            O => \N__11618\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__874\ : InMux
    port map (
            O => \N__11613\,
            I => \un1_M_this_map_address_q_cry_0\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__11610\,
            I => \N__11607\
        );

    \I__872\ : CascadeBuf
    port map (
            O => \N__11607\,
            I => \N__11604\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__11604\,
            I => \N__11601\
        );

    \I__870\ : InMux
    port map (
            O => \N__11601\,
            I => \N__11598\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__11598\,
            I => \N__11594\
        );

    \I__868\ : InMux
    port map (
            O => \N__11597\,
            I => \N__11591\
        );

    \I__867\ : Span4Mux_h
    port map (
            O => \N__11594\,
            I => \N__11588\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__11591\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__11588\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__864\ : IoInMux
    port map (
            O => \N__11583\,
            I => \N__11580\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__11580\,
            I => port_data_rw_i_i
        );

    \I__862\ : IoInMux
    port map (
            O => \N__11577\,
            I => \N__11574\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__11574\,
            I => \N__11571\
        );

    \I__860\ : Odrv12
    port map (
            O => \N__11571\,
            I => port_nmib_0_i
        );

    \I__859\ : IoInMux
    port map (
            O => \N__11568\,
            I => \N__11565\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__11565\,
            I => \N__11562\
        );

    \I__857\ : Odrv12
    port map (
            O => \N__11562\,
            I => this_vga_signals_vvisibility_i
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_20_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_6_0_\
        );

    \IN_MUX_bfv_20_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_vaddress_q_cry_7\,
            carryinitout => \bfn_20_7_0_\
        );

    \IN_MUX_bfv_19_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_5_0_\
        );

    \IN_MUX_bfv_19_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_haddress_q_cry_7\,
            carryinitout => \bfn_19_6_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_21_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_22_0_\
        );

    \IN_MUX_bfv_21_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \M_this_data_count_q_cry_7\,
            carryinitout => \bfn_21_23_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_24_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_11_0_\
        );

    \IN_MUX_bfv_21_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_6_0_\
        );

    \IN_MUX_bfv_21_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_vaddress_q_3_cry_7\,
            carryinitout => \bfn_21_7_0_\
        );

    \IN_MUX_bfv_19_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_7_0_\
        );

    \IN_MUX_bfv_19_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_haddress_q_2_cry_7\,
            carryinitout => \bfn_19_8_0_\
        );

    \IN_MUX_bfv_19_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_22_0_\
        );

    \IN_MUX_bfv_19_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_sprites_address_q_cry_7\,
            carryinitout => \bfn_19_23_0_\
        );

    \IN_MUX_bfv_10_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_27_0_\
        );

    \IN_MUX_bfv_10_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_map_address_q_cry_7\,
            carryinitout => \bfn_10_28_0_\
        );

    \IN_MUX_bfv_26_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_26_21_0_\
        );

    \IN_MUX_bfv_26_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \M_this_external_address_q_cry_7\,
            carryinitout => \bfn_26_22_0_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI67JU6_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14700\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_1332_g\
        );

    \this_reset_cond.M_stage_q_RNIC5C7_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__29698\,
            GLOBALBUFFEROUTPUT => \M_this_reset_cond_out_g_0\
        );

    \this_reset_cond.M_stage_q_RNIC5C7_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__25017\,
            GLOBALBUFFEROUTPUT => \N_404_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_vga_signals.port_data_rw_i_i_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__25547\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24980\,
            lcout => port_data_rw_i_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNINGI76_7_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__24979\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20603\,
            lcout => port_nmib_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_0_7_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20604\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => this_vga_signals_vvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12036\,
            in2 => \_gnd_net_\,
            in3 => \N__12276\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12018\,
            in2 => \_gnd_net_\,
            in3 => \N__12275\,
            lcout => rgb_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12477\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12268\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_4_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32417\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25294\,
            lcout => \M_this_map_ram_write_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI88JG2_9_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__20593\,
            in1 => \N__15831\,
            in2 => \N__11979\,
            in3 => \N__15678\,
            lcout => \N_393_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__12195\,
            in1 => \N__12258\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rgb_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_0_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25346\,
            in1 => \N__11657\,
            in2 => \N__25291\,
            in3 => \N__25295\,
            lcout => \M_this_map_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_27_0_\,
            carryout => \un1_M_this_map_address_q_cry_0\,
            clk => \N__36963\,
            ce => 'H',
            sr => \N__32207\
        );

    \M_this_map_address_q_1_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25352\,
            in1 => \N__11627\,
            in2 => \_gnd_net_\,
            in3 => \N__11613\,
            lcout => \M_this_map_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_0\,
            carryout => \un1_M_this_map_address_q_cry_1\,
            clk => \N__36963\,
            ce => 'H',
            sr => \N__32207\
        );

    \M_this_map_address_q_2_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25347\,
            in1 => \N__11597\,
            in2 => \_gnd_net_\,
            in3 => \N__11967\,
            lcout => \M_this_map_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_1\,
            carryout => \un1_M_this_map_address_q_cry_2\,
            clk => \N__36963\,
            ce => 'H',
            sr => \N__32207\
        );

    \M_this_map_address_q_3_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25353\,
            in1 => \N__11951\,
            in2 => \_gnd_net_\,
            in3 => \N__11937\,
            lcout => \M_this_map_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_2\,
            carryout => \un1_M_this_map_address_q_cry_3\,
            clk => \N__36963\,
            ce => 'H',
            sr => \N__32207\
        );

    \M_this_map_address_q_4_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25348\,
            in1 => \N__11921\,
            in2 => \_gnd_net_\,
            in3 => \N__11907\,
            lcout => \M_this_map_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_3\,
            carryout => \un1_M_this_map_address_q_cry_4\,
            clk => \N__36963\,
            ce => 'H',
            sr => \N__32207\
        );

    \M_this_map_address_q_5_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25350\,
            in1 => \N__11891\,
            in2 => \_gnd_net_\,
            in3 => \N__11877\,
            lcout => \M_this_map_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_4\,
            carryout => \un1_M_this_map_address_q_cry_5\,
            clk => \N__36963\,
            ce => 'H',
            sr => \N__32207\
        );

    \M_this_map_address_q_6_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25349\,
            in1 => \N__11861\,
            in2 => \_gnd_net_\,
            in3 => \N__11847\,
            lcout => \M_this_map_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_5\,
            carryout => \un1_M_this_map_address_q_cry_6\,
            clk => \N__36963\,
            ce => 'H',
            sr => \N__32207\
        );

    \M_this_map_address_q_7_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25351\,
            in1 => \N__11831\,
            in2 => \_gnd_net_\,
            in3 => \N__11817\,
            lcout => \M_this_map_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_6\,
            carryout => \un1_M_this_map_address_q_cry_7\,
            clk => \N__36963\,
            ce => 'H',
            sr => \N__32207\
        );

    \M_this_map_address_q_8_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25357\,
            in1 => \N__11801\,
            in2 => \_gnd_net_\,
            in3 => \N__11787\,
            lcout => \M_this_map_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_10_28_0_\,
            carryout => \un1_M_this_map_address_q_cry_8\,
            clk => \N__36966\,
            ce => 'H',
            sr => \N__32205\
        );

    \M_this_map_address_q_9_LC_10_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__11768\,
            in1 => \N__25358\,
            in2 => \_gnd_net_\,
            in3 => \N__11784\,
            lcout => \M_this_map_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36966\,
            ce => 'H',
            sr => \N__32205\
        );

    \this_vga_signals.un5_vaddress_g0_39_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010101011010"
        )
    port map (
            in0 => \N__17331\,
            in1 => \N__17160\,
            in2 => \N__16505\,
            in3 => \N__17058\,
            lcout => \this_vga_signals.N_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_5_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16783\,
            in2 => \_gnd_net_\,
            in3 => \N__16367\,
            lcout => \this_vga_signals.g2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12262\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12861\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001110111"
        )
    port map (
            in0 => \N__12403\,
            in1 => \N__12338\,
            in2 => \N__12440\,
            in3 => \N__12369\,
            lcout => OPEN,
            ltout => \this_vga_ramdac.i2_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__12032\,
            in1 => \N__29685\,
            in2 => \N__12039\,
            in3 => \N__12895\,
            lcout => \this_vga_ramdac.N_3300_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36909\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111011"
        )
    port map (
            in0 => \N__12404\,
            in1 => \N__12339\,
            in2 => \N__12441\,
            in3 => \N__12370\,
            lcout => OPEN,
            ltout => \this_vga_ramdac.m6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__12011\,
            in1 => \N__29684\,
            in2 => \N__12021\,
            in3 => \N__12894\,
            lcout => \this_vga_ramdac.N_3299_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36909\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_0_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12293\,
            lcout => \this_pixel_clk_M_counter_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36920\,
            ce => 'H',
            sr => \N__36028\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12456\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12244\,
            lcout => rgb_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15599\,
            in2 => \_gnd_net_\,
            in3 => \N__15069\,
            lcout => \this_vga_signals.N_729\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__15597\,
            in1 => \N__15825\,
            in2 => \_gnd_net_\,
            in3 => \N__15672\,
            lcout => \N_495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001111"
        )
    port map (
            in0 => \N__14945\,
            in1 => \N__14873\,
            in2 => \N__16811\,
            in3 => \N__16909\,
            lcout => OPEN,
            ltout => \this_vga_signals.un2_vsynclt8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__12066\,
            in1 => \N__12060\,
            in2 => \N__12093\,
            in3 => \N__16447\,
            lcout => this_vga_signals_vsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__14946\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17412\,
            lcout => \this_vga_signals.vsync_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__16765\,
            in1 => \N__16350\,
            in2 => \N__14797\,
            in3 => \N__16224\,
            lcout => \this_vga_signals.vsync_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_40_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110110110111"
        )
    port map (
            in0 => \N__16223\,
            in1 => \N__17411\,
            in2 => \N__16476\,
            in3 => \N__14783\,
            lcout => \this_vga_signals.if_m8_0_a3_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_2_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010010011"
        )
    port map (
            in0 => \N__16764\,
            in1 => \N__16446\,
            in2 => \N__16377\,
            in3 => \N__17140\,
            lcout => \this_vga_signals.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_38_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010000001111"
        )
    port map (
            in0 => \N__17139\,
            in1 => \N__17302\,
            in2 => \N__12165\,
            in3 => \N__17045\,
            lcout => \this_vga_signals.mult1_un47_sum_c3_1_1_0\,
            ltout => \this_vga_signals.mult1_un47_sum_c3_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_36_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__17303\,
            in1 => \_gnd_net_\,
            in2 => \N__12054\,
            in3 => \N__16795\,
            lcout => \this_vga_signals.g1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_2_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17313\,
            in2 => \_gnd_net_\,
            in3 => \N__15406\,
            lcout => \this_vga_signals.g0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_2_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__15408\,
            in1 => \N__16478\,
            in2 => \_gnd_net_\,
            in3 => \N__16365\,
            lcout => \this_vga_signals.vaddress_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101111010111"
        )
    port map (
            in0 => \N__17395\,
            in1 => \N__14367\,
            in2 => \N__16222\,
            in3 => \N__14753\,
            lcout => \this_vga_signals.if_m8_0_a3_1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_1_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__15407\,
            in1 => \N__16477\,
            in2 => \_gnd_net_\,
            in3 => \N__16366\,
            lcout => \this_vga_signals.vaddress_5_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_7_0_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110101"
        )
    port map (
            in0 => \N__12156\,
            in1 => \N__12150\,
            in2 => \N__12144\,
            in3 => \N__17314\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_37_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__16766\,
            in1 => \N__12135\,
            in2 => \N__12129\,
            in3 => \N__16109\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_4_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_34_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16110\,
            in1 => \N__12126\,
            in2 => \N__12117\,
            in3 => \N__14505\,
            lcout => \this_vga_signals.N_3_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16368\,
            in1 => \N__16217\,
            in2 => \N__16506\,
            in3 => \N__17406\,
            lcout => \this_vga_signals.M_vcounter_d7lto8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_7_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13359\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36893\,
            ce => \N__14157\,
            sr => \N__14109\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x0_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__17311\,
            in1 => \N__16148\,
            in2 => \N__16793\,
            in3 => \N__16093\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_8_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12636\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36893\,
            ce => \N__14157\,
            sr => \N__14109\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__16364\,
            in1 => \N__12216\,
            in2 => \_gnd_net_\,
            in3 => \N__15405\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001110"
        )
    port map (
            in0 => \N__15909\,
            in1 => \N__17310\,
            in2 => \N__12210\,
            in3 => \N__17118\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x1_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__17312\,
            in1 => \N__16789\,
            in2 => \N__12207\,
            in3 => \N__16094\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_31_N_4L6_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011100011000"
        )
    port map (
            in0 => \N__12204\,
            in1 => \N__17315\,
            in2 => \N__16819\,
            in3 => \N__16121\,
            lcout => \this_vga_signals.g0_31_N_4L6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__12171\,
            in1 => \N__29711\,
            in2 => \N__12191\,
            in3 => \N__12896\,
            lcout => \this_vga_ramdac.N_3301_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36897\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIBCAC_6_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16501\,
            in2 => \_gnd_net_\,
            in3 => \N__15710\,
            lcout => OPEN,
            ltout => \this_vga_signals.vvisibility_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_7_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100111"
        )
    port map (
            in0 => \N__16218\,
            in1 => \N__17407\,
            in2 => \N__12174\,
            in3 => \N__14798\,
            lcout => this_vga_signals_vvisibility,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000110110111"
        )
    port map (
            in0 => \N__12430\,
            in1 => \N__12398\,
            in2 => \N__12371\,
            in3 => \N__12334\,
            lcout => \this_vga_ramdac.m16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001101001101"
        )
    port map (
            in0 => \N__12337\,
            in1 => \N__12368\,
            in2 => \N__12405\,
            in3 => \N__12433\,
            lcout => OPEN,
            ltout => \this_vga_ramdac.m19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__12467\,
            in1 => \N__29680\,
            in2 => \N__12480\,
            in3 => \N__12891\,
            lcout => \this_vga_ramdac.N_3302_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36903\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001001110"
        )
    port map (
            in0 => \N__12892\,
            in1 => \N__12452\,
            in2 => \N__29699\,
            in3 => \N__12309\,
            lcout => \this_vga_ramdac.N_3303_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36903\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__12431\,
            in1 => \N__12397\,
            in2 => \_gnd_net_\,
            in3 => \N__12336\,
            lcout => \this_vga_ramdac.N_24_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_2_RNIH7PG8_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12726\,
            in1 => \N__13606\,
            in2 => \_gnd_net_\,
            in3 => \N__13568\,
            lcout => \M_pcounter_q_ret_2_RNIH7PG8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101100011"
        )
    port map (
            in0 => \N__12432\,
            in1 => \N__12399\,
            in2 => \N__12372\,
            in3 => \N__12335\,
            lcout => \this_vga_ramdac.i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_1_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36087\,
            in1 => \N__12303\,
            in2 => \_gnd_net_\,
            in3 => \N__12294\,
            lcout => \this_pixel_clk_M_counter_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.G_394_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__12302\,
            in1 => \N__12292\,
            in2 => \_gnd_net_\,
            in3 => \N__36086\,
            lcout => \this_vga_signals.GZ0Z_394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_q_ret_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__29715\,
            in1 => \N__13260\,
            in2 => \N__12257\,
            in3 => \N__12900\,
            lcout => \this_vga_ramdac.N_880_i_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36921\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3SF72_9_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__15827\,
            in1 => \N__15673\,
            in2 => \N__20589\,
            in3 => \N__15598\,
            lcout => \N_880_0\,
            ltout => \N_880_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIITNT4_9_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12573\,
            in3 => \N__13818\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNILLQLK_9_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__13258\,
            in1 => \N__13782\,
            in2 => \_gnd_net_\,
            in3 => \N__13668\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIS7VH6_9_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13259\,
            in2 => \_gnd_net_\,
            in3 => \N__14019\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_1_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12513\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36926\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_0_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12525\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36926\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_1_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33311\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25229\,
            lcout => \M_this_map_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_5_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36360\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25230\,
            lcout => \M_this_map_ram_write_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17682\,
            in1 => \N__12718\,
            in2 => \N__13923\,
            in3 => \N__13921\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            clk => \N__36861\,
            ce => 'H',
            sr => \N__14106\
        );

    \this_vga_signals.M_vcounter_q_1_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17684\,
            in1 => \N__14872\,
            in2 => \_gnd_net_\,
            in3 => \N__12483\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            clk => \N__36861\,
            ce => 'H',
            sr => \N__14106\
        );

    \this_vga_signals.M_vcounter_q_2_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17683\,
            in1 => \N__14944\,
            in2 => \_gnd_net_\,
            in3 => \N__12597\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            clk => \N__36861\,
            ce => 'H',
            sr => \N__14106\
        );

    \this_vga_signals.M_vcounter_q_3_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17685\,
            in1 => \N__16908\,
            in2 => \_gnd_net_\,
            in3 => \N__12594\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            clk => \N__36861\,
            ce => 'H',
            sr => \N__14106\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16718\,
            in2 => \_gnd_net_\,
            in3 => \N__12591\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16375\,
            in2 => \_gnd_net_\,
            in3 => \N__12588\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16495\,
            in2 => \_gnd_net_\,
            in3 => \N__12585\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17421\,
            in2 => \_gnd_net_\,
            in3 => \N__12582\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16233\,
            in2 => \_gnd_net_\,
            in3 => \N__12579\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_9_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14790\,
            in2 => \_gnd_net_\,
            in3 => \N__12576\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36869\,
            ce => \N__14154\,
            sr => \N__14108\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_8_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12632\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36869\,
            ce => \N__14154\,
            sr => \N__14108\
        );

    \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12631\,
            lcout => \this_vga_signals.M_vcounter_q_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36869\,
            ce => \N__14154\,
            sr => \N__14108\
        );

    \this_vga_signals.un5_vaddress_g0_18_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011010010001"
        )
    port map (
            in0 => \N__14415\,
            in1 => \N__17309\,
            in2 => \N__14406\,
            in3 => \N__17138\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__13383\,
            in1 => \N__13290\,
            in2 => \N__14214\,
            in3 => \N__12618\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100011101"
        )
    port map (
            in0 => \N__13407\,
            in1 => \N__14240\,
            in2 => \N__12612\,
            in3 => \N__14752\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010110000"
        )
    port map (
            in0 => \N__14366\,
            in1 => \N__12603\,
            in2 => \N__12609\,
            in3 => \N__15703\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100011000011"
        )
    port map (
            in0 => \N__15906\,
            in1 => \N__17308\,
            in2 => \N__12606\,
            in3 => \N__17026\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__13382\,
            in1 => \_gnd_net_\,
            in2 => \N__14213\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.vaddress_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100101010"
        )
    port map (
            in0 => \N__13406\,
            in1 => \N__14239\,
            in2 => \N__14770\,
            in3 => \N__14365\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__14876\,
            in1 => \N__14985\,
            in2 => \_gnd_net_\,
            in3 => \N__12642\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_i1_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIIADJ4E2_7_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__15531\,
            in1 => \N__13518\,
            in2 => \N__12699\,
            in3 => \N__12675\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_31_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101011010"
        )
    port map (
            in0 => \N__14316\,
            in1 => \N__12738\,
            in2 => \N__14973\,
            in3 => \N__13445\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_5_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_22_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001110000011"
        )
    port map (
            in0 => \N__12720\,
            in1 => \N__14875\,
            in2 => \N__12678\,
            in3 => \N__12660\,
            lcout => \this_vga_signals.mult1_un82_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_2_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13499\,
            in1 => \N__14500\,
            in2 => \N__16980\,
            in3 => \N__16114\,
            lcout => \this_vga_signals.g0_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_0_0_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16791\,
            in2 => \_gnd_net_\,
            in3 => \N__13500\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_i_x4_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_23_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011110000"
        )
    port map (
            in0 => \N__16952\,
            in1 => \N__12669\,
            in2 => \N__12663\,
            in3 => \N__12768\,
            lcout => \this_vga_signals.N_3_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_24_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16790\,
            in1 => \N__14499\,
            in2 => \N__16981\,
            in3 => \N__15348\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_12_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111110111"
        )
    port map (
            in0 => \N__14981\,
            in1 => \N__14085\,
            in2 => \N__12654\,
            in3 => \N__12651\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_1_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__16554\,
            in1 => \N__14307\,
            in2 => \N__12645\,
            in3 => \N__13446\,
            lcout => \this_vga_signals.N_5_i_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_2_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__16948\,
            in1 => \N__14073\,
            in2 => \_gnd_net_\,
            in3 => \N__16122\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_16_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110111010111"
        )
    port map (
            in0 => \N__14948\,
            in1 => \N__14497\,
            in2 => \N__12771\,
            in3 => \N__13498\,
            lcout => \this_vga_signals.N_5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_ns_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12762\,
            in2 => \N__14634\,
            in3 => \N__12756\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_ns\,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc3_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_31_N_2L1_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12750\,
            in3 => \N__15999\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_31_N_2L1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_31_N_5L8_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111010111101"
        )
    port map (
            in0 => \N__14498\,
            in1 => \N__12747\,
            in2 => \N__12741\,
            in3 => \N__16953\,
            lcout => \this_vga_signals.g0_31_N_5L8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__13896\,
            in1 => \N__13587\,
            in2 => \_gnd_net_\,
            in3 => \N__13556\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_pcounter_q_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__17615\,
            in1 => \_gnd_net_\,
            in2 => \N__12732\,
            in3 => \N__12822\,
            lcout => \this_vga_signals.N_2_0\,
            ltout => \this_vga_signals.N_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_2_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12729\,
            in3 => \N__13608\,
            lcout => \this_vga_signals.M_this_vga_signals_pixel_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36898\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14874\,
            in2 => \_gnd_net_\,
            in3 => \N__12719\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_d7lt3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIK8V32_2_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__14947\,
            in1 => \N__16947\,
            in2 => \N__12909\,
            in3 => \N__16794\,
            lcout => \this_vga_signals.M_vcounter_d7lt9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__12906\,
            in1 => \N__29679\,
            in2 => \N__12860\,
            in3 => \N__12893\,
            lcout => \this_vga_ramdac.N_3298_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36898\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__13588\,
            in1 => \N__12820\,
            in2 => \N__12839\,
            in3 => \N__13897\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_pcounter_q_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12835\,
            in2 => \N__12843\,
            in3 => \N__17614\,
            lcout => \this_vga_signals.N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_1_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__13590\,
            in1 => \N__12821\,
            in2 => \N__12840\,
            in3 => \N__13899\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36904\,
            ce => \N__17669\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_0_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__13898\,
            in1 => \N__13589\,
            in2 => \_gnd_net_\,
            in3 => \N__13557\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36904\,
            ce => \N__17669\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIS3ODH5_9_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__13262\,
            in1 => \N__13209\,
            in2 => \_gnd_net_\,
            in3 => \N__13725\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_1_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13629\,
            in1 => \N__13218\,
            in2 => \N__13200\,
            in3 => \N__13716\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un89_sum_axbxc3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI15V0FA_9_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__13261\,
            in1 => \N__13208\,
            in2 => \N__12789\,
            in3 => \N__13724\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIDAFV71_9_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__13266\,
            in1 => \N__13680\,
            in2 => \_gnd_net_\,
            in3 => \N__13179\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c2_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111000101011"
        )
    port map (
            in0 => \N__15332\,
            in1 => \N__13679\,
            in2 => \N__17760\,
            in3 => \N__13178\,
            lcout => \this_vga_signals.mult1_un82_sum_c2_0\,
            ltout => \this_vga_signals.mult1_un82_sum_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c3_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13196\,
            in2 => \N__13212\,
            in3 => \N__13628\,
            lcout => \this_vga_signals.mult1_un82_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m1_0_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15196\,
            in2 => \_gnd_net_\,
            in3 => \N__14007\,
            lcout => \this_vga_signals.if_m7_0_x4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc1_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13771\,
            in1 => \N__15331\,
            in2 => \N__15272\,
            in3 => \N__13667\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_2_0_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13842\,
            in2 => \_gnd_net_\,
            in3 => \N__14006\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_2_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100000011110"
        )
    port map (
            in0 => \N__15195\,
            in1 => \N__13811\,
            in2 => \N__13185\,
            in3 => \N__15126\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_0_2\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13640\,
            in2 => \N__13182\,
            in3 => \N__13770\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI1VTU_4_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__13167\,
            in1 => \N__13149\,
            in2 => \N__33939\,
            in3 => \N__33792\,
            lcout => \M_this_ppu_sprites_addr_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_0_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31263\,
            in2 => \_gnd_net_\,
            in3 => \N__25276\,
            lcout => \M_this_map_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_7_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25277\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34581\,
            lcout => \M_this_map_ram_write_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_4_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14254\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36856\,
            ce => \N__14155\,
            sr => \N__14104\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_4_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14255\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36856\,
            ce => \N__14155\,
            sr => \N__14104\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_5_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14273\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36856\,
            ce => \N__14155\,
            sr => \N__14104\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_6_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14168\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36856\,
            ce => \N__14155\,
            sr => \N__14104\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_7_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13354\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36862\,
            ce => \N__14150\,
            sr => \N__14107\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011111"
        )
    port map (
            in0 => \N__13381\,
            in1 => \_gnd_net_\,
            in2 => \N__14206\,
            in3 => \N__13278\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_1_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_8_rep1_esr_RNIE4021_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110101111"
        )
    port map (
            in0 => \N__14353\,
            in1 => \N__14771\,
            in2 => \N__13272\,
            in3 => \N__13405\,
            lcout => \this_vga_signals.SUM_2_i_1_2_3\,
            ltout => \this_vga_signals.SUM_2_i_1_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001101010"
        )
    port map (
            in0 => \N__15516\,
            in1 => \N__15489\,
            in2 => \N__13269\,
            in3 => \N__15426\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIG08B1_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110111011101"
        )
    port map (
            in0 => \N__14742\,
            in1 => \N__13404\,
            in2 => \N__14364\,
            in3 => \N__14237\,
            lcout => \this_vga_signals.SUM_2_i_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14196\,
            in1 => \N__14741\,
            in2 => \N__14241\,
            in3 => \N__13403\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13380\,
            in2 => \N__13362\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13355\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36862\,
            ce => \N__14150\,
            sr => \N__14107\
        );

    \this_vga_signals.un5_vaddress_g0_8_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000111101011"
        )
    port map (
            in0 => \N__13434\,
            in1 => \N__14382\,
            in2 => \N__13338\,
            in3 => \N__16166\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13326\,
            in2 => \N__13320\,
            in3 => \N__14373\,
            lcout => \this_vga_signals.N_4_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_x1_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000110110"
        )
    port map (
            in0 => \N__16720\,
            in1 => \N__16092\,
            in2 => \N__17327\,
            in3 => \N__14532\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_654_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110000110100"
        )
    port map (
            in0 => \N__17280\,
            in1 => \N__17027\,
            in2 => \N__15907\,
            in3 => \N__17114\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un47_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_x0_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010010001011"
        )
    port map (
            in0 => \N__16719\,
            in1 => \N__17282\,
            in2 => \N__13317\,
            in3 => \N__16091\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_654_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x0_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110111110"
        )
    port map (
            in0 => \N__16931\,
            in1 => \N__15992\,
            in2 => \N__16596\,
            in3 => \N__14580\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m2_1_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010000011001"
        )
    port map (
            in0 => \N__17028\,
            in1 => \N__15899\,
            in2 => \N__17141\,
            in3 => \N__17281\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1\,
            ltout => \this_vga_signals.mult1_un54_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m4_0_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16721\,
            in2 => \N__13455\,
            in3 => \N__16910\,
            lcout => \this_vga_signals.if_i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_ns_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14493\,
            in2 => \N__14571\,
            in3 => \N__13452\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110100101"
        )
    port map (
            in0 => \N__14624\,
            in1 => \N__16161\,
            in2 => \N__16376\,
            in3 => \N__13433\,
            lcout => \this_vga_signals.mult1_un61_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_1_x0_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010001001011"
        )
    port map (
            in0 => \N__17325\,
            in1 => \N__14536\,
            in2 => \N__16982\,
            in3 => \N__16107\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_1_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_1_ns_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__16108\,
            in1 => \N__16961\,
            in2 => \N__13422\,
            in3 => \N__13539\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_10_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101110110111"
        )
    port map (
            in0 => \N__13494\,
            in1 => \N__14972\,
            in2 => \N__13419\,
            in3 => \N__14492\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_0_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001111000000"
        )
    port map (
            in0 => \N__16932\,
            in1 => \N__13416\,
            in2 => \N__13410\,
            in3 => \N__14300\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__14625\,
            in1 => \N__17324\,
            in2 => \_gnd_net_\,
            in3 => \N__16732\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_x0_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16969\,
            in1 => \N__13496\,
            in2 => \N__14986\,
            in3 => \N__15995\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_axbxc3_0_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_ns_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14496\,
            in2 => \N__13533\,
            in3 => \N__13512\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_0\,
            ltout => \this_vga_signals.mult1_un82_sum_axbxc3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIVJPKIE_3_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14511\,
            in1 => \N__13506\,
            in2 => \N__13530\,
            in3 => \N__13461\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI2J0JQ31_3_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011010010"
        )
    port map (
            in0 => \N__13527\,
            in1 => \N__14832\,
            in2 => \N__13521\,
            in3 => \N__14430\,
            lcout => \this_vga_signals.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_x1_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13497\,
            in1 => \N__16962\,
            in2 => \N__14987\,
            in3 => \N__15993\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_0_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI6FOR21_3_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16788\,
            in1 => \N__14495\,
            in2 => \N__16983\,
            in3 => \N__16123\,
            lcout => \this_vga_signals.g1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14494\,
            in1 => \N__13495\,
            in2 => \N__16984\,
            in3 => \N__15994\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1\,
            ltout => \this_vga_signals.mult1_un68_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_c2_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001011111"
        )
    port map (
            in0 => \N__14980\,
            in1 => \N__16970\,
            in2 => \N__13464\,
            in3 => \N__14299\,
            lcout => \this_vga_signals.mult1_un68_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13607\,
            lcout => \this_vga_signals.M_pcounter_q_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_e_0_RNISGJ64_1_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001010101"
        )
    port map (
            in0 => \N__13866\,
            in1 => \N__16528\,
            in2 => \N__14825\,
            in3 => \N__14792\,
            lcout => \this_vga_signals.M_lcounter_d_0_sqmuxa\,
            ltout => \this_vga_signals.M_lcounter_d_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_0_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110001010101010"
        )
    port map (
            in0 => \N__13952\,
            in1 => \N__17681\,
            in2 => \N__13572\,
            in3 => \N__13908\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNIPGBM_0_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__13865\,
            in1 => \N__13951\,
            in2 => \_gnd_net_\,
            in3 => \N__14791\,
            lcout => \this_vga_signals.line_clk_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_0_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__18882\,
            in1 => \N__29678\,
            in2 => \N__19671\,
            in3 => \N__18861\,
            lcout => \this_ppu.M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13569\,
            lcout => \this_vga_signals.M_pcounter_q_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36894\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__14687\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17628\,
            lcout => \this_vga_signals.N_966_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__17560\,
            in1 => \N__15256\,
            in2 => \N__17759\,
            in3 => \N__14673\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_hcounter_d7lt7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000000000"
        )
    port map (
            in0 => \N__15656\,
            in1 => \N__13827\,
            in2 => \N__13545\,
            in3 => \N__15818\,
            lcout => \this_vga_signals.M_hcounter_d7_0\,
            ltout => \this_vga_signals.M_hcounter_d7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13542\,
            in3 => \N__17627\,
            lcout => \this_vga_signals.M_vcounter_q_501_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_0_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001100111001"
        )
    port map (
            in0 => \N__15197\,
            in1 => \N__13791\,
            in2 => \N__15263\,
            in3 => \N__14015\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_1_1_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13666\,
            in1 => \N__15253\,
            in2 => \_gnd_net_\,
            in3 => \N__13695\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_axbxc3_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13627\,
            in1 => \N__13710\,
            in2 => \N__13728\,
            in3 => \N__13769\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_m2_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100101101111"
        )
    port map (
            in0 => \N__15325\,
            in1 => \N__13626\,
            in2 => \N__17758\,
            in3 => \N__13701\,
            lcout => \this_vga_signals.mult1_un89_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000111010100"
        )
    port map (
            in0 => \N__15318\,
            in1 => \N__13768\,
            in2 => \N__15265\,
            in3 => \N__13664\,
            lcout => \this_vga_signals.mult1_un75_sum_c2_0\,
            ltout => \this_vga_signals.mult1_un75_sum_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_o4_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000110110111"
        )
    port map (
            in0 => \N__13694\,
            in1 => \N__17748\,
            in2 => \N__13704\,
            in3 => \N__17561\,
            lcout => \this_vga_signals.if_N_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110110010"
        )
    port map (
            in0 => \N__15317\,
            in1 => \N__13833\,
            in2 => \N__15264\,
            in3 => \N__13693\,
            lcout => \this_vga_signals.mult1_un75_sum_c3\,
            ltout => \this_vga_signals.mult1_un75_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13665\,
            in1 => \N__13778\,
            in2 => \N__13644\,
            in3 => \N__13641\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110101010111"
        )
    port map (
            in0 => \N__15635\,
            in1 => \N__15566\,
            in2 => \N__15064\,
            in3 => \N__15794\,
            lcout => \this_vga_signals.SUM_3_i_1_0\,
            ltout => \this_vga_signals.SUM_3_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_1_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011001101101"
        )
    port map (
            in0 => \N__15058\,
            in1 => \N__15114\,
            in2 => \N__13845\,
            in3 => \N__14033\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_0_1\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010000101101"
        )
    port map (
            in0 => \N__15180\,
            in1 => \N__13810\,
            in2 => \N__13836\,
            in3 => \N__15120\,
            lcout => \this_vga_signals.if_N_8_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17670\,
            in2 => \_gnd_net_\,
            in3 => \N__17497\,
            lcout => \this_vga_signals.N_966_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000001"
        )
    port map (
            in0 => \N__15115\,
            in1 => \N__15567\,
            in2 => \N__15065\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_hcounter_d7lto7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100100011"
        )
    port map (
            in0 => \N__15059\,
            in1 => \N__14034\,
            in2 => \N__15125\,
            in3 => \N__14052\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15178\,
            in2 => \N__13794\,
            in3 => \N__15119\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc1\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_3_0_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110101001111"
        )
    port map (
            in0 => \N__15235\,
            in1 => \N__15181\,
            in2 => \N__13785\,
            in3 => \N__14008\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIR18F4_9_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__15798\,
            in1 => \N__14058\,
            in2 => \N__15655\,
            in3 => \N__13983\,
            lcout => \M_hcounter_q_esr_RNIR18F4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15255\,
            in1 => \N__15327\,
            in2 => \N__17565\,
            in3 => \N__17756\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_473_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIEVMV1_6_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15056\,
            in1 => \N__15191\,
            in2 => \N__14061\,
            in3 => \N__15112\,
            lcout => \this_vga_signals.N_554\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110101000010"
        )
    port map (
            in0 => \N__15636\,
            in1 => \N__15568\,
            in2 => \N__15814\,
            in3 => \N__15054\,
            lcout => \this_vga_signals.N_735_0\,
            ltout => \this_vga_signals.N_735_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_2_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001100001"
        )
    port map (
            in0 => \N__15055\,
            in1 => \N__14051\,
            in2 => \N__14040\,
            in3 => \N__15110\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111010000"
        )
    port map (
            in0 => \N__15111\,
            in1 => \N__15177\,
            in2 => \N__14037\,
            in3 => \N__14032\,
            lcout => \this_vga_signals.mult1_un61_sum_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIL6NV1_7_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__15057\,
            in1 => \N__15581\,
            in2 => \N__13977\,
            in3 => \N__15113\,
            lcout => \this_vga_signals.hsync_1_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__15198\,
            in1 => \N__17757\,
            in2 => \N__15336\,
            in3 => \N__15273\,
            lcout => \this_vga_signals.N_507_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_6_LC_14_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34455\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25293\,
            lcout => \M_this_map_ram_write_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_e_0_1_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000010101010"
        )
    port map (
            in0 => \N__13859\,
            in1 => \N__13959\,
            in2 => \N__13938\,
            in3 => \N__13922\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36851\,
            ce => \N__17688\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_6_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14178\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36857\,
            ce => \N__14156\,
            sr => \N__14105\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__15385\,
            in1 => \N__16410\,
            in2 => \_gnd_net_\,
            in3 => \N__16302\,
            lcout => \this_vga_signals.vaddress_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_5_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14283\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36857\,
            ce => \N__14156\,
            sr => \N__14105\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15384\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16301\,
            lcout => \this_vga_signals.vaddress_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14262\,
            lcout => \this_vga_signals.M_vcounter_q_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36857\,
            ce => \N__14156\,
            sr => \N__14105\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010010101"
        )
    port map (
            in0 => \N__14238\,
            in1 => \N__14205\,
            in2 => \N__15394\,
            in3 => \N__14354\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14177\,
            lcout => \this_vga_signals.M_vcounter_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36857\,
            ce => \N__14156\,
            sr => \N__14105\
        );

    \this_vga_signals.un5_vaddress_g0_27_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__14544\,
            in1 => \_gnd_net_\,
            in2 => \N__16809\,
            in3 => \N__17244\,
            lcout => \this_vga_signals.g1_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_2_1_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110110"
        )
    port map (
            in0 => \N__17243\,
            in1 => \N__14626\,
            in2 => \N__14538\,
            in3 => \N__16779\,
            lcout => \this_vga_signals.g0_2_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_14_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110011001100"
        )
    port map (
            in0 => \N__15428\,
            in1 => \N__15518\,
            in2 => \N__15464\,
            in3 => \N__15494\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_21_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001101010"
        )
    port map (
            in0 => \N__15517\,
            in1 => \N__15490\,
            in2 => \N__15460\,
            in3 => \N__15427\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_i_2\,
            ltout => \this_vga_signals.mult1_un40_sum_axb1_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_19_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001101000011"
        )
    port map (
            in0 => \N__17143\,
            in1 => \N__14396\,
            in2 => \N__14385\,
            in3 => \N__17241\,
            lcout => \this_vga_signals.mult1_un47_sum_c3_2\,
            ltout => \this_vga_signals.mult1_un47_sum_c3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_0_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100101101100"
        )
    port map (
            in0 => \N__17242\,
            in1 => \N__16971\,
            in2 => \N__14376\,
            in3 => \N__16778\,
            lcout => \this_vga_signals.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_RNID73S_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15386\,
            in2 => \N__16335\,
            in3 => \N__14355\,
            lcout => \this_vga_signals.vaddress_6\,
            ltout => \this_vga_signals.vaddress_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000001111"
        )
    port map (
            in0 => \N__17240\,
            in1 => \N__17142\,
            in2 => \N__14322\,
            in3 => \N__17029\,
            lcout => \this_vga_signals.mult1_un47_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16035\,
            in1 => \N__16026\,
            in2 => \N__16592\,
            in3 => \N__15987\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__14488\,
            in1 => \_gnd_net_\,
            in2 => \N__14319\,
            in3 => \N__15951\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14487\,
            in2 => \N__16591\,
            in3 => \N__15985\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_ns_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14630\,
            in2 => \N__14598\,
            in3 => \N__14589\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_654_ns\,
            ltout => \this_vga_signals.mult1_un68_sum_axb1_654_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m1_3_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16957\,
            in2 => \N__14583\,
            in3 => \N__16784\,
            lcout => \this_vga_signals.if_m1_3\,
            ltout => \this_vga_signals.if_m1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x1_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111011010"
        )
    port map (
            in0 => \N__15986\,
            in1 => \N__16985\,
            in2 => \N__14574\,
            in3 => \N__16582\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_20_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000001111"
        )
    port map (
            in0 => \N__17322\,
            in1 => \N__17165\,
            in2 => \N__14559\,
            in3 => \N__17049\,
            lcout => \this_vga_signals.mult1_un47_sum_c3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111001"
        )
    port map (
            in0 => \N__15870\,
            in1 => \N__17323\,
            in2 => \N__16810\,
            in3 => \N__14537\,
            lcout => \this_vga_signals.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_0_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15003\,
            in1 => \N__14501\,
            in2 => \N__15918\,
            in3 => \N__16125\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_9_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14994\,
            in1 => \N__14421\,
            in2 => \N__14439\,
            in3 => \N__14436\,
            lcout => \this_vga_signals.N_3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_28_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__15864\,
            in1 => \N__16499\,
            in2 => \N__16821\,
            in3 => \N__17166\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_11_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_11_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__17326\,
            in1 => \N__15933\,
            in2 => \N__14424\,
            in3 => \N__15846\,
            lcout => \this_vga_signals.N_4_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__16029\,
            in1 => \N__16167\,
            in2 => \N__16820\,
            in3 => \N__16124\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_1_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010101111"
        )
    port map (
            in0 => \N__16973\,
            in1 => \_gnd_net_\,
            in2 => \N__14997\,
            in3 => \N__16818\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_7_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__18881\,
            in1 => \N__17847\,
            in2 => \_gnd_net_\,
            in3 => \N__21523\,
            lcout => \this_ppu.M_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36884\,
            ce => 'H',
            sr => \N__36015\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIGR3I_9_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15826\,
            in2 => \_gnd_net_\,
            in3 => \N__14793\,
            lcout => \this_vga_signals.g0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m5_s_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__14988\,
            in1 => \N__14883\,
            in2 => \_gnd_net_\,
            in3 => \N__14838\,
            lcout => \this_vga_signals.if_m5_s\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000000000"
        )
    port map (
            in0 => \N__17487\,
            in1 => \N__16536\,
            in2 => \N__14826\,
            in3 => \N__14799\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNI670G_1_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18758\,
            in1 => \N__17833\,
            in2 => \N__17811\,
            in3 => \N__17776\,
            lcout => \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI4I6I_2_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15316\,
            in2 => \_gnd_net_\,
            in3 => \N__15179\,
            lcout => \this_vga_signals.M_hcounter_d7lto4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14667\,
            in1 => \N__14652\,
            in2 => \_gnd_net_\,
            in3 => \N__28109\,
            lcout => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17548\,
            in2 => \N__17749\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17674\,
            in1 => \N__15326\,
            in2 => \_gnd_net_\,
            in3 => \N__15276\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__36905\,
            ce => 'H',
            sr => \N__17515\
        );

    \this_vga_signals.M_hcounter_q_3_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17671\,
            in1 => \N__15254\,
            in2 => \_gnd_net_\,
            in3 => \N__15201\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__36905\,
            ce => 'H',
            sr => \N__17515\
        );

    \this_vga_signals.M_hcounter_q_4_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17675\,
            in1 => \N__15190\,
            in2 => \_gnd_net_\,
            in3 => \N__15129\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__36905\,
            ce => 'H',
            sr => \N__17515\
        );

    \this_vga_signals.M_hcounter_q_5_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17672\,
            in1 => \N__15124\,
            in2 => \_gnd_net_\,
            in3 => \N__15072\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \N__36905\,
            ce => 'H',
            sr => \N__17515\
        );

    \this_vga_signals.M_hcounter_q_6_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17676\,
            in1 => \N__15063\,
            in2 => \_gnd_net_\,
            in3 => \N__15012\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \N__36905\,
            ce => 'H',
            sr => \N__17515\
        );

    \this_vga_signals.M_hcounter_q_7_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17673\,
            in1 => \N__15580\,
            in2 => \_gnd_net_\,
            in3 => \N__15009\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \N__36905\,
            ce => 'H',
            sr => \N__17515\
        );

    \this_vga_signals.M_hcounter_q_8_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17677\,
            in1 => \N__15654\,
            in2 => \_gnd_net_\,
            in3 => \N__15006\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \N__36905\,
            ce => 'H',
            sr => \N__17515\
        );

    \this_vga_signals.M_hcounter_q_esr_9_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15810\,
            in2 => \_gnd_net_\,
            in3 => \N__15834\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36911\,
            ce => \N__15759\,
            sr => \N__17517\
        );

    \this_sprites_ram.mem_mem_3_0_wclke_3_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__34995\,
            in1 => \N__34914\,
            in2 => \N__34820\,
            in3 => \N__34678\,
            lcout => \this_sprites_ram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_2_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35137\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25290\,
            lcout => \M_this_map_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI65531_7_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101111110"
        )
    port map (
            in0 => \N__16236\,
            in1 => \N__17427\,
            in2 => \N__16472\,
            in3 => \N__15714\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI3SF72_7_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__15690\,
            in1 => \N__15677\,
            in2 => \N__15603\,
            in3 => \N__15600\,
            lcout => \this_vga_signals.g0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001101010"
        )
    port map (
            in0 => \N__15519\,
            in1 => \N__15498\,
            in2 => \N__15468\,
            in3 => \N__15435\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_0_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__16466\,
            in1 => \N__16360\,
            in2 => \_gnd_net_\,
            in3 => \N__15393\,
            lcout => \this_vga_signals.vaddress_0_0_6\,
            ltout => \this_vga_signals.vaddress_0_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_25_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010010011001"
        )
    port map (
            in0 => \N__17259\,
            in1 => \N__17153\,
            in2 => \N__15351\,
            in3 => \N__17064\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_30_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__16467\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16750\,
            lcout => \this_vga_signals.g0_i_i_a5_1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__16027\,
            in1 => \N__16165\,
            in2 => \N__16792\,
            in3 => \N__16115\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_1\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16972\,
            in2 => \N__16038\,
            in3 => \N__16754\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16028\,
            in1 => \N__16589\,
            in2 => \N__16002\,
            in3 => \N__15988\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_29_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__17161\,
            in1 => \N__17304\,
            in2 => \N__15945\,
            in3 => \N__15859\,
            lcout => \this_vga_signals.g0_i_i_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHT721_5_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__16756\,
            in1 => \N__16468\,
            in2 => \_gnd_net_\,
            in3 => \N__16362\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_7_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100011000011"
        )
    port map (
            in0 => \N__17164\,
            in1 => \N__17307\,
            in2 => \N__15927\,
            in3 => \N__15924\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000001111"
        )
    port map (
            in0 => \N__17305\,
            in1 => \N__17162\,
            in2 => \N__15908\,
            in3 => \N__17062\,
            lcout => \this_vga_signals.mult1_un47_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_17_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101110110111"
        )
    port map (
            in0 => \N__16361\,
            in1 => \N__16755\,
            in2 => \N__16494\,
            in3 => \N__15860\,
            lcout => \this_vga_signals.N_7_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_26_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100010100101"
        )
    port map (
            in0 => \N__17306\,
            in1 => \N__17163\,
            in2 => \N__17073\,
            in3 => \N__17063\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_axb1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_0_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001001001011"
        )
    port map (
            in0 => \N__16986\,
            in1 => \N__16757\,
            in2 => \N__16599\,
            in3 => \N__16590\,
            lcout => \this_vga_signals.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNINAB95_1_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__19897\,
            in1 => \N__18950\,
            in2 => \N__19684\,
            in3 => \N__19711\,
            lcout => \this_ppu.un13_0\,
            ltout => \this_ppu.un13_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_6_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000000010"
        )
    port map (
            in0 => \N__18831\,
            in1 => \N__17346\,
            in2 => \N__16542\,
            in3 => \N__18663\,
            lcout => \this_ppu.M_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010001010"
        )
    port map (
            in0 => \N__16251\,
            in1 => \N__16235\,
            in2 => \N__16260\,
            in3 => \N__17423\,
            lcout => \this_ppu.M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIO1JM4_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__19709\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19896\,
            lcout => \this_ppu.M_line_clk_out_0\,
            ltout => \this_ppu.M_line_clk_out_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIC69A5_1_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19673\,
            in1 => \N__27714\,
            in2 => \N__16539\,
            in3 => \N__27802\,
            lcout => \this_ppu.un1_M_vaddress_q_2_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_5_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__16535\,
            in1 => \N__16500\,
            in2 => \_gnd_net_\,
            in3 => \N__16363\,
            lcout => \this_vga_signals.un4_lvisibility_1\,
            ltout => \this_vga_signals.un4_lvisibility_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIV6084_7_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010001010"
        )
    port map (
            in0 => \N__16250\,
            in1 => \N__16234\,
            in2 => \N__16170\,
            in3 => \N__17422\,
            lcout => \M_this_vga_signals_line_clk_0\,
            ltout => \M_this_vga_signals_line_clk_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIN5VV4_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__19710\,
            in1 => \_gnd_net_\,
            in2 => \N__17364\,
            in3 => \N__19672\,
            lcout => \this_ppu.M_count_d_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18580\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => \this_ppu.un1_M_count_q_1_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28749\,
            in2 => \N__17781\,
            in3 => \N__17361\,
            lcout => \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_0_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17834\,
            in2 => \N__28807\,
            in3 => \N__17358\,
            lcout => \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_1_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28753\,
            in2 => \N__18759\,
            in3 => \N__17355\,
            lcout => \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_2_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17809\,
            in2 => \N__28808\,
            in3 => \N__17352\,
            lcout => \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_3_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28757\,
            in2 => \N__18606\,
            in3 => \N__17349\,
            lcout => \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_4_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18662\,
            in2 => \N__28809\,
            in3 => \N__17337\,
            lcout => \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_5_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_7_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000011110"
        )
    port map (
            in0 => \N__18951\,
            in1 => \N__21519\,
            in2 => \N__18644\,
            in3 => \N__17334\,
            lcout => \this_ppu.M_count_q_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_2_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000000010"
        )
    port map (
            in0 => \N__18829\,
            in1 => \N__17841\,
            in2 => \N__18794\,
            in3 => \N__17835\,
            lcout => \this_ppu.M_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_4_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000000010"
        )
    port map (
            in0 => \N__18830\,
            in1 => \N__17817\,
            in2 => \N__18795\,
            in3 => \N__17810\,
            lcout => \this_ppu.M_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_1_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100100000000"
        )
    port map (
            in0 => \N__17780\,
            in1 => \N__18787\,
            in2 => \N__17790\,
            in3 => \N__18828\,
            lcout => \this_ppu.M_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_1_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__17556\,
            in1 => \N__17686\,
            in2 => \_gnd_net_\,
            in3 => \N__17732\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36892\,
            ce => 'H',
            sr => \N__17516\
        );

    \this_vga_signals.M_hcounter_q_0_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17687\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17555\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36892\,
            ce => 'H',
            sr => \N__17516\
        );

    \this_delay_clk.M_pipe_q_3_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17457\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_2_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17466\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36896\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__34994\,
            in1 => \N__34912\,
            in2 => \N__34819\,
            in3 => \N__34699\,
            lcout => \this_sprites_ram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_substate_q_RNO_0_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100111111111"
        )
    port map (
            in0 => \N__25711\,
            in1 => \N__25665\,
            in2 => \N__25833\,
            in3 => \N__31638\,
            lcout => \M_this_substate_q_s_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_i_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24900\,
            in2 => \_gnd_net_\,
            in3 => \N__36095\,
            lcout => \N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_464_tz_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__26430\,
            in1 => \N__31147\,
            in2 => \N__23536\,
            in3 => \N__26519\,
            lcout => \N_1294_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_7_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110011"
        )
    port map (
            in0 => \N__27050\,
            in1 => \N__26125\,
            in2 => \N__23782\,
            in3 => \N__26205\,
            lcout => \M_this_sprites_address_qc_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_7_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000101"
        )
    port map (
            in0 => \N__23748\,
            in1 => \N__27052\,
            in2 => \N__31337\,
            in3 => \N__31149\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_7_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000110000"
        )
    port map (
            in0 => \N__25503\,
            in1 => \N__23705\,
            in2 => \N__17877\,
            in3 => \N__26438\,
            lcout => OPEN,
            ltout => \N_597_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_7_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__23706\,
            in1 => \N__17865\,
            in2 => \N__17874\,
            in3 => \N__17871\,
            lcout => \M_this_sprites_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36919\,
            ce => 'H',
            sr => \N__32203\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_468_tz_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110000"
        )
    port map (
            in0 => \N__31148\,
            in1 => \N__26553\,
            in2 => \N__23783\,
            in3 => \N__26436\,
            lcout => \N_1298_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_8_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__26437\,
            in1 => \N__25504\,
            in2 => \N__20397\,
            in3 => \N__23468\,
            lcout => OPEN,
            ltout => \N_602_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_8_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__23469\,
            in1 => \N__17859\,
            in2 => \N__17850\,
            in3 => \N__18561\,
            lcout => \M_this_sprites_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36919\,
            ce => 'H',
            sr => \N__32203\
        );

    \M_this_sprites_address_q_RNO_0_8_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110101000101"
        )
    port map (
            in0 => \N__26204\,
            in1 => \N__23510\,
            in2 => \N__26130\,
            in3 => \N__27051\,
            lcout => \M_this_sprites_address_qc_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27054\,
            in2 => \_gnd_net_\,
            in3 => \N__31146\,
            lcout => \this_vga_signals.N_415_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_3_LC_16_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35830\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25266\,
            lcout => \M_this_map_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19469\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI0VTU_0_4_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__18543\,
            in1 => \N__33773\,
            in2 => \N__18531\,
            in3 => \N__33863\,
            lcout => \M_this_ppu_sprites_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIEH4G1_2_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__33772\,
            in1 => \N__27605\,
            in2 => \N__33888\,
            in3 => \N__19596\,
            lcout => \M_this_ppu_sprites_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19485\,
            in2 => \_gnd_net_\,
            in3 => \N__18123\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__19484\,
            in1 => \N__18132\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIBD3G1_1_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__27713\,
            in1 => \N__33771\,
            in2 => \N__33846\,
            in3 => \N__19611\,
            lcout => \M_this_ppu_sprites_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19486\,
            in2 => \_gnd_net_\,
            in3 => \N__18675\,
            lcout => \this_reset_cond.M_stage_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_1_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20686\,
            in1 => \N__18944\,
            in2 => \N__33845\,
            in3 => \N__36097\,
            lcout => OPEN,
            ltout => \this_ppu.M_state_q_srsts_i_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_1_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__20646\,
            in1 => \N__19740\,
            in2 => \N__18666\,
            in3 => \N__18857\,
            lcout => \this_ppu.M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNIEF0G_7_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18661\,
            in1 => \N__18605\,
            in2 => \N__18645\,
            in3 => \N__18582\,
            lcout => \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_5\,
            ltout => \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_2_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__18945\,
            in1 => \N__18906\,
            in2 => \N__18618\,
            in3 => \N__36103\,
            lcout => \this_ppu.M_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_1_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__27788\,
            in1 => \N__19683\,
            in2 => \N__27715\,
            in3 => \N__18856\,
            lcout => \this_ppu.M_vaddress_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36876\,
            ce => 'H',
            sr => \N__21484\
        );

    \this_ppu.M_vaddress_q_0_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001110011001100"
        )
    port map (
            in0 => \N__19715\,
            in1 => \N__27787\,
            in2 => \N__19688\,
            in3 => \N__19905\,
            lcout => \M_this_ppu_vram_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36876\,
            ce => 'H',
            sr => \N__21484\
        );

    \this_ppu.M_count_q_5_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000010"
        )
    port map (
            in0 => \N__18827\,
            in1 => \N__18604\,
            in2 => \N__18615\,
            in3 => \N__18786\,
            lcout => \this_ppu.M_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_0_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__18581\,
            in1 => \N__18777\,
            in2 => \_gnd_net_\,
            in3 => \N__18826\,
            lcout => \this_ppu.M_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_9_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__18957\,
            in1 => \_gnd_net_\,
            in2 => \N__19509\,
            in3 => \_gnd_net_\,
            lcout => \M_this_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_8_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__18681\,
            in1 => \N__19501\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_reset_cond.M_stage_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIKRC91_1_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18946\,
            in1 => \N__18915\,
            in2 => \_gnd_net_\,
            in3 => \N__18905\,
            lcout => \this_ppu.M_count_d_0_sqmuxa_1\,
            ltout => \this_ppu.M_count_d_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIN6OG6_0_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__19670\,
            in1 => \N__29662\,
            in2 => \N__18864\,
            in3 => \N__18849\,
            lcout => \this_ppu.N_1417_0\,
            ltout => \this_ppu.N_1417_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_3_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010010000"
        )
    port map (
            in0 => \N__18804\,
            in1 => \N__18751\,
            in2 => \N__18798\,
            in3 => \N__18778\,
            lcout => \this_ppu.M_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_6_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19507\,
            in2 => \_gnd_net_\,
            in3 => \N__19434\,
            lcout => \this_reset_cond.M_stage_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28086\,
            in1 => \N__18729\,
            in2 => \_gnd_net_\,
            in3 => \N__18714\,
            lcout => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_4_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__19505\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18696\,
            lcout => \this_reset_cond.M_stage_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_7_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19508\,
            in2 => \_gnd_net_\,
            in3 => \N__18687\,
            lcout => \this_reset_cond.M_stage_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_5_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__19506\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19440\,
            lcout => \this_reset_cond.M_stage_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36895\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28068\,
            in1 => \N__19428\,
            in2 => \_gnd_net_\,
            in3 => \N__19410\,
            lcout => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_11_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__33785\,
            in1 => \N__19395\,
            in2 => \N__19374\,
            in3 => \N__33906\,
            lcout => \this_sprites_ram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36899\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_13_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__33786\,
            in1 => \N__19353\,
            in2 => \N__19335\,
            in3 => \N__33907\,
            lcout => \this_sprites_ram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36899\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28069\,
            in1 => \N__19311\,
            in2 => \_gnd_net_\,
            in3 => \N__19296\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__21662\,
            in1 => \N__21757\,
            in2 => \N__19284\,
            in3 => \N__19281\,
            lcout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI0VTU_4_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__19275\,
            in1 => \N__19251\,
            in2 => \N__33927\,
            in3 => \N__33784\,
            lcout => \M_this_ppu_sprites_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18990\,
            in1 => \N__18975\,
            in2 => \_gnd_net_\,
            in3 => \N__28070\,
            lcout => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_substate_q_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110100010"
        )
    port map (
            in0 => \N__31555\,
            in1 => \N__23377\,
            in2 => \N__19539\,
            in3 => \N__25533\,
            lcout => \M_this_substate_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36906\,
            ce => 'H',
            sr => \N__36018\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_480_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000001"
        )
    port map (
            in0 => \N__22128\,
            in1 => \N__24359\,
            in2 => \N__22203\,
            in3 => \N__26555\,
            lcout => OPEN,
            ltout => \M_this_sprites_address_q_0_0_i_480_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_4_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000100"
        )
    port map (
            in0 => \N__19515\,
            in1 => \N__19527\,
            in2 => \N__19530\,
            in3 => \N__19521\,
            lcout => \M_this_sprites_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36912\,
            ce => 'H',
            sr => \N__32210\
        );

    \M_this_sprites_address_q_RNO_0_4_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100110001"
        )
    port map (
            in0 => \N__24275\,
            in1 => \N__26216\,
            in2 => \N__22202\,
            in3 => \N__26413\,
            lcout => \M_this_sprites_address_qc_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_4_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__25468\,
            in1 => \N__22127\,
            in2 => \_gnd_net_\,
            in3 => \N__27049\,
            lcout => \N_511_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_4_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001101"
        )
    port map (
            in0 => \N__22170\,
            in1 => \N__31103\,
            in2 => \N__32441\,
            in3 => \N__26412\,
            lcout => \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_5_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000010"
        )
    port map (
            in0 => \N__20277\,
            in1 => \N__20349\,
            in2 => \N__19584\,
            in3 => \N__20283\,
            lcout => \M_this_sprites_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36912\,
            ce => 'H',
            sr => \N__32210\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_484_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000001"
        )
    port map (
            in0 => \N__22421\,
            in1 => \N__24358\,
            in2 => \N__22392\,
            in3 => \N__26537\,
            lcout => \M_this_sprites_address_q_0_0_i_484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_492_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101011"
        )
    port map (
            in0 => \N__26536\,
            in1 => \N__22926\,
            in2 => \N__24367\,
            in3 => \N__22887\,
            lcout => \M_this_sprites_address_q_0_0_i_492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_3_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001101"
        )
    port map (
            in0 => \N__22422\,
            in1 => \N__31115\,
            in2 => \N__35831\,
            in3 => \N__26435\,
            lcout => \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_5_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000011"
        )
    port map (
            in0 => \N__26434\,
            in1 => \N__21919\,
            in2 => \N__36356\,
            in3 => \N__31117\,
            lcout => \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_i_0_0_a4_4_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31178\,
            in2 => \_gnd_net_\,
            in3 => \N__31116\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_659_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_4_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__25829\,
            in1 => \N__25744\,
            in2 => \N__19575\,
            in3 => \N__27073\,
            lcout => \M_this_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36922\,
            ce => 'H',
            sr => \N__36023\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_2_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000110000"
        )
    port map (
            in0 => \N__25505\,
            in1 => \N__22625\,
            in2 => \N__19563\,
            in3 => \N__27053\,
            lcout => OPEN,
            ltout => \N_572_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_2_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__22626\,
            in1 => \N__19626\,
            in2 => \N__19572\,
            in3 => \N__19569\,
            lcout => \M_this_sprites_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36927\,
            ce => 'H',
            sr => \N__32206\
        );

    \M_this_sprites_address_q_RNO_0_2_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001111"
        )
    port map (
            in0 => \N__26432\,
            in1 => \N__22691\,
            in2 => \N__24280\,
            in3 => \N__26206\,
            lcout => \M_this_sprites_address_qc_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_2_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001011"
        )
    port map (
            in0 => \N__31144\,
            in1 => \N__22703\,
            in2 => \N__35238\,
            in3 => \N__26431\,
            lcout => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_3_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001111"
        )
    port map (
            in0 => \N__26433\,
            in1 => \N__22420\,
            in2 => \N__24281\,
            in3 => \N__26207\,
            lcout => OPEN,
            ltout => \M_this_sprites_address_qc_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_3_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__19554\,
            in1 => \N__19548\,
            in2 => \N__19542\,
            in3 => \N__20403\,
            lcout => \M_this_sprites_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36927\,
            ce => 'H',
            sr => \N__32206\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0_6_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__25663\,
            in1 => \N__25746\,
            in2 => \_gnd_net_\,
            in3 => \N__25803\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_0_0_a2_1_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__25662\,
            in1 => \N__31646\,
            in2 => \_gnd_net_\,
            in3 => \N__23382\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_488_tz_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__24345\,
            in1 => \N__22690\,
            in2 => \_gnd_net_\,
            in3 => \N__26548\,
            lcout => \N_1318_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_10_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100110001"
        )
    port map (
            in0 => \N__26105\,
            in1 => \N__26217\,
            in2 => \N__24493\,
            in3 => \N__27045\,
            lcout => \M_this_sprites_address_qc_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_11_LC_17_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100110001"
        )
    port map (
            in0 => \N__26106\,
            in1 => \N__26218\,
            in2 => \N__34676\,
            in3 => \N__27046\,
            lcout => \M_this_sprites_address_qc_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_vscroll_cry_0_c_inv_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19617\,
            in2 => \N__27823\,
            in3 => \N__27868\,
            lcout => \this_ppu.M_this_oam_ram_read_data_i_16\,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \this_ppu.un2_vscroll_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19590\,
            in2 => \N__27720\,
            in3 => \N__19602\,
            lcout => \this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un2_vscroll_cry_0\,
            carryout => \this_ppu.un2_vscroll_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__27539\,
            in1 => \N__27604\,
            in2 => \_gnd_net_\,
            in3 => \N__19599\,
            lcout => \this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27659\,
            lcout => \M_this_oam_ram_read_data_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_0_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100011011000011"
        )
    port map (
            in0 => \N__33725\,
            in1 => \N__34267\,
            in2 => \N__20642\,
            in3 => \N__19842\,
            lcout => \M_this_ppu_vram_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36864\,
            ce => 'H',
            sr => \N__21068\
        );

    \this_ppu.M_state_q_RNIQKAOF_3_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20669\,
            in2 => \_gnd_net_\,
            in3 => \N__19841\,
            lcout => \this_ppu.N_124\,
            ltout => \this_ppu.N_124_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_4_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000110010"
        )
    port map (
            in0 => \N__20687\,
            in1 => \N__29697\,
            in2 => \N__19734\,
            in3 => \N__24852\,
            lcout => \this_ppu.M_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_2_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__27789\,
            in1 => \N__27703\,
            in2 => \N__27602\,
            in3 => \N__21528\,
            lcout => \this_ppu.M_vaddress_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36877\,
            ce => 'H',
            sr => \N__21494\
        );

    \this_ppu.M_vaddress_q_6_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__27249\,
            in1 => \N__27319\,
            in2 => \_gnd_net_\,
            in3 => \N__19727\,
            lcout => \M_this_ppu_map_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36877\,
            ce => 'H',
            sr => \N__21494\
        );

    \this_ppu.M_vaddress_q_RNI3FOP5_4_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27461\,
            in1 => \N__27399\,
            in2 => \N__27606\,
            in3 => \N__20620\,
            lcout => \this_ppu.un1_M_vaddress_q_2_c5\,
            ltout => \this_ppu.un1_M_vaddress_q_2_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_5_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19731\,
            in3 => \N__27317\,
            lcout => \M_this_ppu_map_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36886\,
            ce => 'H',
            sr => \N__21474\
        );

    \this_ppu.M_vaddress_q_7_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__27250\,
            in1 => \N__27318\,
            in2 => \N__27958\,
            in3 => \N__19728\,
            lcout => \M_this_ppu_map_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36886\,
            ce => 'H',
            sr => \N__21474\
        );

    \this_ppu.M_vaddress_q_3_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__20621\,
            in1 => \N__27601\,
            in2 => \_gnd_net_\,
            in3 => \N__27462\,
            lcout => \M_this_ppu_map_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36886\,
            ce => 'H',
            sr => \N__21474\
        );

    \this_ppu.line_clk.M_last_q_RNI3BB75_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__19716\,
            in1 => \N__36098\,
            in2 => \N__19689\,
            in3 => \N__19904\,
            lcout => \this_ppu.M_last_q_RNI3BB75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28094\,
            in1 => \N__19881\,
            in2 => \_gnd_net_\,
            in3 => \N__19860\,
            lcout => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.vram_en_i_a2_0_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19796\,
            in1 => \N__21716\,
            in2 => \N__20006\,
            in3 => \N__19751\,
            lcout => \this_ppu.vram_en_i_a2Z0Z_0\,
            ltout => \this_ppu.vram_en_i_a2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIUTM1G_3_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33760\,
            in2 => \N__19824\,
            in3 => \N__20670\,
            lcout => \M_this_ppu_vram_en_0\,
            ltout => \M_this_ppu_vram_en_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNINDU1G_1_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33031\,
            in2 => \N__19821\,
            in3 => \N__34283\,
            lcout => \this_ppu.un1_M_haddress_q_3_c2\,
            ltout => \this_ppu.un1_M_haddress_q_3_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI4T92G_4_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21416\,
            in1 => \N__21334\,
            in2 => \N__19818\,
            in3 => \N__32743\,
            lcout => \this_ppu.un1_M_haddress_q_3_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__19815\,
            in1 => \N__20235\,
            in2 => \N__21766\,
            in3 => \N__19809\,
            lcout => \M_this_ppu_vram_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__21753\,
            in1 => \N__19785\,
            in2 => \N__21666\,
            in3 => \N__19779\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__21765\,
            in1 => \N__19773\,
            in2 => \N__19761\,
            in3 => \N__28020\,
            lcout => \M_this_ppu_vram_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28088\,
            in1 => \N__20268\,
            in2 => \_gnd_net_\,
            in3 => \N__20250\,
            lcout => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIITVO4_0_7_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24951\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => dma_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28087\,
            in1 => \N__20052\,
            in2 => \_gnd_net_\,
            in3 => \N__20037\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__21661\,
            in1 => \N__21763\,
            in2 => \N__20019\,
            in3 => \N__21831\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__21764\,
            in1 => \N__19911\,
            in2 => \N__20016\,
            in3 => \N__19950\,
            lcout => \M_this_ppu_vram_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28089\,
            in1 => \N__19983\,
            in2 => \_gnd_net_\,
            in3 => \N__19965\,
            lcout => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19944\,
            in1 => \N__19929\,
            in2 => \_gnd_net_\,
            in3 => \N__28090\,
            lcout => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_9_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__25047\,
            in1 => \N__25118\,
            in2 => \N__27180\,
            in3 => \N__25162\,
            lcout => \M_this_state_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36913\,
            ce => 'H',
            sr => \N__36016\
        );

    \this_vga_signals.un1_M_this_state_q_19_i_0_o2_0_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__25119\,
            in1 => \N__25155\,
            in2 => \_gnd_net_\,
            in3 => \N__25046\,
            lcout => \this_vga_signals.N_419_0\,
            ltout => \this_vga_signals.N_419_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_19_i_0_o2_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__25599\,
            in1 => \N__25568\,
            in2 => \N__20313\,
            in3 => \N__35253\,
            lcout => \N_440_0\,
            ltout => \N_440_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_19_i_0_o4_0_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20310\,
            in3 => \N__31639\,
            lcout => \this_vga_signals.N_467_0\,
            ltout => \this_vga_signals.N_467_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_5_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__20385\,
            in1 => \N__28192\,
            in2 => \N__20307\,
            in3 => \N__31126\,
            lcout => \M_this_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36913\,
            ce => 'H',
            sr => \N__36016\
        );

    \M_this_state_q_6_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__31125\,
            in1 => \N__20304\,
            in2 => \N__20298\,
            in3 => \N__29316\,
            lcout => \M_this_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36913\,
            ce => 'H',
            sr => \N__36016\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_7_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__29315\,
            in1 => \N__30404\,
            in2 => \_gnd_net_\,
            in3 => \N__26241\,
            lcout => \this_vga_signals.N_732\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_19_i_0_o4_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111101110"
        )
    port map (
            in0 => \N__25815\,
            in1 => \N__25664\,
            in2 => \_gnd_net_\,
            in3 => \N__25745\,
            lcout => \this_vga_signals.N_459_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_5_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__25483\,
            in1 => \N__21884\,
            in2 => \_gnd_net_\,
            in3 => \N__27048\,
            lcout => \N_510_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_5_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100110001"
        )
    port map (
            in0 => \N__24268\,
            in1 => \N__26214\,
            in2 => \N__21936\,
            in3 => \N__26403\,
            lcout => \M_this_sprites_address_qc_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0Z0Z_0_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000110000"
        )
    port map (
            in0 => \N__25482\,
            in1 => \N__23123\,
            in2 => \N__20334\,
            in3 => \N__27047\,
            lcout => OPEN,
            ltout => \N_562_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_0_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100000011"
        )
    port map (
            in0 => \N__23184\,
            in1 => \N__26215\,
            in2 => \N__20352\,
            in3 => \N__26404\,
            lcout => \M_this_sprites_address_qc_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_476_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000001"
        )
    port map (
            in0 => \N__21935\,
            in1 => \N__21885\,
            in2 => \N__24368\,
            in3 => \N__26554\,
            lcout => \M_this_sprites_address_q_0_0_i_476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_496_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000001"
        )
    port map (
            in0 => \N__23183\,
            in1 => \N__23127\,
            in2 => \N__24369\,
            in3 => \N__26538\,
            lcout => OPEN,
            ltout => \M_this_sprites_address_q_0_0_i_496_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_0_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100000000"
        )
    port map (
            in0 => \N__23185\,
            in1 => \N__24279\,
            in2 => \N__20343\,
            in3 => \N__20340\,
            lcout => \M_this_sprites_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36928\,
            ce => 'H',
            sr => \N__32211\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_0_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001101"
        )
    port map (
            in0 => \N__23182\,
            in1 => \N__31111\,
            in2 => \N__31355\,
            in3 => \N__26417\,
            lcout => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_0_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001000"
        )
    port map (
            in0 => \N__26416\,
            in1 => \N__25472\,
            in2 => \N__31143\,
            in3 => \N__27043\,
            lcout => \N_773\,
            ltout => \N_773_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_1_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100100011"
        )
    port map (
            in0 => \N__22925\,
            in1 => \N__26219\,
            in2 => \N__20325\,
            in3 => \N__26418\,
            lcout => OPEN,
            ltout => \M_this_sprites_address_qc_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_1_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__20370\,
            in1 => \N__20322\,
            in2 => \N__20316\,
            in3 => \N__20409\,
            lcout => \M_this_sprites_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36928\,
            ce => 'H',
            sr => \N__32211\
        );

    \M_this_sprites_address_q_13_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__26253\,
            in1 => \N__23400\,
            in2 => \N__26268\,
            in3 => \N__24378\,
            lcout => \M_this_sprites_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36931\,
            ce => 'H',
            sr => \N__32208\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_13_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000101"
        )
    port map (
            in0 => \N__34771\,
            in1 => \N__27006\,
            in2 => \N__34439\,
            in3 => \N__31120\,
            lcout => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_1_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__25498\,
            in1 => \N__22883\,
            in2 => \_gnd_net_\,
            in3 => \N__27017\,
            lcout => \N_896_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_3_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__25484\,
            in1 => \N__22385\,
            in2 => \_gnd_net_\,
            in3 => \N__27007\,
            lcout => \N_512_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_8_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001011"
        )
    port map (
            in0 => \N__31121\,
            in1 => \N__23518\,
            in2 => \N__33372\,
            in3 => \N__27016\,
            lcout => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1_5_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__25743\,
            in1 => \N__25649\,
            in2 => \_gnd_net_\,
            in3 => \N__25828\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_11_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001011"
        )
    port map (
            in0 => \N__31122\,
            in1 => \N__34651\,
            in2 => \N__32426\,
            in3 => \N__27044\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_11_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__26420\,
            in1 => \N__25501\,
            in2 => \N__20373\,
            in3 => \N__23444\,
            lcout => \N_617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_1_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000011"
        )
    port map (
            in0 => \N__26419\,
            in1 => \N__22947\,
            in2 => \N__33360\,
            in3 => \N__31123\,
            lcout => \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_456_tz_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__26415\,
            in1 => \N__24459\,
            in2 => \N__31145\,
            in3 => \N__26556\,
            lcout => OPEN,
            ltout => \N_1286_tz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_10_LC_18_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__20361\,
            in1 => \N__24396\,
            in2 => \N__20355\,
            in3 => \N__24414\,
            lcout => \M_this_sprites_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36941\,
            ce => 'H',
            sr => \N__32204\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_7_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010100000"
        )
    port map (
            in0 => \N__27038\,
            in1 => \N__31127\,
            in2 => \N__25499\,
            in3 => \N__26414\,
            lcout => \N_762\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_11_LC_18_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__20421\,
            in1 => \N__20415\,
            in2 => \N__24003\,
            in3 => \N__23448\,
            lcout => \M_this_sprites_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36941\,
            ce => 'H',
            sr => \N__32204\
        );

    \this_ppu.un1_M_haddress_q_cry_0_c_LC_19_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32798\,
            in2 => \N__20535\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_19_5_0_\,
            carryout => \this_ppu.un1_M_haddress_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_1_c_LC_19_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20514\,
            in2 => \N__32000\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_0\,
            carryout => \this_ppu.un1_M_haddress_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_2_c_LC_19_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20496\,
            in2 => \N__33130\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_1\,
            carryout => \this_ppu.un1_M_haddress_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_3_c_LC_19_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31811\,
            in2 => \N__20481\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_2\,
            carryout => \this_ppu.un1_M_haddress_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_4_c_LC_19_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31839\,
            in2 => \N__20460\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_3\,
            carryout => \this_ppu.un1_M_haddress_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_5_c_LC_19_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31743\,
            in2 => \N__20442\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_4\,
            carryout => \this_ppu.un1_M_haddress_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_6_c_LC_19_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31770\,
            in2 => \N__20739\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_5\,
            carryout => \this_ppu.un1_M_haddress_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_7_c_LC_19_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31875\,
            in2 => \N__20718\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_6\,
            carryout => \this_ppu.un1_M_haddress_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_7_THRU_LUT4_0_LC_19_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20538\,
            lcout => \this_ppu.un1_M_haddress_q_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32799\,
            in2 => \N__20531\,
            in3 => \N__34297\,
            lcout => \this_ppu.M_this_ppu_vram_addr_i_0\,
            ltout => OPEN,
            carryin => \bfn_19_7_0_\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_19_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32001\,
            in2 => \N__20513\,
            in3 => \N__33060\,
            lcout => \this_ppu.M_this_ppu_vram_addr_i_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_0\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20492\,
            in2 => \N__33135\,
            in3 => \N__32720\,
            lcout => \this_ppu.M_this_ppu_vram_addr_i_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_1\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24825\,
            in2 => \N__20477\,
            in3 => \N__21361\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_2\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_19_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20453\,
            in2 => \N__24390\,
            in3 => \N__21424\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_3\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_19_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31902\,
            in2 => \N__20438\,
            in3 => \N__21235\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_4\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_19_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31722\,
            in2 => \N__20735\,
            in3 => \N__21160\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_3\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_5\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21290\,
            in1 => \N__31854\,
            in2 => \N__20714\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_4\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_6\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_7_THRU_LUT4_0_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20697\,
            lcout => \this_ppu.un1_M_haddress_q_2_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_5_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36355\,
            lcout => \M_this_data_tmp_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36849\,
            ce => \N__30229\,
            sr => \N__36027\
        );

    \this_ppu.M_state_q_3_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__20694\,
            in1 => \N__36105\,
            in2 => \_gnd_net_\,
            in3 => \N__24848\,
            lcout => \this_ppu.M_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI6GOI_3_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33713\,
            in2 => \_gnd_net_\,
            in3 => \N__20665\,
            lcout => \this_ppu.N_122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_5_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33844\,
            in2 => \_gnd_net_\,
            in3 => \N__36104\,
            lcout => \this_ppu.M_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36872\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_4_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__27472\,
            in1 => \N__27585\,
            in2 => \N__27400\,
            in3 => \N__20625\,
            lcout => \M_this_ppu_map_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36878\,
            ce => 'H',
            sr => \N__21495\
        );

    \this_ppu.M_haddress_q_2_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__33039\,
            in1 => \N__34290\,
            in2 => \N__32737\,
            in3 => \N__21092\,
            lcout => \M_this_ppu_vram_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36887\,
            ce => 'H',
            sr => \N__21067\
        );

    \this_ppu.line_clk.M_last_q_RNIQRTEB_LC_19_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001100"
        )
    port map (
            in0 => \N__20585\,
            in1 => \N__29700\,
            in2 => \N__24939\,
            in3 => \N__21524\,
            lcout => \this_ppu.M_last_q_RNIQRTEB\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_4_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__21384\,
            in1 => \N__21336\,
            in2 => \N__32738\,
            in3 => \N__21417\,
            lcout => \M_this_ppu_map_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36900\,
            ce => 'H',
            sr => \N__21069\
        );

    \this_ppu.M_haddress_q_3_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__21335\,
            in1 => \N__32721\,
            in2 => \_gnd_net_\,
            in3 => \N__21383\,
            lcout => \M_this_ppu_map_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36900\,
            ce => 'H',
            sr => \N__21069\
        );

    \this_ppu.M_haddress_q_7_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__21258\,
            in1 => \N__21280\,
            in2 => \N__21219\,
            in3 => \N__21135\,
            lcout => \M_this_ppu_map_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36900\,
            ce => 'H',
            sr => \N__21069\
        );

    \this_ppu.M_haddress_q_5_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21202\,
            in2 => \_gnd_net_\,
            in3 => \N__21256\,
            lcout => \M_this_ppu_map_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36900\,
            ce => 'H',
            sr => \N__21069\
        );

    \this_ppu.M_haddress_q_6_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__21257\,
            in1 => \_gnd_net_\,
            in2 => \N__21218\,
            in3 => \N__21134\,
            lcout => \M_this_ppu_map_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36900\,
            ce => 'H',
            sr => \N__21069\
        );

    \this_ppu.M_haddress_q_1_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__33032\,
            in1 => \N__34303\,
            in2 => \_gnd_net_\,
            in3 => \N__21085\,
            lcout => \M_this_ppu_vram_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36900\,
            ce => 'H',
            sr => \N__21069\
        );

    \M_this_state_q_fast_9_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__27179\,
            in1 => \N__25164\,
            in2 => \N__25117\,
            in3 => \N__25056\,
            lcout => \M_this_state_q_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36907\,
            ce => 'H',
            sr => \N__36008\
        );

    \this_ppu.M_state_q_RNI0VTU_1_4_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__33776\,
            in1 => \N__21036\,
            in2 => \N__33934\,
            in3 => \N__21015\,
            lcout => \M_this_ppu_sprites_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28096\,
            in1 => \N__21807\,
            in2 => \_gnd_net_\,
            in3 => \N__21789\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__21660\,
            in1 => \N__21767\,
            in2 => \N__21771\,
            in3 => \N__21609\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__21768\,
            in1 => \N__21534\,
            in2 => \N__21723\,
            in3 => \N__21567\,
            lcout => \M_this_ppu_vram_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_12_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__33777\,
            in1 => \N__21699\,
            in2 => \N__33935\,
            in3 => \N__21684\,
            lcout => \this_sprites_ram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28095\,
            in1 => \N__21633\,
            in2 => \_gnd_net_\,
            in3 => \N__21618\,
            lcout => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21603\,
            in1 => \N__21585\,
            in2 => \_gnd_net_\,
            in3 => \N__28097\,
            lcout => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28098\,
            in1 => \N__21561\,
            in2 => \_gnd_net_\,
            in3 => \N__21552\,
            lcout => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_9_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001011"
        )
    port map (
            in0 => \N__30945\,
            in1 => \N__25951\,
            in2 => \N__35224\,
            in3 => \N__27042\,
            lcout => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_tr30_0_0_a2_0_a2_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__30944\,
            in1 => \_gnd_net_\,
            in2 => \N__29376\,
            in3 => \_gnd_net_\,
            lcout => \M_this_map_ram_write_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_4_LC_19_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21870\,
            lcout => \M_this_delay_clk_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28108\,
            in1 => \N__21861\,
            in2 => \_gnd_net_\,
            in3 => \N__21846\,
            lcout => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_6_0_0_m2_LC_19_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001011101"
        )
    port map (
            in0 => \N__26240\,
            in1 => \N__26518\,
            in2 => \N__30416\,
            in3 => \N__30943\,
            lcout => \this_vga_signals.N_505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_LC_19_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__25108\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25054\,
            lcout => \this_start_data_delay_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36923\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_i_a4_2_0_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__31624\,
            in1 => \N__29299\,
            in2 => \N__25173\,
            in3 => \N__27125\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_i_i_a4_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_q_0_i_a2_9_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__29297\,
            in1 => \N__35229\,
            in2 => \N__26787\,
            in3 => \N__30946\,
            lcout => \this_vga_signals.N_746\,
            ltout => \this_vga_signals.N_746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_6_0_0_i_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110011"
        )
    port map (
            in0 => \N__36325\,
            in1 => \N__29298\,
            in2 => \N__21825\,
            in3 => \N__21822\,
            lcout => \un1_M_this_state_q_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_i_a4_4_0_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__31213\,
            in1 => \N__28191\,
            in2 => \N__21816\,
            in3 => \N__26509\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_i_i_a4_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_3_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__30948\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27126\,
            lcout => \this_vga_signals.N_648\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_i_1_0_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010101"
        )
    port map (
            in0 => \N__31625\,
            in1 => \N__23388\,
            in2 => \N__23381\,
            in3 => \N__30947\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_i_i_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNIRO0N6_0_LC_19_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23181\,
            in2 => \N__23142\,
            in3 => \N__23141\,
            lcout => \M_this_sprites_address_q_RNIRO0N6Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_19_22_0_\,
            carryout => \un1_M_this_sprites_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22924\,
            in2 => \_gnd_net_\,
            in3 => \N__22872\,
            lcout => \un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_0\,
            carryout => \un1_M_this_sprites_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_19_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22775\,
            in3 => \N__22611\,
            lcout => \un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_1\,
            carryout => \un1_M_this_sprites_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22448\,
            in2 => \_gnd_net_\,
            in3 => \N__22371\,
            lcout => \un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_2\,
            carryout => \un1_M_this_sprites_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_19_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22204\,
            in2 => \_gnd_net_\,
            in3 => \N__22113\,
            lcout => \un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_3\,
            carryout => \un1_M_this_sprites_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_19_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21947\,
            in2 => \_gnd_net_\,
            in3 => \N__21876\,
            lcout => \un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_4\,
            carryout => \un1_M_this_sprites_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_19_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24071\,
            in2 => \_gnd_net_\,
            in3 => \N__21873\,
            lcout => \un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_5\,
            carryout => \un1_M_this_sprites_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_19_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23811\,
            in2 => \_gnd_net_\,
            in3 => \N__23691\,
            lcout => \un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_6\,
            carryout => \un1_M_this_sprites_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23517\,
            in2 => \_gnd_net_\,
            in3 => \N__23457\,
            lcout => \un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0\,
            ltout => OPEN,
            carryin => \bfn_19_23_0_\,
            carryout => \un1_M_this_sprites_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25875\,
            in2 => \_gnd_net_\,
            in3 => \N__23454\,
            lcout => \un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_8\,
            carryout => \un1_M_this_sprites_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24492\,
            in2 => \_gnd_net_\,
            in3 => \N__23451\,
            lcout => \un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_9\,
            carryout => \un1_M_this_sprites_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34675\,
            in2 => \_gnd_net_\,
            in3 => \N__23433\,
            lcout => \un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_10\,
            carryout => \un1_M_this_sprites_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_19_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34953\,
            in2 => \_gnd_net_\,
            in3 => \N__23430\,
            lcout => \un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_11\,
            carryout => \un1_M_this_sprites_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_19_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34748\,
            in2 => \_gnd_net_\,
            in3 => \N__23427\,
            lcout => \un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_9_LC_19_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__26424\,
            in1 => \N__25486\,
            in2 => \N__23424\,
            in3 => \N__23990\,
            lcout => \N_607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_13_LC_19_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__25485\,
            in1 => \N__26425\,
            in2 => \N__23409\,
            in3 => \N__23399\,
            lcout => \N_627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_6_LC_19_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__26989\,
            in1 => \N__25502\,
            in2 => \_gnd_net_\,
            in3 => \N__24305\,
            lcout => OPEN,
            ltout => \N_509_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_6_LC_19_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000100"
        )
    port map (
            in0 => \N__24288\,
            in1 => \N__24009\,
            in2 => \N__24372\,
            in3 => \N__24294\,
            lcout => \M_this_sprites_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36942\,
            ce => 'H',
            sr => \N__32209\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_472_LC_19_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101011"
        )
    port map (
            in0 => \N__26550\,
            in1 => \N__24366\,
            in2 => \N__24109\,
            in3 => \N__24306\,
            lcout => \M_this_sprites_address_q_0_0_i_472\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_6_LC_19_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000011"
        )
    port map (
            in0 => \N__26422\,
            in1 => \N__34445\,
            in2 => \N__24153\,
            in3 => \N__31105\,
            lcout => \this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_6_LC_19_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100010001"
        )
    port map (
            in0 => \N__26184\,
            in1 => \N__24282\,
            in2 => \N__26439\,
            in3 => \N__24108\,
            lcout => \M_this_sprites_address_qc_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_452_tz_LC_19_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__26421\,
            in1 => \N__31104\,
            in2 => \N__34677\,
            in3 => \N__26549\,
            lcout => \N_1282_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_460_tz_LC_19_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001010000"
        )
    port map (
            in0 => \N__26551\,
            in1 => \N__31124\,
            in2 => \N__25953\,
            in3 => \N__26423\,
            lcout => OPEN,
            ltout => \N_1290_tz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_9_LC_19_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__23991\,
            in1 => \N__25839\,
            in2 => \N__23979\,
            in3 => \N__23976\,
            lcout => \M_this_sprites_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36942\,
            ce => 'H',
            sr => \N__32209\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_10_LC_19_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001011"
        )
    port map (
            in0 => \N__31102\,
            in1 => \N__24455\,
            in2 => \N__35863\,
            in3 => \N__27005\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_10_LC_19_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000110000"
        )
    port map (
            in0 => \N__25500\,
            in1 => \N__24413\,
            in2 => \N__24399\,
            in3 => \N__26429\,
            lcout => \N_612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_address_q_0_i_a4_9_LC_19_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36344\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31706\,
            lcout => \N_560\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_axbxc1_LC_20_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31838\,
            in2 => \_gnd_net_\,
            in3 => \N__31810\,
            lcout => \this_ppu.un1_M_haddress_q_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_0_c_LC_20_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27870\,
            in2 => \N__27738\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_20_6_0_\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_1_c_LC_20_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27660\,
            in2 => \N__27624\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_0\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_2_c_LC_20_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27498\,
            in2 => \N__27543\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_1\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_3_c_LC_20_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32070\,
            in2 => \N__27435\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_2\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_4_c_LC_20_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32103\,
            in2 => \N__27362\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_3\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_5_c_LC_20_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27290\,
            in2 => \N__32142\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_4\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_6_c_LC_20_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29241\,
            in2 => \N__27222\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_5\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_7_c_LC_20_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29214\,
            in2 => \N__27927\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_6\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIF7IO_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__27903\,
            in1 => \N__24870\,
            in2 => \N__24864\,
            in3 => \N__24855\,
            lcout => \this_ppu.vscroll8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_20_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31815\,
            lcout => \M_this_oam_ram_read_data_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_2_LC_20_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35136\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36853\,
            ce => \N__30228\,
            sr => \N__36024\
        );

    \M_this_oam_address_q_0_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__30844\,
            in1 => \N__30648\,
            in2 => \_gnd_net_\,
            in3 => \N__33239\,
            lcout => \M_this_oam_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36879\,
            ce => 'H',
            sr => \N__32214\
        );

    \this_ppu.M_vaddress_q_RNINGCA_0_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27815\,
            in2 => \_gnd_net_\,
            in3 => \N__27869\,
            lcout => \this_ppu.un2_vscroll_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIO1A21_0_LC_20_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000001"
        )
    port map (
            in0 => \N__24819\,
            in1 => \N__33748\,
            in2 => \N__33897\,
            in3 => \N__27816\,
            lcout => \M_this_ppu_sprites_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI0A0E_6_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29334\,
            in2 => \_gnd_net_\,
            in3 => \N__27037\,
            lcout => \M_this_state_q_RNI0A0EZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI244K2_6_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__28143\,
            in1 => \N__24996\,
            in2 => \N__24879\,
            in3 => \N__29552\,
            lcout => OPEN,
            ltout => \M_this_state_q_RNI244K2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIITVO4_7_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001100"
        )
    port map (
            in0 => \N__25518\,
            in1 => \N__24885\,
            in2 => \N__24987\,
            in3 => \N__30376\,
            lcout => dma_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_address_q_0_i_o3_0_a4_5_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__35233\,
            in1 => \N__36334\,
            in2 => \_gnd_net_\,
            in3 => \N__29762\,
            lcout => \N_661\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_82_i_0_o2_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__27169\,
            in1 => \N__25163\,
            in2 => \N__25127\,
            in3 => \N__25055\,
            lcout => \this_vga_signals.N_428_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_a2_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__29363\,
            in1 => \N__24909\,
            in2 => \_gnd_net_\,
            in3 => \N__30586\,
            lcout => \N_861\,
            ltout => \N_861_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIG5R81_10_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__29418\,
            in1 => \N__28009\,
            in2 => \N__24888\,
            in3 => \N__27168\,
            lcout => dma_c4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un20_i_a2_4_a3_0_a4_2_1_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28008\,
            in1 => \N__30375\,
            in2 => \N__29374\,
            in3 => \N__27123\,
            lcout => this_vga_signals_un20_i_a2_4_a3_0_a4_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_13_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__30597\,
            in1 => \N__31002\,
            in2 => \N__27197\,
            in3 => \N__29417\,
            lcout => \M_this_state_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36924\,
            ce => 'H',
            sr => \N__36009\
        );

    \this_vga_signals.M_this_state_q_ns_i_0_0_o2_13_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31539\,
            in2 => \_gnd_net_\,
            in3 => \N__30285\,
            lcout => \N_460_0\,
            ltout => \N_460_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_11_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000100010"
        )
    port map (
            in0 => \N__29373\,
            in1 => \N__31001\,
            in2 => \N__25365\,
            in3 => \N__28010\,
            lcout => \M_this_state_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36924\,
            ce => 'H',
            sr => \N__36009\
        );

    \M_this_state_q_10_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__28011\,
            in1 => \N__30488\,
            in2 => \N__25362\,
            in3 => \N__25205\,
            lcout => \M_this_state_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36924\,
            ce => 'H',
            sr => \N__36009\
        );

    \this_vga_signals.M_this_external_address_qlde_i_0_a2_0_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__26775\,
            in1 => \N__29318\,
            in2 => \_gnd_net_\,
            in3 => \N__30966\,
            lcout => \this_vga_signals.N_745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_0_0_o2_1_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__25126\,
            in1 => \N__25153\,
            in2 => \_gnd_net_\,
            in3 => \N__25044\,
            lcout => \N_888_0\,
            ltout => \N_888_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_address_q_0_i_o3_0_a2_5_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26776\,
            in1 => \N__35218\,
            in2 => \N__25176\,
            in3 => \N__29319\,
            lcout => \M_this_oam_address_q_0_i_o3_0_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_i_a2_0_0_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__36313\,
            in1 => \_gnd_net_\,
            in2 => \N__26783\,
            in3 => \N__35219\,
            lcout => \this_vga_signals.N_779\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_en_1_sqmuxa_i_0_o4_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__30593\,
            in1 => \N__25154\,
            in2 => \N__25128\,
            in3 => \N__25045\,
            lcout => \N_413_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28193\,
            in2 => \_gnd_net_\,
            in3 => \N__29317\,
            lcout => \un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36092\,
            lcout => \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_5L8_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__25658\,
            in1 => \N__25595\,
            in2 => \N__25726\,
            in3 => \N__25817\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_5LZ0Z8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__35337\,
            in1 => \N__25569\,
            in2 => \N__25536\,
            in3 => \N__35346\,
            lcout => \M_this_substate_d_0_sqmuxa\,
            ltout => \M_this_substate_d_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_1_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__26316\,
            in1 => \_gnd_net_\,
            in2 => \N__25521\,
            in3 => \N__31003\,
            lcout => \M_this_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36932\,
            ce => 'H',
            sr => \N__36012\
        );

    \M_this_state_q_RNITB0L_3_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__28202\,
            in1 => \N__27124\,
            in2 => \_gnd_net_\,
            in3 => \N__26315\,
            lcout => dma_c4_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0_2_LC_20_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__25707\,
            in1 => \N__25816\,
            in2 => \_gnd_net_\,
            in3 => \N__31566\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_12_LC_20_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__26314\,
            in1 => \N__25506\,
            in2 => \N__25374\,
            in3 => \N__25391\,
            lcout => OPEN,
            ltout => \N_622_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_12_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__25392\,
            in1 => \N__25380\,
            in2 => \N__25383\,
            in3 => \N__26562\,
            lcout => \M_this_sprites_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36936\,
            ce => 'H',
            sr => \N__32212\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_448_tz_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__26313\,
            in1 => \N__31101\,
            in2 => \N__26552\,
            in3 => \N__34955\,
            lcout => \N_1278_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_12_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110001"
        )
    port map (
            in0 => \N__34954\,
            in1 => \N__36314\,
            in2 => \N__31142\,
            in3 => \N__26941\,
            lcout => \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_12_LC_20_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000011"
        )
    port map (
            in0 => \N__26942\,
            in1 => \N__26123\,
            in2 => \N__26220\,
            in3 => \N__34956\,
            lcout => \M_this_sprites_address_qc_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_i_o2_2_0_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26939\,
            in2 => \_gnd_net_\,
            in3 => \N__26311\,
            lcout => \this_vga_signals.N_427_0\,
            ltout => \this_vga_signals.N_427_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_444_tz_LC_20_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001100"
        )
    port map (
            in0 => \N__26312\,
            in1 => \N__34831\,
            in2 => \N__26271\,
            in3 => \N__31097\,
            lcout => \N_1274_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_13_LC_20_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000101"
        )
    port map (
            in0 => \N__26173\,
            in1 => \N__26940\,
            in2 => \N__26129\,
            in3 => \N__34818\,
            lcout => \M_this_sprites_address_qc_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_6_0_0_o2_LC_20_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27154\,
            in2 => \_gnd_net_\,
            in3 => \N__27110\,
            lcout => \this_vga_signals.N_889_0\,
            ltout => \this_vga_signals.N_889_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_LC_20_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__36323\,
            in1 => \N__31702\,
            in2 => \N__26223\,
            in3 => \N__30431\,
            lcout => \N_750\,
            ltout => \N_750_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_9_LC_20_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100001101"
        )
    port map (
            in0 => \N__26124\,
            in1 => \N__25952\,
            in2 => \N__25842\,
            in3 => \N__26985\,
            lcout => \M_this_sprites_address_qc_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_3_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__25818\,
            in1 => \N__25755\,
            in2 => \N__25742\,
            in3 => \N__27080\,
            lcout => \M_this_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36943\,
            ce => 'H',
            sr => \N__36019\
        );

    \M_this_state_q_8_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__31084\,
            in1 => \N__30377\,
            in2 => \N__27204\,
            in3 => \N__27161\,
            lcout => \M_this_state_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36943\,
            ce => 'H',
            sr => \N__36019\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_i_i_o2_0_LC_20_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100001111"
        )
    port map (
            in0 => \N__27160\,
            in1 => \N__27111\,
            in2 => \N__30442\,
            in3 => \N__31082\,
            lcout => \this_vga_signals.N_431_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_2_LC_20_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__31083\,
            in1 => \N__27090\,
            in2 => \N__27036\,
            in3 => \N__27081\,
            lcout => \M_this_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36943\,
            ce => 'H',
            sr => \N__36019\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_3_LC_20_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__28523\,
            in1 => \N__35826\,
            in2 => \N__34577\,
            in3 => \N__28547\,
            lcout => \N_250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_3_0_LC_20_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32383\,
            in1 => \N__34573\,
            in2 => \N__35846\,
            in3 => \N__31324\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_0_LC_20_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34444\,
            in2 => \N__26790\,
            in3 => \N__33355\,
            lcout => \this_vga_signals.N_743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_1_LC_20_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__33354\,
            in1 => \N__28545\,
            in2 => \N__36348\,
            in3 => \N__28521\,
            lcout => \N_228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_2_LC_20_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__28522\,
            in1 => \N__34443\,
            in2 => \N__35207\,
            in3 => \N__28546\,
            lcout => \N_248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_6_LC_21_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34441\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36848\,
            ce => \N__30230\,
            sr => \N__36029\
        );

    \M_this_data_tmp_q_esr_1_LC_21_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33411\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36848\,
            ce => \N__30230\,
            sr => \N__36029\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_21_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27864\,
            in2 => \N__27737\,
            in3 => \N__27825\,
            lcout => \this_ppu.M_this_ppu_vram_addr_i_7\,
            ltout => OPEN,
            carryin => \bfn_21_6_0_\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_21_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27716\,
            in1 => \N__27655\,
            in2 => \N__27623\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.M_vaddress_q_i_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_0\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_21_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27603\,
            in1 => \N__27497\,
            in2 => \N__27538\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.M_vaddress_q_i_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_1\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_21_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27882\,
            in2 => \N__27434\,
            in3 => \N__27476\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_5\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_2\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_21_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29142\,
            in2 => \N__27363\,
            in3 => \N__27404\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_6\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_3\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_21_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32031\,
            in2 => \N__27291\,
            in3 => \N__27335\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_7\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_4\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_21_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29265\,
            in2 => \N__27221\,
            in3 => \N__27272\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_8\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_5\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_21_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29178\,
            in2 => \N__27923\,
            in3 => \N__27968\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_9\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_6\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_21_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27906\,
            lcout => \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a4_16_LC_21_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27876\,
            in2 => \_gnd_net_\,
            in3 => \N__35707\,
            lcout => \M_this_oam_ram_write_data_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_21_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32066\,
            lcout => \M_this_oam_ram_read_data_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_16_LC_21_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31350\,
            lcout => \M_this_data_tmp_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36854\,
            ce => \N__34019\,
            sr => \N__36025\
        );

    \M_this_data_tmp_q_esr_17_LC_21_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33407\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36854\,
            ce => \N__34019\,
            sr => \N__36025\
        );

    \M_this_data_tmp_q_esr_23_LC_21_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34542\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36854\,
            ce => \N__34019\,
            sr => \N__36025\
        );

    \M_this_data_tmp_q_esr_3_LC_21_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35868\,
            lcout => \M_this_data_tmp_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36866\,
            ce => \N__30215\,
            sr => \N__36020\
        );

    \M_this_data_tmp_q_esr_7_LC_21_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34514\,
            lcout => \M_this_data_tmp_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36866\,
            ce => \N__30215\,
            sr => \N__36020\
        );

    \M_this_oam_address_q_RNI24IA1_1_1_LC_21_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__30558\,
            in1 => \N__30658\,
            in2 => \N__30853\,
            in3 => \N__36102\,
            lcout => \N_1412_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un20_i_a2_0_a3_0_a4_2_2_LC_21_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31205\,
            in1 => \N__29402\,
            in2 => \N__30605\,
            in3 => \N__30378\,
            lcout => this_vga_signals_un20_i_a2_0_a3_0_a4_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_6_0_0_a2_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__35220\,
            in1 => \N__36333\,
            in2 => \_gnd_net_\,
            in3 => \N__29763\,
            lcout => \this_vga_signals.N_747\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_en_iv_i_0_0_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28510\,
            in2 => \_gnd_net_\,
            in3 => \N__30438\,
            lcout => \N_25_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_21_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28137\,
            in1 => \N__28122\,
            in2 => \_gnd_net_\,
            in3 => \N__28110\,
            lcout => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_qlde_i_o2_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__29416\,
            in1 => \N__28007\,
            in2 => \_gnd_net_\,
            in3 => \N__30361\,
            lcout => \this_vga_signals.N_433_0\,
            ltout => \this_vga_signals.N_433_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_qlde_i_o2_0_LC_21_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27987\,
            in3 => \N__30279\,
            lcout => \this_vga_signals.N_442_0\,
            ltout => \this_vga_signals.N_442_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_qlde_i_a4_0_LC_21_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__29329\,
            in1 => \N__28203\,
            in2 => \N__27984\,
            in3 => \N__31000\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_719_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_qlde_i_1_LC_21_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__29548\,
            in1 => \N__30323\,
            in2 => \N__27981\,
            in3 => \N__30480\,
            lcout => \this_vga_signals.M_this_data_count_qlde_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_2_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__28215\,
            in1 => \N__31670\,
            in2 => \N__28233\,
            in3 => \N__31486\,
            lcout => \M_this_data_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36933\,
            ce => \N__31392\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_a3_0_a4_0_2_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__28195\,
            in1 => \_gnd_net_\,
            in2 => \N__36332\,
            in3 => \N__36090\,
            lcout => \this_vga_signals_M_this_data_count_q_3_0_a3_0_a4_0_2\,
            ltout => \this_vga_signals_M_this_data_count_q_3_0_a3_0_a4_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_i_i_10_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001111011111"
        )
    port map (
            in0 => \N__29751\,
            in1 => \N__35211\,
            in2 => \N__28209\,
            in3 => \N__28260\,
            lcout => OPEN,
            ltout => \N_307_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_10_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111000011011"
        )
    port map (
            in0 => \N__31487\,
            in1 => \N__28302\,
            in2 => \N__28206\,
            in3 => \N__29518\,
            lcout => \M_this_data_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36933\,
            ce => \N__31392\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_i_i_a2_10_LC_21_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__36089\,
            in1 => \N__28194\,
            in2 => \_gnd_net_\,
            in3 => \N__31076\,
            lcout => \N_755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_0_a4_0_1_13_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__36303\,
            in1 => \N__29750\,
            in2 => \N__35228\,
            in3 => \N__36088\,
            lcout => \this_vga_signals.N_665_1\,
            ltout => \this_vga_signals.N_665_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_q_3_0_0_13_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36302\,
            in2 => \N__28149\,
            in3 => \N__28259\,
            lcout => OPEN,
            ltout => \M_this_data_count_q_3_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_13_LC_21_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111000011011"
        )
    port map (
            in0 => \N__31488\,
            in1 => \N__29136\,
            in2 => \N__28146\,
            in3 => \N__29819\,
            lcout => \M_this_data_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36933\,
            ce => \N__31392\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_11_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__28290\,
            in1 => \N__31479\,
            in2 => \N__35847\,
            in3 => \N__28263\,
            lcout => \M_this_data_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36937\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_12_LC_21_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__28278\,
            in1 => \N__31480\,
            in2 => \N__32413\,
            in3 => \N__28264\,
            lcout => \M_this_data_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36937\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_14_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__28261\,
            in1 => \N__28578\,
            in2 => \N__34442\,
            in3 => \N__31483\,
            lcout => \M_this_data_count_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36937\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_15_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__28563\,
            in1 => \N__31481\,
            in2 => \N__34569\,
            in3 => \N__28265\,
            lcout => \M_this_data_count_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36937\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_8_LC_21_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__28262\,
            in1 => \N__28329\,
            in2 => \N__31362\,
            in3 => \N__31484\,
            lcout => \M_this_data_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36937\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_9_LC_21_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__28317\,
            in1 => \N__31482\,
            in2 => \N__33391\,
            in3 => \N__28266\,
            lcout => \M_this_data_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36937\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_0_LC_21_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31485\,
            in2 => \_gnd_net_\,
            in3 => \N__29586\,
            lcout => \M_this_data_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36937\,
            ce => \N__31400\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_c_0_LC_21_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29585\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_21_22_0_\,
            carryout => \M_this_data_count_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_0_THRU_LUT4_0_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28980\,
            in2 => \N__30030\,
            in3 => \N__28236\,
            lcout => \M_this_data_count_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_0\,
            carryout => \M_this_data_count_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_2_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29601\,
            in2 => \N__29046\,
            in3 => \N__28221\,
            lcout => \M_this_data_count_q_s_2\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_1\,
            carryout => \M_this_data_count_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_2_THRU_LUT4_0_LC_21_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28981\,
            in2 => \N__30000\,
            in3 => \N__28218\,
            lcout => \M_this_data_count_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_2\,
            carryout => \M_this_data_count_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_3_THRU_LUT4_0_LC_21_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29969\,
            in2 => \N__29047\,
            in3 => \N__28341\,
            lcout => \M_this_data_count_q_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_3\,
            carryout => \M_this_data_count_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_4_THRU_LUT4_0_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28985\,
            in2 => \N__29946\,
            in3 => \N__28338\,
            lcout => \M_this_data_count_q_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_4\,
            carryout => \M_this_data_count_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_5_THRU_LUT4_0_LC_21_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29917\,
            in2 => \N__29048\,
            in3 => \N__28335\,
            lcout => \M_this_data_count_q_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_5\,
            carryout => \M_this_data_count_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_6_THRU_LUT4_0_LC_21_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28989\,
            in2 => \N__31431\,
            in3 => \N__28332\,
            lcout => \M_this_data_count_q_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_6\,
            carryout => \M_this_data_count_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_8_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29003\,
            in2 => \N__29460\,
            in3 => \N__28320\,
            lcout => \M_this_data_count_q_s_8\,
            ltout => OPEN,
            carryin => \bfn_21_23_0_\,
            carryout => \M_this_data_count_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_9_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29496\,
            in2 => \N__29063\,
            in3 => \N__28305\,
            lcout => \M_this_data_count_q_s_9\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_8\,
            carryout => \M_this_data_count_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_9_THRU_LUT4_0_LC_21_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29010\,
            in2 => \N__29526\,
            in3 => \N__28293\,
            lcout => \M_this_data_count_q_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_9\,
            carryout => \M_this_data_count_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_11_LC_21_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29480\,
            in2 => \N__29062\,
            in3 => \N__28281\,
            lcout => \M_this_data_count_q_s_11\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_10\,
            carryout => \M_this_data_count_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_12_LC_21_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29001\,
            in2 => \N__29781\,
            in3 => \N__28269\,
            lcout => \M_this_data_count_q_s_12\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_11\,
            carryout => \M_this_data_count_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_12_THRU_LUT4_0_LC_21_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29820\,
            in2 => \N__29064\,
            in3 => \N__29127\,
            lcout => \M_this_data_count_q_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_12\,
            carryout => \M_this_data_count_q_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_14_LC_21_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29002\,
            in2 => \N__29838\,
            in3 => \N__28569\,
            lcout => \M_this_data_count_q_s_14\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_13\,
            carryout => \M_this_data_count_q_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_15_LC_21_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29799\,
            in2 => \_gnd_net_\,
            in3 => \N__28566\,
            lcout => \M_this_data_count_q_s_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_0_LC_21_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__31356\,
            in1 => \N__28551\,
            in2 => \N__32405\,
            in3 => \N__28527\,
            lcout => \N_226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_6_LC_22_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28401\,
            in2 => \_gnd_net_\,
            in3 => \N__35690\,
            lcout => \M_this_oam_ram_write_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_2_LC_22_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28383\,
            in2 => \_gnd_net_\,
            in3 => \N__35689\,
            lcout => \M_this_oam_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_1_LC_22_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28359\,
            in2 => \_gnd_net_\,
            in3 => \N__35688\,
            lcout => \M_this_oam_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_4_LC_22_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__30066\,
            in1 => \N__33257\,
            in2 => \_gnd_net_\,
            in3 => \N__30770\,
            lcout => \M_this_oam_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36850\,
            ce => 'H',
            sr => \N__32217\
        );

    \M_this_oam_address_q_5_LC_22_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__30771\,
            in1 => \N__30106\,
            in2 => \N__33261\,
            in3 => \N__30067\,
            lcout => \M_this_oam_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36850\,
            ce => 'H',
            sr => \N__32217\
        );

    \this_ppu.un1_oam_data_ac0_1_LC_22_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32098\,
            in2 => \_gnd_net_\,
            in3 => \N__32064\,
            lcout => \this_ppu.un1_oam_data_c2\,
            ltout => \this_ppu.un1_oam_data_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_axbxc3_LC_22_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__29239\,
            in1 => \_gnd_net_\,
            in2 => \N__29268\,
            in3 => \N__32137\,
            lcout => \this_ppu.un1_M_vaddress_q_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_23_LC_22_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29259\,
            in2 => \_gnd_net_\,
            in3 => \N__35627\,
            lcout => \M_this_oam_ram_write_data_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_axbxc4_LC_22_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__29240\,
            in1 => \N__32138\,
            in2 => \N__29213\,
            in3 => \N__29184\,
            lcout => \this_ppu.un1_M_vaddress_q_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_25_LC_22_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33359\,
            in2 => \_gnd_net_\,
            in3 => \N__35626\,
            lcout => \M_this_oam_ram_write_data_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a4_17_LC_22_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__35628\,
            in1 => \_gnd_net_\,
            in2 => \N__29163\,
            in3 => \_gnd_net_\,
            lcout => \M_this_oam_ram_write_data_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_axbxc1_LC_22_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32099\,
            in2 => \_gnd_net_\,
            in3 => \N__32065\,
            lcout => \this_ppu.un1_M_vaddress_q_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_22_LC_22_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34440\,
            lcout => \M_this_data_tmp_qZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36858\,
            ce => \N__34018\,
            sr => \N__36022\
        );

    \M_this_data_tmp_q_esr_21_LC_22_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36252\,
            lcout => \M_this_data_tmp_qZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36858\,
            ce => \N__34018\,
            sr => \N__36022\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_24_LC_22_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31351\,
            in2 => \_gnd_net_\,
            in3 => \N__35625\,
            lcout => \M_this_oam_ram_write_data_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI24IA1_0_1_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__30556\,
            in1 => \N__30669\,
            in2 => \N__30845\,
            in3 => \N__36101\,
            lcout => \N_1404_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI24IA1_1_LC_22_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__30552\,
            in1 => \N__30668\,
            in2 => \N__30852\,
            in3 => \N__36100\,
            lcout => \N_1396_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_1_LC_22_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__30547\,
            in1 => \N__30666\,
            in2 => \N__30855\,
            in3 => \N__33250\,
            lcout => \M_this_oam_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36915\,
            ce => 'H',
            sr => \N__32213\
        );

    \M_this_state_q_12_LC_22_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__33227\,
            in1 => \N__29406\,
            in2 => \N__30854\,
            in3 => \N__30489\,
            lcout => \M_this_state_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36925\,
            ce => 'H',
            sr => \N__36005\
        );

    \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_o2_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30604\,
            in2 => \_gnd_net_\,
            in3 => \N__29375\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_469_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_qlde_i_0_m2_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000010111111"
        )
    port map (
            in0 => \N__31214\,
            in1 => \N__30444\,
            in2 => \N__29340\,
            in3 => \N__31118\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_qlde_i_0_i_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__29727\,
            in1 => \N__36099\,
            in2 => \N__29337\,
            in3 => \N__29330\,
            lcout => \N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_qlde_i_o2_1_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__30280\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31538\,
            lcout => \this_vga_signals.N_461_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNI60TF_15_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29831\,
            in1 => \N__29815\,
            in2 => \N__29798\,
            in3 => \N__29774\,
            lcout => \M_this_state_d62_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_qlde_i_0_a2_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__35164\,
            in1 => \N__36324\,
            in2 => \_gnd_net_\,
            in3 => \N__29761\,
            lcout => \this_vga_signals.M_this_external_address_qlde_i_0_aZ0Z2\,
            ltout => \this_vga_signals.M_this_external_address_qlde_i_0_aZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_qlde_i_i_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011111111"
        )
    port map (
            in0 => \N__29721\,
            in1 => \N__29710\,
            in2 => \N__29610\,
            in3 => \N__29607\,
            lcout => \N_364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIQ9QL_0_LC_22_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29597\,
            in1 => \N__30025\,
            in2 => \N__29999\,
            in3 => \N__29584\,
            lcout => OPEN,
            ltout => \M_this_state_d62_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNII1EE2_10_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29568\,
            in1 => \N__29442\,
            in2 => \N__29559\,
            in3 => \N__29436\,
            lcout => \M_this_state_d62\,
            ltout => \M_this_state_d62_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_716_i_LC_22_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29556\,
            in2 => \N__29529\,
            in3 => \N__36096\,
            lcout => \N_716_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNI8TRI_10_LC_22_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29519\,
            in1 => \N__29492\,
            in2 => \N__29481\,
            in3 => \N__29453\,
            lcout => \M_this_state_d62_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNIAQQL_4_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29919\,
            in1 => \N__29941\,
            in2 => \N__31427\,
            in3 => \N__29968\,
            lcout => \M_this_state_d62_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_1_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__30036\,
            in1 => \N__31489\,
            in2 => \_gnd_net_\,
            in3 => \N__30029\,
            lcout => \M_this_data_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36947\,
            ce => \N__31393\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_3_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000101"
        )
    port map (
            in0 => \N__31490\,
            in1 => \_gnd_net_\,
            in2 => \N__30009\,
            in3 => \N__29998\,
            lcout => \M_this_data_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36947\,
            ce => \N__31393\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_4_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__29976\,
            in1 => \N__31491\,
            in2 => \_gnd_net_\,
            in3 => \N__29970\,
            lcout => \M_this_data_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36947\,
            ce => \N__31393\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_5_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__31492\,
            in1 => \N__29952\,
            in2 => \_gnd_net_\,
            in3 => \N__29945\,
            lcout => \M_this_data_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36947\,
            ce => \N__31393\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_6_LC_22_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__29925\,
            in1 => \N__31493\,
            in2 => \_gnd_net_\,
            in3 => \N__29918\,
            lcout => \M_this_data_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36947\,
            ce => \N__31393\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_4_LC_23_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30249\,
            in2 => \_gnd_net_\,
            in3 => \N__35699\,
            lcout => \M_this_oam_ram_write_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_7_LC_23_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29886\,
            in2 => \_gnd_net_\,
            in3 => \N__35700\,
            lcout => \M_this_oam_ram_write_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a4_8_LC_23_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30867\,
            in2 => \_gnd_net_\,
            in3 => \N__35701\,
            lcout => \M_this_oam_ram_write_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_0_LC_23_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30243\,
            in2 => \_gnd_net_\,
            in3 => \N__35698\,
            lcout => \M_this_oam_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_4_LC_23_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32448\,
            lcout => \M_this_data_tmp_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36855\,
            ce => \N__30237\,
            sr => \N__36026\
        );

    \M_this_data_tmp_q_esr_0_LC_23_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31361\,
            lcout => \M_this_data_tmp_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36855\,
            ce => \N__30237\,
            sr => \N__36026\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_3_LC_23_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35630\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30174\,
            lcout => \M_this_oam_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_10_LC_23_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30138\,
            in2 => \_gnd_net_\,
            in3 => \N__35629\,
            lcout => \M_this_oam_ram_write_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_10_LC_23_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35203\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36867\,
            ce => \N__36143\,
            sr => \N__36021\
        );

    \M_this_data_tmp_q_esr_12_LC_23_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32444\,
            lcout => \M_this_data_tmp_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36867\,
            ce => \N__36143\,
            sr => \N__36021\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a4_11_LC_23_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30042\,
            in2 => \_gnd_net_\,
            in3 => \N__35642\,
            lcout => \M_this_oam_ram_write_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNIOKR51_5_LC_23_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30110\,
            in1 => \N__30077\,
            in2 => \_gnd_net_\,
            in3 => \N__30764\,
            lcout => \un1_M_this_oam_address_q_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_11_LC_23_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35864\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36880\,
            ce => \N__36141\,
            sr => \N__36013\
        );

    \M_this_data_tmp_q_esr_8_LC_23_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31303\,
            lcout => \M_this_data_tmp_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36888\,
            ce => \N__36128\,
            sr => \N__36010\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_0_a2_1_a2_LC_23_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30811\,
            in1 => \N__30557\,
            in2 => \_gnd_net_\,
            in3 => \N__30667\,
            lcout => \M_this_oam_ram_write_data_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNILNG41_3_LC_23_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30727\,
            in1 => \N__30690\,
            in2 => \_gnd_net_\,
            in3 => \N__30505\,
            lcout => \un1_M_this_oam_address_q_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_3_LC_23_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__30507\,
            in1 => \N__30728\,
            in2 => \N__33251\,
            in3 => \N__30692\,
            lcout => \M_this_oam_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36908\,
            ce => 'H',
            sr => \N__32215\
        );

    \M_this_oam_address_q_2_LC_23_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__30691\,
            in1 => \N__33240\,
            in2 => \_gnd_net_\,
            in3 => \N__30506\,
            lcout => \M_this_oam_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36908\,
            ce => 'H',
            sr => \N__32215\
        );

    \M_this_oam_address_q_RNIMU531_1_LC_23_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30665\,
            in1 => \N__30606\,
            in2 => \N__30548\,
            in3 => \N__31106\,
            lcout => \un1_M_this_oam_address_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_7_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__30374\,
            in1 => \N__30481\,
            in2 => \N__30459\,
            in3 => \N__30443\,
            lcout => \M_this_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36938\,
            ce => 'H',
            sr => \N__36006\
        );

    \M_this_state_q_0_LC_23_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101011100000011"
        )
    port map (
            in0 => \N__30327\,
            in1 => \N__30312\,
            in2 => \N__30300\,
            in3 => \N__30284\,
            lcout => led_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36938\,
            ce => 'H',
            sr => \N__36006\
        );

    \this_vga_signals.M_this_external_address_q_3_i_i_14_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__31677\,
            in1 => \N__35038\,
            in2 => \N__34424\,
            in3 => \N__31707\,
            lcout => \N_312_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0_12_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__36284\,
            in1 => \N__31209\,
            in2 => \_gnd_net_\,
            in3 => \N__36093\,
            lcout => \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0Z0Z_12\,
            ltout => \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_3_0_0_12_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__32406\,
            in1 => \N__31671\,
            in2 => \N__31656\,
            in3 => \N__35040\,
            lcout => \M_this_external_address_q_3_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_3L4_LC_23_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__31589\,
            in1 => \N__31562\,
            in2 => \_gnd_net_\,
            in3 => \N__31531\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_3LZ0Z4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_3_i_0_0_15_LC_23_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101010101"
        )
    port map (
            in0 => \N__36094\,
            in1 => \N__34552\,
            in2 => \N__31215\,
            in3 => \N__31119\,
            lcout => \this_vga_signals_M_this_external_address_q_3_i_0_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_7_LC_23_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__31506\,
            in1 => \N__31494\,
            in2 => \_gnd_net_\,
            in3 => \N__31420\,
            lcout => \M_this_data_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36948\,
            ce => \N__31401\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_8_LC_23_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__36495\,
            in1 => \N__37107\,
            in2 => \N__31360\,
            in3 => \N__35035\,
            lcout => \M_this_external_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36951\,
            ce => \N__36561\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_3_0_0_a2_12_LC_23_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31184\,
            in1 => \N__36091\,
            in2 => \_gnd_net_\,
            in3 => \N__31107\,
            lcout => \N_760\,
            ltout => \N_760_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_11_LC_23_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__35839\,
            in1 => \N__37106\,
            in2 => \N__30870\,
            in3 => \N__36372\,
            lcout => \M_this_external_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36951\,
            ce => \N__36561\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_12_LC_23_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010010111110"
        )
    port map (
            in0 => \N__37105\,
            in1 => \N__37317\,
            in2 => \N__37343\,
            in3 => \N__31938\,
            lcout => \M_this_external_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36951\,
            ce => \N__36561\,
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_5_0_wclke_3_LC_23_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__34993\,
            in1 => \N__34910\,
            in2 => \N__34830\,
            in3 => \N__34682\,
            lcout => \this_sprites_ram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_axbxc2_LC_24_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__31737\,
            in1 => \N__31831\,
            in2 => \_gnd_net_\,
            in3 => \N__31797\,
            lcout => \this_ppu.un1_M_haddress_q_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_13_LC_24_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36159\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35705\,
            lcout => \M_this_oam_ram_write_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_15_LC_24_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35706\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34467\,
            lcout => \M_this_oam_ram_write_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_axbxc4_LC_24_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__31763\,
            in1 => \N__31739\,
            in2 => \N__31871\,
            in3 => \N__31776\,
            lcout => \this_ppu.un1_M_haddress_q_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_ac0_1_LC_24_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31830\,
            in2 => \_gnd_net_\,
            in3 => \N__31796\,
            lcout => \this_ppu.un1_oam_data_1_c2\,
            ltout => \this_ppu.un1_oam_data_1_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_axbxc3_LC_24_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31762\,
            in2 => \N__31746\,
            in3 => \N__31738\,
            lcout => \this_ppu.un1_M_haddress_q_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_12_LC_24_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32157\,
            in2 => \_gnd_net_\,
            in3 => \N__35702\,
            lcout => \M_this_oam_ram_write_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_axbxc2_LC_24_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__32128\,
            in1 => \N__32097\,
            in2 => \_gnd_net_\,
            in3 => \N__32063\,
            lcout => \this_ppu.un1_M_vaddress_q_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_5_LC_24_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32022\,
            in2 => \_gnd_net_\,
            in3 => \N__35703\,
            lcout => \M_this_oam_ram_write_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_0_RNISG75_LC_24_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31984\,
            lcout => \M_this_oam_ram_read_data_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a4_9_LC_24_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32166\,
            in2 => \_gnd_net_\,
            in3 => \N__35704\,
            lcout => \M_this_oam_ram_write_data_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_18_LC_24_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32460\,
            in2 => \_gnd_net_\,
            in3 => \N__35695\,
            lcout => \M_this_oam_ram_write_data_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_20_LC_24_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35696\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32454\,
            lcout => \M_this_oam_ram_write_data_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_29_LC_24_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36301\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35692\,
            lcout => \M_this_oam_ram_write_data_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_30_LC_24_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35693\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34417\,
            lcout => \M_this_oam_ram_write_data_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_22_LC_24_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32487\,
            in2 => \_gnd_net_\,
            in3 => \N__35697\,
            lcout => \M_this_oam_ram_write_data_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_31_LC_24_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35694\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34529\,
            lcout => \M_this_oam_ram_write_data_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_18_LC_24_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35234\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36873\,
            ce => \N__34020\,
            sr => \N__36017\
        );

    \M_this_data_tmp_q_esr_20_LC_24_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32442\,
            lcout => \M_this_data_tmp_qZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36873\,
            ce => \N__34020\,
            sr => \N__36017\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_28_LC_24_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32443\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35643\,
            lcout => \M_this_oam_ram_write_data_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_21_LC_24_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35644\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32289\,
            lcout => \M_this_oam_ram_write_data_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_6_LC_24_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__32266\,
            in1 => \N__33245\,
            in2 => \_gnd_net_\,
            in3 => \N__32249\,
            lcout => \M_this_oam_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36881\,
            ce => 'H',
            sr => \N__32216\
        );

    \M_this_oam_address_q_7_LC_24_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__32267\,
            in1 => \N__33246\,
            in2 => \N__32237\,
            in3 => \N__32250\,
            lcout => \M_this_oam_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36881\,
            ce => 'H',
            sr => \N__32216\
        );

    \M_this_data_tmp_q_esr_9_LC_24_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33371\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36889\,
            ce => \N__36142\,
            sr => \N__36011\
        );

    \this_ppu.un2_hscroll_cry_0_c_inv_LC_24_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33153\,
            in2 => \N__34307\,
            in3 => \N__32793\,
            lcout => \this_ppu.M_this_oam_ram_read_data_iZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_24_11_0_\,
            carryout => \this_ppu.un2_hscroll_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_24_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33147\,
            in2 => \N__33066\,
            in3 => \N__33138\,
            lcout => \this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un2_hscroll_cry_0\,
            carryout => \this_ppu.un2_hscroll_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_24_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__33131\,
            in1 => \N__32739\,
            in2 => \_gnd_net_\,
            in3 => \N__33093\,
            lcout => \this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_26_LC_24_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35168\,
            in2 => \_gnd_net_\,
            in3 => \N__35540\,
            lcout => \M_this_oam_ram_write_data_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a4_19_LC_24_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35541\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34029\,
            lcout => \M_this_oam_ram_write_data_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI0O061_1_LC_24_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__33790\,
            in1 => \N__33064\,
            in2 => \N__33933\,
            in3 => \N__32994\,
            lcout => \M_this_ppu_sprites_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI88B5_0_LC_24_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__32794\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34301\,
            lcout => \this_ppu.un2_hscroll_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI3S161_2_LC_24_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__33775\,
            in1 => \N__33917\,
            in2 => \N__32747\,
            in3 => \N__32670\,
            lcout => \M_this_ppu_sprites_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNIRG7O_0_LC_24_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000001"
        )
    port map (
            in0 => \N__34320\,
            in1 => \N__33774\,
            in2 => \N__33932\,
            in3 => \N__34302\,
            lcout => \M_this_ppu_sprites_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_19_LC_24_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35848\,
            lcout => \M_this_data_tmp_qZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36916\,
            ce => \N__34005\,
            sr => \N__36007\
        );

    \this_ppu.M_state_q_RNI0VTU_2_4_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__33975\,
            in1 => \N__33960\,
            in2 => \N__33931\,
            in3 => \N__33791\,
            lcout => \M_this_ppu_sprites_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34996\,
            in1 => \N__34905\,
            in2 => \N__34832\,
            in3 => \N__34709\,
            lcout => \this_sprites_ram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__34710\,
            in1 => \N__34821\,
            in2 => \N__34913\,
            in3 => \N__34997\,
            lcout => \this_sprites_ram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__34998\,
            in1 => \N__34889\,
            in2 => \N__34833\,
            in3 => \N__34708\,
            lcout => \this_sprites_ram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_9_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__35039\,
            in1 => \N__36453\,
            in2 => \N__33400\,
            in3 => \N__37116\,
            lcout => \M_this_external_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36944\,
            ce => \N__36560\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_15_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__37115\,
            in1 => \N__33267\,
            in2 => \N__37176\,
            in3 => \N__33244\,
            lcout => \M_this_external_address_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36944\,
            ce => \N__36560\,
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__34906\,
            in1 => \N__34991\,
            in2 => \N__34828\,
            in3 => \N__34693\,
            lcout => \this_sprites_ram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_external_address_q_3_0_0_13_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__36259\,
            in1 => \N__35037\,
            in2 => \_gnd_net_\,
            in3 => \N__35361\,
            lcout => \M_this_external_address_q_3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_4L6_LC_24_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35285\,
            in1 => \N__35270\,
            in2 => \N__35307\,
            in3 => \N__35352\,
            lcout => \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_4LZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_19_i_0_o2_4_LC_24_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35327\,
            in1 => \N__35306\,
            in2 => \N__35289\,
            in3 => \N__35271\,
            lcout => \this_vga_signals.un1_M_this_state_q_19_i_0_o2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_10_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37114\,
            in1 => \N__36411\,
            in2 => \N__35172\,
            in3 => \N__35036\,
            lcout => \M_this_external_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36954\,
            ce => \N__36576\,
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__34992\,
            in1 => \N__34911\,
            in2 => \N__34829\,
            in3 => \N__34683\,
            lcout => \this_sprites_ram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_14_LC_26_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34329\,
            in2 => \_gnd_net_\,
            in3 => \N__35691\,
            lcout => \M_this_oam_ram_write_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_15_LC_26_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34513\,
            lcout => \M_this_data_tmp_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36882\,
            ce => \N__36147\,
            sr => \N__36014\
        );

    \M_this_data_tmp_q_esr_14_LC_26_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34391\,
            lcout => \M_this_data_tmp_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36882\,
            ce => \N__36147\,
            sr => \N__36014\
        );

    \M_this_data_tmp_q_esr_13_LC_26_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36300\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36882\,
            ce => \N__36147\,
            sr => \N__36014\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_27_LC_26_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35838\,
            in2 => \_gnd_net_\,
            in3 => \N__35641\,
            lcout => \M_this_oam_ram_write_data_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_13_LC_26_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010010111110"
        )
    port map (
            in0 => \N__37113\,
            in1 => \N__37272\,
            in2 => \N__37298\,
            in3 => \N__35502\,
            lcout => \M_this_external_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36957\,
            ce => \N__36574\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_14_LC_26_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010010111110"
        )
    port map (
            in0 => \N__37112\,
            in1 => \N__37227\,
            in2 => \N__37253\,
            in3 => \N__35493\,
            lcout => \M_this_external_address_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36957\,
            ce => \N__36574\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_0_LC_26_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37108\,
            in1 => \N__35471\,
            in2 => \_gnd_net_\,
            in3 => \N__35460\,
            lcout => \M_this_external_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_26_21_0_\,
            carryout => \M_this_external_address_q_cry_0\,
            clk => \N__36958\,
            ce => \N__36575\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_1_LC_26_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37079\,
            in1 => \N__35450\,
            in2 => \_gnd_net_\,
            in3 => \N__35439\,
            lcout => \M_this_external_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_0\,
            carryout => \M_this_external_address_q_cry_1\,
            clk => \N__36958\,
            ce => \N__36575\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_2_LC_26_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37109\,
            in1 => \N__35423\,
            in2 => \_gnd_net_\,
            in3 => \N__35412\,
            lcout => \M_this_external_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_1\,
            carryout => \M_this_external_address_q_cry_2\,
            clk => \N__36958\,
            ce => \N__36575\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_3_LC_26_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37080\,
            in1 => \N__35396\,
            in2 => \_gnd_net_\,
            in3 => \N__35385\,
            lcout => \M_this_external_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_2\,
            carryout => \M_this_external_address_q_cry_3\,
            clk => \N__36958\,
            ce => \N__36575\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_4_LC_26_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37110\,
            in1 => \N__35372\,
            in2 => \_gnd_net_\,
            in3 => \N__37161\,
            lcout => \M_this_external_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_3\,
            carryout => \M_this_external_address_q_cry_4\,
            clk => \N__36958\,
            ce => \N__36575\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_5_LC_26_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37081\,
            in1 => \N__37154\,
            in2 => \_gnd_net_\,
            in3 => \N__37143\,
            lcout => \M_this_external_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_4\,
            carryout => \M_this_external_address_q_cry_5\,
            clk => \N__36958\,
            ce => \N__36575\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_6_LC_26_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37111\,
            in1 => \N__37130\,
            in2 => \_gnd_net_\,
            in3 => \N__37119\,
            lcout => \M_this_external_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_5\,
            carryout => \M_this_external_address_q_cry_6\,
            clk => \N__36958\,
            ce => \N__36575\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_7_LC_26_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37082\,
            in1 => \N__36992\,
            in2 => \_gnd_net_\,
            in3 => \N__36981\,
            lcout => \M_this_external_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_6\,
            carryout => \M_this_external_address_q_cry_7\,
            clk => \N__36958\,
            ce => \N__36575\,
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_RNO_0_8_LC_26_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36512\,
            in2 => \_gnd_net_\,
            in3 => \N__36486\,
            lcout => \M_this_external_address_q_s_8\,
            ltout => OPEN,
            carryin => \bfn_26_22_0_\,
            carryout => \M_this_external_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_RNO_0_9_LC_26_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36476\,
            in2 => \_gnd_net_\,
            in3 => \N__36441\,
            lcout => \M_this_external_address_q_s_9\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_8\,
            carryout => \M_this_external_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_RNO_0_10_LC_26_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36428\,
            in2 => \_gnd_net_\,
            in3 => \N__36402\,
            lcout => \M_this_external_address_q_s_10\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_9\,
            carryout => \M_this_external_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_RNO_0_11_LC_26_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36386\,
            in2 => \_gnd_net_\,
            in3 => \N__36363\,
            lcout => \M_this_external_address_q_s_11\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_10\,
            carryout => \M_this_external_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_cry_11_THRU_LUT4_0_LC_26_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37342\,
            in2 => \_gnd_net_\,
            in3 => \N__37308\,
            lcout => \M_this_external_address_q_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_11\,
            carryout => \M_this_external_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_cry_12_THRU_LUT4_0_LC_26_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37297\,
            in2 => \_gnd_net_\,
            in3 => \N__37263\,
            lcout => \M_this_external_address_q_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_12\,
            carryout => \M_this_external_address_q_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_cry_13_THRU_LUT4_0_LC_26_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37252\,
            in2 => \_gnd_net_\,
            in3 => \N__37218\,
            lcout => \M_this_external_address_q_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_external_address_q_cry_13\,
            carryout => \M_this_external_address_q_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_RNO_0_15_LC_26_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37202\,
            in2 => \_gnd_net_\,
            in3 => \N__37179\,
            lcout => \M_this_external_address_q_s_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
