// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     May 10 2022 20:23:05

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    debug,
    rgb,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    clk);

    inout [15:0] port_address;
    input [7:0] port_data;
    output [1:0] debug;
    output [5:0] rgb;
    output vsync;
    output vblank;
    input rst_n;
    inout port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    input clk;

    wire N__22316;
    wire N__22315;
    wire N__22314;
    wire N__22305;
    wire N__22304;
    wire N__22303;
    wire N__22296;
    wire N__22295;
    wire N__22294;
    wire N__22287;
    wire N__22286;
    wire N__22285;
    wire N__22278;
    wire N__22277;
    wire N__22276;
    wire N__22269;
    wire N__22268;
    wire N__22267;
    wire N__22260;
    wire N__22259;
    wire N__22258;
    wire N__22251;
    wire N__22250;
    wire N__22249;
    wire N__22242;
    wire N__22241;
    wire N__22240;
    wire N__22233;
    wire N__22232;
    wire N__22231;
    wire N__22224;
    wire N__22223;
    wire N__22222;
    wire N__22215;
    wire N__22214;
    wire N__22213;
    wire N__22206;
    wire N__22205;
    wire N__22204;
    wire N__22197;
    wire N__22196;
    wire N__22195;
    wire N__22188;
    wire N__22187;
    wire N__22186;
    wire N__22179;
    wire N__22178;
    wire N__22177;
    wire N__22170;
    wire N__22169;
    wire N__22168;
    wire N__22161;
    wire N__22160;
    wire N__22159;
    wire N__22152;
    wire N__22151;
    wire N__22150;
    wire N__22143;
    wire N__22142;
    wire N__22141;
    wire N__22134;
    wire N__22133;
    wire N__22132;
    wire N__22125;
    wire N__22124;
    wire N__22123;
    wire N__22116;
    wire N__22115;
    wire N__22114;
    wire N__22107;
    wire N__22106;
    wire N__22105;
    wire N__22098;
    wire N__22097;
    wire N__22096;
    wire N__22089;
    wire N__22088;
    wire N__22087;
    wire N__22080;
    wire N__22079;
    wire N__22078;
    wire N__22071;
    wire N__22070;
    wire N__22069;
    wire N__22062;
    wire N__22061;
    wire N__22060;
    wire N__22053;
    wire N__22052;
    wire N__22051;
    wire N__22044;
    wire N__22043;
    wire N__22042;
    wire N__22035;
    wire N__22034;
    wire N__22033;
    wire N__22026;
    wire N__22025;
    wire N__22024;
    wire N__22017;
    wire N__22016;
    wire N__22015;
    wire N__22008;
    wire N__22007;
    wire N__22006;
    wire N__21999;
    wire N__21998;
    wire N__21997;
    wire N__21990;
    wire N__21989;
    wire N__21988;
    wire N__21981;
    wire N__21980;
    wire N__21979;
    wire N__21972;
    wire N__21971;
    wire N__21970;
    wire N__21963;
    wire N__21962;
    wire N__21961;
    wire N__21954;
    wire N__21953;
    wire N__21952;
    wire N__21945;
    wire N__21944;
    wire N__21943;
    wire N__21936;
    wire N__21935;
    wire N__21934;
    wire N__21927;
    wire N__21926;
    wire N__21925;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21898;
    wire N__21895;
    wire N__21892;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21863;
    wire N__21860;
    wire N__21859;
    wire N__21858;
    wire N__21857;
    wire N__21856;
    wire N__21855;
    wire N__21854;
    wire N__21853;
    wire N__21852;
    wire N__21851;
    wire N__21850;
    wire N__21849;
    wire N__21848;
    wire N__21847;
    wire N__21846;
    wire N__21845;
    wire N__21844;
    wire N__21843;
    wire N__21842;
    wire N__21841;
    wire N__21840;
    wire N__21839;
    wire N__21838;
    wire N__21837;
    wire N__21836;
    wire N__21835;
    wire N__21830;
    wire N__21821;
    wire N__21820;
    wire N__21819;
    wire N__21810;
    wire N__21801;
    wire N__21792;
    wire N__21783;
    wire N__21782;
    wire N__21775;
    wire N__21772;
    wire N__21767;
    wire N__21762;
    wire N__21761;
    wire N__21758;
    wire N__21751;
    wire N__21748;
    wire N__21747;
    wire N__21746;
    wire N__21743;
    wire N__21736;
    wire N__21733;
    wire N__21728;
    wire N__21727;
    wire N__21724;
    wire N__21719;
    wire N__21718;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21706;
    wire N__21703;
    wire N__21698;
    wire N__21693;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21653;
    wire N__21652;
    wire N__21651;
    wire N__21650;
    wire N__21649;
    wire N__21648;
    wire N__21647;
    wire N__21646;
    wire N__21645;
    wire N__21644;
    wire N__21643;
    wire N__21642;
    wire N__21641;
    wire N__21640;
    wire N__21639;
    wire N__21638;
    wire N__21637;
    wire N__21636;
    wire N__21635;
    wire N__21634;
    wire N__21633;
    wire N__21632;
    wire N__21631;
    wire N__21630;
    wire N__21629;
    wire N__21628;
    wire N__21627;
    wire N__21626;
    wire N__21625;
    wire N__21624;
    wire N__21623;
    wire N__21622;
    wire N__21621;
    wire N__21620;
    wire N__21619;
    wire N__21618;
    wire N__21617;
    wire N__21616;
    wire N__21615;
    wire N__21614;
    wire N__21613;
    wire N__21612;
    wire N__21611;
    wire N__21610;
    wire N__21609;
    wire N__21608;
    wire N__21607;
    wire N__21606;
    wire N__21605;
    wire N__21604;
    wire N__21603;
    wire N__21602;
    wire N__21601;
    wire N__21600;
    wire N__21599;
    wire N__21598;
    wire N__21597;
    wire N__21596;
    wire N__21595;
    wire N__21594;
    wire N__21593;
    wire N__21592;
    wire N__21591;
    wire N__21590;
    wire N__21589;
    wire N__21588;
    wire N__21587;
    wire N__21586;
    wire N__21585;
    wire N__21584;
    wire N__21583;
    wire N__21582;
    wire N__21581;
    wire N__21580;
    wire N__21579;
    wire N__21578;
    wire N__21577;
    wire N__21576;
    wire N__21575;
    wire N__21574;
    wire N__21573;
    wire N__21572;
    wire N__21571;
    wire N__21570;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21394;
    wire N__21393;
    wire N__21392;
    wire N__21391;
    wire N__21390;
    wire N__21389;
    wire N__21388;
    wire N__21387;
    wire N__21386;
    wire N__21385;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21359;
    wire N__21354;
    wire N__21351;
    wire N__21350;
    wire N__21349;
    wire N__21348;
    wire N__21347;
    wire N__21346;
    wire N__21345;
    wire N__21344;
    wire N__21343;
    wire N__21342;
    wire N__21341;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21205;
    wire N__21202;
    wire N__21201;
    wire N__21198;
    wire N__21197;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21118;
    wire N__21115;
    wire N__21112;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21065;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21034;
    wire N__21031;
    wire N__21028;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21016;
    wire N__21013;
    wire N__21010;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20998;
    wire N__20995;
    wire N__20992;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20977;
    wire N__20974;
    wire N__20971;
    wire N__20970;
    wire N__20967;
    wire N__20964;
    wire N__20961;
    wire N__20958;
    wire N__20953;
    wire N__20950;
    wire N__20947;
    wire N__20942;
    wire N__20939;
    wire N__20938;
    wire N__20935;
    wire N__20932;
    wire N__20929;
    wire N__20926;
    wire N__20921;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20902;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20879;
    wire N__20878;
    wire N__20877;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20855;
    wire N__20852;
    wire N__20851;
    wire N__20848;
    wire N__20845;
    wire N__20844;
    wire N__20843;
    wire N__20838;
    wire N__20835;
    wire N__20834;
    wire N__20831;
    wire N__20830;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20815;
    wire N__20810;
    wire N__20805;
    wire N__20802;
    wire N__20801;
    wire N__20798;
    wire N__20793;
    wire N__20790;
    wire N__20783;
    wire N__20782;
    wire N__20779;
    wire N__20776;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20761;
    wire N__20760;
    wire N__20759;
    wire N__20752;
    wire N__20751;
    wire N__20750;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20735;
    wire N__20734;
    wire N__20731;
    wire N__20730;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20712;
    wire N__20707;
    wire N__20704;
    wire N__20699;
    wire N__20696;
    wire N__20687;
    wire N__20686;
    wire N__20685;
    wire N__20682;
    wire N__20681;
    wire N__20680;
    wire N__20679;
    wire N__20676;
    wire N__20675;
    wire N__20672;
    wire N__20665;
    wire N__20664;
    wire N__20663;
    wire N__20660;
    wire N__20655;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20609;
    wire N__20606;
    wire N__20597;
    wire N__20596;
    wire N__20595;
    wire N__20594;
    wire N__20591;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20567;
    wire N__20566;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20554;
    wire N__20551;
    wire N__20550;
    wire N__20543;
    wire N__20538;
    wire N__20535;
    wire N__20530;
    wire N__20527;
    wire N__20526;
    wire N__20521;
    wire N__20518;
    wire N__20513;
    wire N__20512;
    wire N__20511;
    wire N__20510;
    wire N__20503;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20493;
    wire N__20490;
    wire N__20489;
    wire N__20488;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20470;
    wire N__20459;
    wire N__20456;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20437;
    wire N__20436;
    wire N__20435;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20427;
    wire N__20424;
    wire N__20421;
    wire N__20420;
    wire N__20419;
    wire N__20416;
    wire N__20415;
    wire N__20414;
    wire N__20409;
    wire N__20406;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20394;
    wire N__20393;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20382;
    wire N__20381;
    wire N__20376;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20362;
    wire N__20361;
    wire N__20360;
    wire N__20357;
    wire N__20356;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20344;
    wire N__20343;
    wire N__20340;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20324;
    wire N__20323;
    wire N__20322;
    wire N__20319;
    wire N__20318;
    wire N__20317;
    wire N__20316;
    wire N__20313;
    wire N__20312;
    wire N__20309;
    wire N__20308;
    wire N__20307;
    wire N__20306;
    wire N__20305;
    wire N__20298;
    wire N__20295;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20272;
    wire N__20271;
    wire N__20268;
    wire N__20267;
    wire N__20264;
    wire N__20263;
    wire N__20260;
    wire N__20259;
    wire N__20256;
    wire N__20255;
    wire N__20252;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20234;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20207;
    wire N__20204;
    wire N__20189;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20181;
    wire N__20180;
    wire N__20175;
    wire N__20170;
    wire N__20167;
    wire N__20162;
    wire N__20153;
    wire N__20150;
    wire N__20149;
    wire N__20144;
    wire N__20141;
    wire N__20136;
    wire N__20135;
    wire N__20132;
    wire N__20131;
    wire N__20128;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20103;
    wire N__20096;
    wire N__20093;
    wire N__20088;
    wire N__20083;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20060;
    wire N__20059;
    wire N__20056;
    wire N__20055;
    wire N__20054;
    wire N__20053;
    wire N__20052;
    wire N__20051;
    wire N__20050;
    wire N__20049;
    wire N__20048;
    wire N__20047;
    wire N__20044;
    wire N__20041;
    wire N__20040;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20023;
    wire N__20020;
    wire N__20019;
    wire N__20016;
    wire N__20015;
    wire N__20012;
    wire N__20011;
    wire N__20008;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19996;
    wire N__19995;
    wire N__19990;
    wire N__19983;
    wire N__19966;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19956;
    wire N__19951;
    wire N__19944;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19932;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19911;
    wire N__19908;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19813;
    wire N__19810;
    wire N__19807;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19627;
    wire N__19626;
    wire N__19625;
    wire N__19624;
    wire N__19623;
    wire N__19622;
    wire N__19621;
    wire N__19620;
    wire N__19619;
    wire N__19618;
    wire N__19617;
    wire N__19616;
    wire N__19615;
    wire N__19612;
    wire N__19601;
    wire N__19598;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19580;
    wire N__19571;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19431;
    wire N__19430;
    wire N__19425;
    wire N__19422;
    wire N__19421;
    wire N__19418;
    wire N__19417;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19402;
    wire N__19397;
    wire N__19392;
    wire N__19389;
    wire N__19388;
    wire N__19385;
    wire N__19380;
    wire N__19377;
    wire N__19370;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19213;
    wire N__19212;
    wire N__19211;
    wire N__19210;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19199;
    wire N__19196;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19165;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19054;
    wire N__19053;
    wire N__19048;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19031;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19023;
    wire N__19020;
    wire N__19019;
    wire N__19016;
    wire N__19015;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19005;
    wire N__19002;
    wire N__18999;
    wire N__18996;
    wire N__18989;
    wire N__18980;
    wire N__18979;
    wire N__18976;
    wire N__18975;
    wire N__18972;
    wire N__18969;
    wire N__18966;
    wire N__18963;
    wire N__18960;
    wire N__18957;
    wire N__18952;
    wire N__18949;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18937;
    wire N__18934;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18912;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18895;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18866;
    wire N__18865;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18853;
    wire N__18850;
    wire N__18849;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18831;
    wire N__18826;
    wire N__18823;
    wire N__18818;
    wire N__18815;
    wire N__18810;
    wire N__18805;
    wire N__18800;
    wire N__18799;
    wire N__18798;
    wire N__18797;
    wire N__18796;
    wire N__18795;
    wire N__18794;
    wire N__18793;
    wire N__18792;
    wire N__18791;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18772;
    wire N__18771;
    wire N__18764;
    wire N__18763;
    wire N__18762;
    wire N__18761;
    wire N__18756;
    wire N__18751;
    wire N__18748;
    wire N__18741;
    wire N__18740;
    wire N__18739;
    wire N__18738;
    wire N__18737;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18725;
    wire N__18722;
    wire N__18717;
    wire N__18712;
    wire N__18709;
    wire N__18700;
    wire N__18683;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18661;
    wire N__18658;
    wire N__18655;
    wire N__18650;
    wire N__18647;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18623;
    wire N__18622;
    wire N__18619;
    wire N__18616;
    wire N__18613;
    wire N__18610;
    wire N__18605;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18574;
    wire N__18571;
    wire N__18568;
    wire N__18565;
    wire N__18562;
    wire N__18559;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18547;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18466;
    wire N__18463;
    wire N__18462;
    wire N__18461;
    wire N__18460;
    wire N__18459;
    wire N__18456;
    wire N__18451;
    wire N__18444;
    wire N__18441;
    wire N__18436;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18418;
    wire N__18417;
    wire N__18414;
    wire N__18413;
    wire N__18412;
    wire N__18409;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18393;
    wire N__18390;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18376;
    wire N__18373;
    wire N__18370;
    wire N__18365;
    wire N__18364;
    wire N__18363;
    wire N__18360;
    wire N__18359;
    wire N__18356;
    wire N__18355;
    wire N__18352;
    wire N__18351;
    wire N__18350;
    wire N__18347;
    wire N__18340;
    wire N__18337;
    wire N__18332;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18310;
    wire N__18309;
    wire N__18308;
    wire N__18307;
    wire N__18306;
    wire N__18303;
    wire N__18296;
    wire N__18291;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18274;
    wire N__18271;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18249;
    wire N__18244;
    wire N__18241;
    wire N__18238;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18219;
    wire N__18216;
    wire N__18213;
    wire N__18210;
    wire N__18205;
    wire N__18202;
    wire N__18199;
    wire N__18196;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18184;
    wire N__18181;
    wire N__18180;
    wire N__18177;
    wire N__18176;
    wire N__18175;
    wire N__18172;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18137;
    wire N__18132;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18102;
    wire N__18093;
    wire N__18086;
    wire N__18085;
    wire N__18084;
    wire N__18083;
    wire N__18082;
    wire N__18081;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18073;
    wire N__18070;
    wire N__18069;
    wire N__18066;
    wire N__18063;
    wire N__18060;
    wire N__18057;
    wire N__18052;
    wire N__18051;
    wire N__18050;
    wire N__18047;
    wire N__18046;
    wire N__18045;
    wire N__18042;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18014;
    wire N__18013;
    wire N__18008;
    wire N__18001;
    wire N__17998;
    wire N__17995;
    wire N__17992;
    wire N__17989;
    wire N__17986;
    wire N__17981;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17926;
    wire N__17925;
    wire N__17924;
    wire N__17923;
    wire N__17922;
    wire N__17915;
    wire N__17912;
    wire N__17907;
    wire N__17904;
    wire N__17899;
    wire N__17896;
    wire N__17893;
    wire N__17890;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17777;
    wire N__17776;
    wire N__17775;
    wire N__17772;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17749;
    wire N__17748;
    wire N__17747;
    wire N__17746;
    wire N__17745;
    wire N__17742;
    wire N__17741;
    wire N__17738;
    wire N__17737;
    wire N__17736;
    wire N__17735;
    wire N__17734;
    wire N__17727;
    wire N__17726;
    wire N__17723;
    wire N__17722;
    wire N__17721;
    wire N__17720;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17700;
    wire N__17697;
    wire N__17694;
    wire N__17691;
    wire N__17688;
    wire N__17685;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17666;
    wire N__17661;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17539;
    wire N__17538;
    wire N__17535;
    wire N__17532;
    wire N__17529;
    wire N__17526;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17491;
    wire N__17490;
    wire N__17489;
    wire N__17480;
    wire N__17477;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17363;
    wire N__17360;
    wire N__17357;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17249;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17201;
    wire N__17198;
    wire N__17197;
    wire N__17196;
    wire N__17193;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17177;
    wire N__17174;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17153;
    wire N__17150;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17135;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17096;
    wire N__17093;
    wire N__17090;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17078;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17063;
    wire N__17060;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17035;
    wire N__17032;
    wire N__17031;
    wire N__17028;
    wire N__17025;
    wire N__17022;
    wire N__17017;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16897;
    wire N__16896;
    wire N__16893;
    wire N__16890;
    wire N__16887;
    wire N__16884;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16765;
    wire N__16764;
    wire N__16761;
    wire N__16758;
    wire N__16755;
    wire N__16752;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16633;
    wire N__16632;
    wire N__16629;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16565;
    wire N__16562;
    wire N__16559;
    wire N__16556;
    wire N__16553;
    wire N__16550;
    wire N__16547;
    wire N__16544;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16498;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16406;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16376;
    wire N__16373;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16346;
    wire N__16343;
    wire N__16340;
    wire N__16337;
    wire N__16334;
    wire N__16331;
    wire N__16328;
    wire N__16325;
    wire N__16322;
    wire N__16319;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16307;
    wire N__16304;
    wire N__16303;
    wire N__16300;
    wire N__16297;
    wire N__16294;
    wire N__16291;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16281;
    wire N__16278;
    wire N__16271;
    wire N__16268;
    wire N__16265;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16253;
    wire N__16250;
    wire N__16247;
    wire N__16244;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16226;
    wire N__16223;
    wire N__16220;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16205;
    wire N__16202;
    wire N__16199;
    wire N__16196;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16181;
    wire N__16178;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16163;
    wire N__16160;
    wire N__16157;
    wire N__16154;
    wire N__16153;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16143;
    wire N__16140;
    wire N__16133;
    wire N__16130;
    wire N__16127;
    wire N__16124;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16105;
    wire N__16102;
    wire N__16099;
    wire N__16094;
    wire N__16093;
    wire N__16092;
    wire N__16087;
    wire N__16084;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16055;
    wire N__16054;
    wire N__16053;
    wire N__16052;
    wire N__16049;
    wire N__16046;
    wire N__16041;
    wire N__16036;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16024;
    wire N__16023;
    wire N__16022;
    wire N__16017;
    wire N__16012;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15994;
    wire N__15991;
    wire N__15988;
    wire N__15983;
    wire N__15980;
    wire N__15979;
    wire N__15978;
    wire N__15977;
    wire N__15976;
    wire N__15975;
    wire N__15972;
    wire N__15967;
    wire N__15964;
    wire N__15959;
    wire N__15956;
    wire N__15947;
    wire N__15946;
    wire N__15945;
    wire N__15942;
    wire N__15939;
    wire N__15936;
    wire N__15933;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15907;
    wire N__15904;
    wire N__15901;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15877;
    wire N__15876;
    wire N__15875;
    wire N__15866;
    wire N__15863;
    wire N__15860;
    wire N__15857;
    wire N__15854;
    wire N__15853;
    wire N__15852;
    wire N__15851;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15835;
    wire N__15834;
    wire N__15827;
    wire N__15824;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15803;
    wire N__15800;
    wire N__15799;
    wire N__15798;
    wire N__15797;
    wire N__15788;
    wire N__15785;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15766;
    wire N__15763;
    wire N__15760;
    wire N__15757;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15725;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15701;
    wire N__15698;
    wire N__15697;
    wire N__15694;
    wire N__15691;
    wire N__15686;
    wire N__15685;
    wire N__15682;
    wire N__15679;
    wire N__15676;
    wire N__15671;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15659;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15641;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15617;
    wire N__15616;
    wire N__15615;
    wire N__15612;
    wire N__15607;
    wire N__15602;
    wire N__15601;
    wire N__15598;
    wire N__15595;
    wire N__15590;
    wire N__15587;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15575;
    wire N__15574;
    wire N__15571;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15557;
    wire N__15556;
    wire N__15553;
    wire N__15550;
    wire N__15545;
    wire N__15542;
    wire N__15539;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15527;
    wire N__15526;
    wire N__15523;
    wire N__15520;
    wire N__15515;
    wire N__15514;
    wire N__15511;
    wire N__15508;
    wire N__15505;
    wire N__15500;
    wire N__15499;
    wire N__15496;
    wire N__15493;
    wire N__15488;
    wire N__15485;
    wire N__15482;
    wire N__15479;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15467;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15457;
    wire N__15456;
    wire N__15453;
    wire N__15448;
    wire N__15447;
    wire N__15446;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15436;
    wire N__15435;
    wire N__15432;
    wire N__15429;
    wire N__15422;
    wire N__15419;
    wire N__15410;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15400;
    wire N__15397;
    wire N__15392;
    wire N__15391;
    wire N__15388;
    wire N__15385;
    wire N__15384;
    wire N__15383;
    wire N__15382;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15344;
    wire N__15341;
    wire N__15340;
    wire N__15337;
    wire N__15334;
    wire N__15329;
    wire N__15328;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15317;
    wire N__15316;
    wire N__15313;
    wire N__15308;
    wire N__15307;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15299;
    wire N__15296;
    wire N__15293;
    wire N__15292;
    wire N__15289;
    wire N__15286;
    wire N__15283;
    wire N__15280;
    wire N__15277;
    wire N__15272;
    wire N__15269;
    wire N__15268;
    wire N__15265;
    wire N__15262;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15232;
    wire N__15227;
    wire N__15218;
    wire N__15217;
    wire N__15216;
    wire N__15215;
    wire N__15212;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15204;
    wire N__15201;
    wire N__15198;
    wire N__15197;
    wire N__15194;
    wire N__15193;
    wire N__15190;
    wire N__15187;
    wire N__15184;
    wire N__15183;
    wire N__15180;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15162;
    wire N__15159;
    wire N__15156;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15144;
    wire N__15139;
    wire N__15132;
    wire N__15127;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15115;
    wire N__15112;
    wire N__15109;
    wire N__15098;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15088;
    wire N__15083;
    wire N__15082;
    wire N__15079;
    wire N__15074;
    wire N__15073;
    wire N__15072;
    wire N__15071;
    wire N__15070;
    wire N__15069;
    wire N__15068;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15052;
    wire N__15051;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15037;
    wire N__15034;
    wire N__15029;
    wire N__15024;
    wire N__15021;
    wire N__15018;
    wire N__15011;
    wire N__15008;
    wire N__15007;
    wire N__15004;
    wire N__15003;
    wire N__15000;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14990;
    wire N__14985;
    wire N__14982;
    wire N__14979;
    wire N__14976;
    wire N__14971;
    wire N__14966;
    wire N__14965;
    wire N__14962;
    wire N__14959;
    wire N__14958;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14937;
    wire N__14936;
    wire N__14933;
    wire N__14932;
    wire N__14931;
    wire N__14928;
    wire N__14925;
    wire N__14922;
    wire N__14919;
    wire N__14916;
    wire N__14913;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14878;
    wire N__14875;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14852;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14815;
    wire N__14814;
    wire N__14813;
    wire N__14812;
    wire N__14809;
    wire N__14806;
    wire N__14803;
    wire N__14802;
    wire N__14801;
    wire N__14800;
    wire N__14799;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14791;
    wire N__14790;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14770;
    wire N__14767;
    wire N__14762;
    wire N__14759;
    wire N__14758;
    wire N__14755;
    wire N__14754;
    wire N__14753;
    wire N__14752;
    wire N__14751;
    wire N__14750;
    wire N__14747;
    wire N__14746;
    wire N__14745;
    wire N__14742;
    wire N__14741;
    wire N__14740;
    wire N__14735;
    wire N__14726;
    wire N__14723;
    wire N__14718;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14700;
    wire N__14695;
    wire N__14692;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14672;
    wire N__14667;
    wire N__14664;
    wire N__14653;
    wire N__14644;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14611;
    wire N__14610;
    wire N__14609;
    wire N__14608;
    wire N__14607;
    wire N__14606;
    wire N__14603;
    wire N__14602;
    wire N__14595;
    wire N__14592;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14578;
    wire N__14577;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14565;
    wire N__14564;
    wire N__14561;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14535;
    wire N__14534;
    wire N__14533;
    wire N__14532;
    wire N__14531;
    wire N__14530;
    wire N__14525;
    wire N__14520;
    wire N__14511;
    wire N__14506;
    wire N__14501;
    wire N__14496;
    wire N__14483;
    wire N__14482;
    wire N__14481;
    wire N__14480;
    wire N__14479;
    wire N__14478;
    wire N__14477;
    wire N__14476;
    wire N__14473;
    wire N__14472;
    wire N__14471;
    wire N__14470;
    wire N__14467;
    wire N__14464;
    wire N__14463;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14449;
    wire N__14444;
    wire N__14441;
    wire N__14438;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14423;
    wire N__14418;
    wire N__14415;
    wire N__14412;
    wire N__14409;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14398;
    wire N__14397;
    wire N__14394;
    wire N__14391;
    wire N__14388;
    wire N__14385;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14356;
    wire N__14353;
    wire N__14348;
    wire N__14341;
    wire N__14336;
    wire N__14331;
    wire N__14324;
    wire N__14319;
    wire N__14314;
    wire N__14303;
    wire N__14302;
    wire N__14299;
    wire N__14298;
    wire N__14297;
    wire N__14296;
    wire N__14293;
    wire N__14292;
    wire N__14287;
    wire N__14284;
    wire N__14283;
    wire N__14280;
    wire N__14279;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14271;
    wire N__14268;
    wire N__14267;
    wire N__14266;
    wire N__14265;
    wire N__14264;
    wire N__14263;
    wire N__14260;
    wire N__14259;
    wire N__14258;
    wire N__14255;
    wire N__14252;
    wire N__14249;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14220;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14205;
    wire N__14200;
    wire N__14199;
    wire N__14198;
    wire N__14191;
    wire N__14182;
    wire N__14179;
    wire N__14178;
    wire N__14177;
    wire N__14174;
    wire N__14167;
    wire N__14162;
    wire N__14157;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14126;
    wire N__14123;
    wire N__14120;
    wire N__14119;
    wire N__14118;
    wire N__14117;
    wire N__14116;
    wire N__14115;
    wire N__14114;
    wire N__14113;
    wire N__14112;
    wire N__14111;
    wire N__14108;
    wire N__14103;
    wire N__14102;
    wire N__14099;
    wire N__14098;
    wire N__14097;
    wire N__14094;
    wire N__14093;
    wire N__14092;
    wire N__14087;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14077;
    wire N__14076;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14045;
    wire N__14040;
    wire N__14039;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14027;
    wire N__14020;
    wire N__14015;
    wire N__14012;
    wire N__14007;
    wire N__14002;
    wire N__14001;
    wire N__14000;
    wire N__13999;
    wire N__13994;
    wire N__13985;
    wire N__13980;
    wire N__13975;
    wire N__13972;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13928;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13826;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13808;
    wire N__13807;
    wire N__13806;
    wire N__13805;
    wire N__13804;
    wire N__13803;
    wire N__13800;
    wire N__13799;
    wire N__13798;
    wire N__13797;
    wire N__13796;
    wire N__13795;
    wire N__13794;
    wire N__13791;
    wire N__13790;
    wire N__13785;
    wire N__13776;
    wire N__13773;
    wire N__13768;
    wire N__13763;
    wire N__13760;
    wire N__13757;
    wire N__13752;
    wire N__13739;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13728;
    wire N__13727;
    wire N__13724;
    wire N__13723;
    wire N__13722;
    wire N__13721;
    wire N__13720;
    wire N__13719;
    wire N__13718;
    wire N__13717;
    wire N__13716;
    wire N__13715;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13696;
    wire N__13693;
    wire N__13684;
    wire N__13681;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13654;
    wire N__13651;
    wire N__13648;
    wire N__13647;
    wire N__13642;
    wire N__13641;
    wire N__13640;
    wire N__13637;
    wire N__13636;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13625;
    wire N__13624;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13616;
    wire N__13615;
    wire N__13612;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13595;
    wire N__13594;
    wire N__13593;
    wire N__13592;
    wire N__13587;
    wire N__13584;
    wire N__13581;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13567;
    wire N__13564;
    wire N__13561;
    wire N__13558;
    wire N__13555;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13536;
    wire N__13533;
    wire N__13530;
    wire N__13527;
    wire N__13524;
    wire N__13517;
    wire N__13514;
    wire N__13511;
    wire N__13504;
    wire N__13501;
    wire N__13498;
    wire N__13497;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13470;
    wire N__13467;
    wire N__13464;
    wire N__13461;
    wire N__13454;
    wire N__13453;
    wire N__13452;
    wire N__13449;
    wire N__13446;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13438;
    wire N__13435;
    wire N__13432;
    wire N__13429;
    wire N__13428;
    wire N__13427;
    wire N__13426;
    wire N__13425;
    wire N__13424;
    wire N__13423;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13413;
    wire N__13410;
    wire N__13407;
    wire N__13402;
    wire N__13397;
    wire N__13392;
    wire N__13389;
    wire N__13370;
    wire N__13367;
    wire N__13366;
    wire N__13363;
    wire N__13360;
    wire N__13355;
    wire N__13354;
    wire N__13349;
    wire N__13346;
    wire N__13343;
    wire N__13340;
    wire N__13337;
    wire N__13336;
    wire N__13335;
    wire N__13334;
    wire N__13333;
    wire N__13332;
    wire N__13331;
    wire N__13330;
    wire N__13329;
    wire N__13326;
    wire N__13321;
    wire N__13314;
    wire N__13311;
    wire N__13306;
    wire N__13301;
    wire N__13298;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13282;
    wire N__13281;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13269;
    wire N__13262;
    wire N__13259;
    wire N__13258;
    wire N__13255;
    wire N__13252;
    wire N__13249;
    wire N__13246;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13222;
    wire N__13221;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13209;
    wire N__13202;
    wire N__13201;
    wire N__13200;
    wire N__13199;
    wire N__13198;
    wire N__13197;
    wire N__13196;
    wire N__13195;
    wire N__13194;
    wire N__13193;
    wire N__13192;
    wire N__13185;
    wire N__13182;
    wire N__13181;
    wire N__13178;
    wire N__13173;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13157;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13145;
    wire N__13138;
    wire N__13127;
    wire N__13124;
    wire N__13123;
    wire N__13122;
    wire N__13121;
    wire N__13120;
    wire N__13117;
    wire N__13116;
    wire N__13115;
    wire N__13114;
    wire N__13113;
    wire N__13110;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13093;
    wire N__13090;
    wire N__13087;
    wire N__13086;
    wire N__13081;
    wire N__13080;
    wire N__13077;
    wire N__13068;
    wire N__13065;
    wire N__13062;
    wire N__13059;
    wire N__13056;
    wire N__13051;
    wire N__13040;
    wire N__13037;
    wire N__13036;
    wire N__13035;
    wire N__13034;
    wire N__13033;
    wire N__13032;
    wire N__13029;
    wire N__13028;
    wire N__13027;
    wire N__13026;
    wire N__13025;
    wire N__13022;
    wire N__13021;
    wire N__13020;
    wire N__13019;
    wire N__13018;
    wire N__13017;
    wire N__13014;
    wire N__13011;
    wire N__13010;
    wire N__13007;
    wire N__12996;
    wire N__12993;
    wire N__12990;
    wire N__12987;
    wire N__12984;
    wire N__12981;
    wire N__12976;
    wire N__12971;
    wire N__12968;
    wire N__12963;
    wire N__12956;
    wire N__12947;
    wire N__12938;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12925;
    wire N__12924;
    wire N__12923;
    wire N__12922;
    wire N__12921;
    wire N__12920;
    wire N__12919;
    wire N__12918;
    wire N__12917;
    wire N__12916;
    wire N__12907;
    wire N__12902;
    wire N__12897;
    wire N__12896;
    wire N__12895;
    wire N__12892;
    wire N__12889;
    wire N__12886;
    wire N__12885;
    wire N__12884;
    wire N__12883;
    wire N__12876;
    wire N__12873;
    wire N__12870;
    wire N__12865;
    wire N__12862;
    wire N__12857;
    wire N__12854;
    wire N__12853;
    wire N__12850;
    wire N__12847;
    wire N__12844;
    wire N__12837;
    wire N__12832;
    wire N__12829;
    wire N__12826;
    wire N__12821;
    wire N__12812;
    wire N__12809;
    wire N__12808;
    wire N__12807;
    wire N__12802;
    wire N__12799;
    wire N__12796;
    wire N__12793;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12766;
    wire N__12765;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12746;
    wire N__12743;
    wire N__12742;
    wire N__12739;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12719;
    wire N__12718;
    wire N__12717;
    wire N__12714;
    wire N__12713;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12690;
    wire N__12685;
    wire N__12682;
    wire N__12679;
    wire N__12676;
    wire N__12673;
    wire N__12668;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12644;
    wire N__12641;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12617;
    wire N__12614;
    wire N__12611;
    wire N__12608;
    wire N__12605;
    wire N__12602;
    wire N__12599;
    wire N__12596;
    wire N__12593;
    wire N__12590;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12520;
    wire N__12517;
    wire N__12514;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12502;
    wire N__12499;
    wire N__12496;
    wire N__12491;
    wire N__12490;
    wire N__12489;
    wire N__12488;
    wire N__12487;
    wire N__12484;
    wire N__12481;
    wire N__12474;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12458;
    wire N__12455;
    wire N__12452;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12437;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12425;
    wire N__12422;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12401;
    wire N__12398;
    wire N__12395;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12368;
    wire N__12365;
    wire N__12362;
    wire N__12359;
    wire N__12356;
    wire N__12353;
    wire N__12350;
    wire N__12347;
    wire N__12346;
    wire N__12343;
    wire N__12340;
    wire N__12335;
    wire N__12332;
    wire N__12331;
    wire N__12330;
    wire N__12325;
    wire N__12322;
    wire N__12317;
    wire N__12314;
    wire N__12311;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12287;
    wire N__12284;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12260;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12199;
    wire N__12194;
    wire N__12191;
    wire N__12190;
    wire N__12189;
    wire N__12188;
    wire N__12187;
    wire N__12186;
    wire N__12183;
    wire N__12176;
    wire N__12171;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12149;
    wire N__12148;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12077;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12038;
    wire N__12035;
    wire N__12032;
    wire N__12029;
    wire N__12026;
    wire N__12023;
    wire N__12020;
    wire N__12017;
    wire N__12014;
    wire N__12011;
    wire N__12008;
    wire N__12005;
    wire N__12004;
    wire N__12001;
    wire N__11998;
    wire N__11993;
    wire N__11990;
    wire N__11989;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11972;
    wire N__11969;
    wire N__11964;
    wire N__11961;
    wire N__11958;
    wire N__11953;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11939;
    wire N__11936;
    wire N__11933;
    wire N__11932;
    wire N__11931;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11911;
    wire N__11908;
    wire N__11905;
    wire N__11900;
    wire N__11897;
    wire N__11896;
    wire N__11891;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11879;
    wire N__11878;
    wire N__11875;
    wire N__11872;
    wire N__11871;
    wire N__11870;
    wire N__11863;
    wire N__11860;
    wire N__11857;
    wire N__11854;
    wire N__11849;
    wire N__11846;
    wire N__11843;
    wire N__11840;
    wire N__11837;
    wire N__11836;
    wire N__11835;
    wire N__11832;
    wire N__11827;
    wire N__11822;
    wire N__11821;
    wire N__11818;
    wire N__11815;
    wire N__11810;
    wire N__11807;
    wire N__11804;
    wire N__11803;
    wire N__11802;
    wire N__11799;
    wire N__11794;
    wire N__11789;
    wire N__11788;
    wire N__11785;
    wire N__11782;
    wire N__11777;
    wire N__11774;
    wire N__11773;
    wire N__11772;
    wire N__11769;
    wire N__11764;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11747;
    wire N__11744;
    wire N__11741;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11714;
    wire N__11711;
    wire N__11708;
    wire N__11705;
    wire N__11702;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11690;
    wire N__11687;
    wire N__11684;
    wire N__11681;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11666;
    wire N__11663;
    wire N__11660;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11645;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11602;
    wire N__11601;
    wire N__11598;
    wire N__11595;
    wire N__11592;
    wire N__11589;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11573;
    wire N__11570;
    wire N__11565;
    wire N__11562;
    wire N__11555;
    wire N__11554;
    wire N__11551;
    wire N__11550;
    wire N__11549;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11541;
    wire N__11538;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11514;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11487;
    wire N__11480;
    wire N__11477;
    wire N__11476;
    wire N__11475;
    wire N__11472;
    wire N__11471;
    wire N__11470;
    wire N__11469;
    wire N__11468;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11447;
    wire N__11446;
    wire N__11445;
    wire N__11442;
    wire N__11441;
    wire N__11436;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11406;
    wire N__11397;
    wire N__11394;
    wire N__11391;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11341;
    wire N__11340;
    wire N__11339;
    wire N__11338;
    wire N__11337;
    wire N__11336;
    wire N__11335;
    wire N__11334;
    wire N__11333;
    wire N__11330;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11302;
    wire N__11301;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11289;
    wire N__11284;
    wire N__11281;
    wire N__11276;
    wire N__11273;
    wire N__11272;
    wire N__11271;
    wire N__11268;
    wire N__11263;
    wire N__11260;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11246;
    wire N__11243;
    wire N__11242;
    wire N__11241;
    wire N__11236;
    wire N__11233;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11218;
    wire N__11217;
    wire N__11214;
    wire N__11211;
    wire N__11208;
    wire N__11205;
    wire N__11202;
    wire N__11199;
    wire N__11196;
    wire N__11191;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11179;
    wire N__11178;
    wire N__11175;
    wire N__11172;
    wire N__11169;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11150;
    wire N__11149;
    wire N__11148;
    wire N__11145;
    wire N__11144;
    wire N__11143;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11132;
    wire N__11131;
    wire N__11128;
    wire N__11125;
    wire N__11124;
    wire N__11123;
    wire N__11122;
    wire N__11119;
    wire N__11118;
    wire N__11117;
    wire N__11116;
    wire N__11111;
    wire N__11110;
    wire N__11107;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11093;
    wire N__11092;
    wire N__11089;
    wire N__11088;
    wire N__11087;
    wire N__11086;
    wire N__11085;
    wire N__11084;
    wire N__11081;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11050;
    wire N__11047;
    wire N__11042;
    wire N__11037;
    wire N__11034;
    wire N__11027;
    wire N__11022;
    wire N__11013;
    wire N__11010;
    wire N__10997;
    wire N__10996;
    wire N__10993;
    wire N__10992;
    wire N__10991;
    wire N__10990;
    wire N__10987;
    wire N__10984;
    wire N__10983;
    wire N__10982;
    wire N__10981;
    wire N__10980;
    wire N__10979;
    wire N__10976;
    wire N__10975;
    wire N__10974;
    wire N__10973;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10965;
    wire N__10964;
    wire N__10963;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10932;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10924;
    wire N__10923;
    wire N__10916;
    wire N__10911;
    wire N__10910;
    wire N__10909;
    wire N__10908;
    wire N__10907;
    wire N__10906;
    wire N__10899;
    wire N__10894;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10867;
    wire N__10864;
    wire N__10861;
    wire N__10858;
    wire N__10855;
    wire N__10852;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10834;
    wire N__10831;
    wire N__10826;
    wire N__10821;
    wire N__10814;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10672;
    wire N__10671;
    wire N__10670;
    wire N__10667;
    wire N__10662;
    wire N__10659;
    wire N__10652;
    wire N__10651;
    wire N__10650;
    wire N__10649;
    wire N__10648;
    wire N__10647;
    wire N__10644;
    wire N__10641;
    wire N__10634;
    wire N__10631;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10612;
    wire N__10611;
    wire N__10610;
    wire N__10609;
    wire N__10606;
    wire N__10603;
    wire N__10600;
    wire N__10595;
    wire N__10586;
    wire N__10585;
    wire N__10584;
    wire N__10581;
    wire N__10580;
    wire N__10577;
    wire N__10572;
    wire N__10569;
    wire N__10562;
    wire N__10559;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10447;
    wire N__10446;
    wire N__10445;
    wire N__10444;
    wire N__10441;
    wire N__10440;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10428;
    wire N__10421;
    wire N__10412;
    wire N__10411;
    wire N__10410;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10400;
    wire N__10399;
    wire N__10398;
    wire N__10397;
    wire N__10396;
    wire N__10393;
    wire N__10386;
    wire N__10377;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10255;
    wire N__10252;
    wire N__10251;
    wire N__10250;
    wire N__10247;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10237;
    wire N__10232;
    wire N__10223;
    wire N__10222;
    wire N__10221;
    wire N__10220;
    wire N__10219;
    wire N__10216;
    wire N__10215;
    wire N__10212;
    wire N__10209;
    wire N__10208;
    wire N__10203;
    wire N__10202;
    wire N__10201;
    wire N__10200;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10171;
    wire N__10170;
    wire N__10169;
    wire N__10168;
    wire N__10165;
    wire N__10164;
    wire N__10163;
    wire N__10162;
    wire N__10161;
    wire N__10160;
    wire N__10159;
    wire N__10154;
    wire N__10141;
    wire N__10136;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10111;
    wire N__10094;
    wire N__10093;
    wire N__10090;
    wire N__10087;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10077;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10061;
    wire N__10060;
    wire N__10057;
    wire N__10056;
    wire N__10055;
    wire N__10054;
    wire N__10053;
    wire N__10052;
    wire N__10051;
    wire N__10050;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10034;
    wire N__10033;
    wire N__10032;
    wire N__10029;
    wire N__10028;
    wire N__10027;
    wire N__10026;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10009;
    wire N__10004;
    wire N__10001;
    wire N__9996;
    wire N__9991;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9863;
    wire N__9860;
    wire N__9859;
    wire N__9858;
    wire N__9855;
    wire N__9854;
    wire N__9851;
    wire N__9850;
    wire N__9847;
    wire N__9844;
    wire N__9841;
    wire N__9840;
    wire N__9839;
    wire N__9834;
    wire N__9831;
    wire N__9826;
    wire N__9821;
    wire N__9816;
    wire N__9813;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9796;
    wire N__9795;
    wire N__9794;
    wire N__9793;
    wire N__9792;
    wire N__9791;
    wire N__9790;
    wire N__9787;
    wire N__9786;
    wire N__9785;
    wire N__9782;
    wire N__9781;
    wire N__9780;
    wire N__9779;
    wire N__9774;
    wire N__9769;
    wire N__9764;
    wire N__9757;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9731;
    wire N__9730;
    wire N__9725;
    wire N__9722;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9710;
    wire N__9707;
    wire N__9706;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9694;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9634;
    wire N__9633;
    wire N__9628;
    wire N__9625;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9613;
    wire N__9608;
    wire N__9607;
    wire N__9604;
    wire N__9601;
    wire N__9598;
    wire N__9593;
    wire N__9590;
    wire N__9589;
    wire N__9588;
    wire N__9583;
    wire N__9582;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9570;
    wire N__9563;
    wire N__9560;
    wire N__9559;
    wire N__9558;
    wire N__9555;
    wire N__9550;
    wire N__9549;
    wire N__9544;
    wire N__9541;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9508;
    wire N__9507;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9495;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9466;
    wire N__9463;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9424;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9412;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9397;
    wire N__9394;
    wire N__9393;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9378;
    wire N__9371;
    wire N__9370;
    wire N__9369;
    wire N__9368;
    wire N__9367;
    wire N__9364;
    wire N__9359;
    wire N__9358;
    wire N__9357;
    wire N__9352;
    wire N__9347;
    wire N__9342;
    wire N__9335;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9277;
    wire N__9274;
    wire N__9273;
    wire N__9272;
    wire N__9271;
    wire N__9268;
    wire N__9265;
    wire N__9262;
    wire N__9257;
    wire N__9254;
    wire N__9245;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9233;
    wire N__9232;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9224;
    wire N__9223;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9188;
    wire N__9187;
    wire N__9186;
    wire N__9185;
    wire N__9182;
    wire N__9181;
    wire N__9180;
    wire N__9179;
    wire N__9176;
    wire N__9171;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9146;
    wire N__9145;
    wire N__9144;
    wire N__9143;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9135;
    wire N__9134;
    wire N__9133;
    wire N__9130;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9114;
    wire N__9111;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9069;
    wire N__9068;
    wire N__9063;
    wire N__9062;
    wire N__9059;
    wire N__9058;
    wire N__9055;
    wire N__9054;
    wire N__9051;
    wire N__9048;
    wire N__9045;
    wire N__9042;
    wire N__9039;
    wire N__9036;
    wire N__9033;
    wire N__9030;
    wire N__9023;
    wire N__9020;
    wire N__9011;
    wire N__9010;
    wire N__9007;
    wire N__9006;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8971;
    wire N__8970;
    wire N__8967;
    wire N__8964;
    wire N__8961;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8914;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8888;
    wire N__8887;
    wire N__8886;
    wire N__8885;
    wire N__8884;
    wire N__8883;
    wire N__8882;
    wire N__8877;
    wire N__8872;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8852;
    wire N__8851;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8789;
    wire N__8786;
    wire N__8785;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8777;
    wire N__8776;
    wire N__8775;
    wire N__8774;
    wire N__8771;
    wire N__8766;
    wire N__8763;
    wire N__8758;
    wire N__8755;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8734;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8710;
    wire N__8709;
    wire N__8708;
    wire N__8705;
    wire N__8700;
    wire N__8697;
    wire N__8690;
    wire N__8687;
    wire N__8686;
    wire N__8681;
    wire N__8680;
    wire N__8679;
    wire N__8678;
    wire N__8677;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8665;
    wire N__8664;
    wire N__8663;
    wire N__8662;
    wire N__8659;
    wire N__8656;
    wire N__8649;
    wire N__8642;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8620;
    wire N__8619;
    wire N__8618;
    wire N__8615;
    wire N__8610;
    wire N__8607;
    wire N__8600;
    wire N__8599;
    wire N__8598;
    wire N__8595;
    wire N__8594;
    wire N__8593;
    wire N__8588;
    wire N__8581;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8503;
    wire N__8500;
    wire N__8497;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8443;
    wire N__8440;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8321;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8236;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8216;
    wire N__8213;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8165;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8077;
    wire N__8076;
    wire N__8073;
    wire N__8068;
    wire N__8065;
    wire N__8060;
    wire N__8059;
    wire N__8058;
    wire N__8055;
    wire N__8054;
    wire N__8049;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8037;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7990;
    wire N__7987;
    wire N__7984;
    wire N__7981;
    wire N__7978;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7796;
    wire N__7793;
    wire N__7790;
    wire N__7787;
    wire N__7784;
    wire N__7781;
    wire N__7780;
    wire N__7777;
    wire N__7776;
    wire N__7775;
    wire N__7774;
    wire N__7771;
    wire N__7770;
    wire N__7767;
    wire N__7764;
    wire N__7759;
    wire N__7754;
    wire N__7745;
    wire N__7742;
    wire N__7739;
    wire N__7738;
    wire N__7735;
    wire N__7732;
    wire N__7727;
    wire N__7724;
    wire N__7723;
    wire N__7722;
    wire N__7721;
    wire N__7720;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7708;
    wire N__7703;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7526;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7514;
    wire N__7511;
    wire N__7510;
    wire N__7507;
    wire N__7504;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7486;
    wire N__7483;
    wire N__7480;
    wire N__7477;
    wire N__7474;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7453;
    wire N__7450;
    wire N__7447;
    wire N__7444;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7430;
    wire N__7427;
    wire VCCG0;
    wire N_377_i;
    wire port_nmib_0_i;
    wire port_clk_c;
    wire \this_delay_clk.M_pipe_qZ0Z_0 ;
    wire rgb_c_0;
    wire i7_mux_0;
    wire rgb_c_1;
    wire N_28_0;
    wire rgb_c_5;
    wire \this_vga_signals.new_pixel_1_1_cascade_ ;
    wire debug_c_0_cascade_;
    wire rgb_c_3;
    wire N_37;
    wire rgb_c_4;
    wire \this_vga_signals.new_pixel_1_3_1_cascade_ ;
    wire \this_vga_signals.new_pixel_sx_0 ;
    wire this_vga_signals_vvisibility_i;
    wire N_60;
    wire i7_mux;
    wire N_50_cascade_;
    wire debug_c_0;
    wire rgb_c_2;
    wire M_hcounter_q_esr_RNIH8GJ4_9;
    wire bfn_6_21_0_;
    wire \this_vga_signals.new_pixel_1Z0Z_1 ;
    wire \this_vga_signals.new_pixel_1_cry_0 ;
    wire \this_vga_signals.new_pixel_1_2 ;
    wire \this_vga_signals.new_pixel_1_cry_1 ;
    wire \this_vga_signals.new_pixel_1_3 ;
    wire \this_vga_signals.new_pixel_1_cry_2 ;
    wire \this_vga_signals.new_pixel_1_4 ;
    wire \this_vga_signals.new_pixel_1_cry_3 ;
    wire \this_vga_signals.new_pixel_1_5 ;
    wire \this_vga_signals.new_pixel_1_cry_4 ;
    wire \this_vga_signals.new_pixel_1_6 ;
    wire \this_vga_signals.new_pixel_1_cry_5 ;
    wire \this_vga_signals.M_hcounter_q_i_7 ;
    wire \this_vga_signals.new_pixel_1_7 ;
    wire \this_vga_signals.new_pixel_1_cry_6 ;
    wire \this_vga_signals.new_pixel_1_cry_7 ;
    wire \this_vga_signals.new_pixel_1_8 ;
    wire bfn_6_22_0_;
    wire \this_vga_signals.new_pixel_1_9 ;
    wire \this_vga_signals.new_pixel_1_cry_8 ;
    wire \this_vga_signals.new_pixel_1_10 ;
    wire \this_vga_signals.new_pixel_1_cry_9 ;
    wire \this_vga_signals.new_pixel_1_cry_10 ;
    wire \this_vga_signals.new_pixel_1_11 ;
    wire \this_vga_signals.un4_hsynclt8_0 ;
    wire this_vga_signals_hsync_1_i;
    wire debug_c_i_1;
    wire \this_vga_signals.M_hcounter_q_esr_RNIG53K_1Z0Z_9 ;
    wire \this_vga_signals.un3_hsynclt8_0 ;
    wire \this_vga_signals.new_pixel_1_i_0 ;
    wire \this_vga_signals.M_hcounter_q_RNIUA42NDZ0Z_1 ;
    wire \this_vga_signals.new_pixel_1_cry_0_c_RNOZ0 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNIG53KZ0Z_9 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_4_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_5_cascade_ ;
    wire \this_vga_signals.g0_13_N_3L3_x0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_2_0_0 ;
    wire \this_vga_signals.g0_13_N_3L3_x1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_cascade_ ;
    wire M_this_vga_signals_address_3;
    wire \this_vga_signals.M_hcounter_d6lt9_cascade_ ;
    wire this_pixel_clock_M_counter_q_i_1;
    wire this_pixel_clock_M_counter_q_0;
    wire \this_vga_signals.M_hcounter_d6_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_q_esr_RNIUKG82Z0Z_9 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_1_sx_cascade_ ;
    wire \this_vga_signals.if_m2_0_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axb2_i_1_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_1 ;
    wire \this_vga_signals.N_4_i_1_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_ac0_1_cascade_ ;
    wire \this_vga_signals.N_4_i ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.M_hcounter_q_esr_RNIGF3C6Z0Z_9_cascade_ ;
    wire \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TAZ0Z7 ;
    wire bfn_9_23_0_;
    wire \this_vga_signals.mult1_un75_sum_i_0_3 ;
    wire \this_vga_signals.un1_haddress_0_axb_2_l_ofxZ0 ;
    wire \this_vga_signals.un1_haddress_0_cry_1_c_RNIDP44VZ0Z02 ;
    wire \this_vga_signals.un1_haddress_0_cry_1 ;
    wire \this_vga_signals.un1_haddress_0_axb_3_l_fxZ0 ;
    wire \this_vga_signals.mult1_un68_sum_i_3 ;
    wire \this_vga_signals.un1_haddress_0_cry_2_c_RNIVPNA9DZ0 ;
    wire \this_vga_signals.un1_haddress_0_cry_2 ;
    wire \this_vga_signals.un1_haddress_0_axb_4_l_fxZ0 ;
    wire \this_vga_signals.un1_haddress_0_cry_3_c_RNIBO4TZ0Z72 ;
    wire \this_vga_signals.un1_haddress_0_cry_3 ;
    wire \this_vga_signals.un1_haddress_0_cry_4_c_RNI5SHJLZ0 ;
    wire \this_vga_signals.un1_haddress_0_cry_4 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNIGF3C6Z0Z_9 ;
    wire \this_vga_signals.un1_haddress_0_cry_5_THRU_CO ;
    wire \this_vga_signals.un1_haddress_0_cry_5 ;
    wire \this_vga_signals.un1_haddress_0_axb_7 ;
    wire \this_vga_signals.un1_haddress_0_cry_6_c_RNI5KQUZ0 ;
    wire \this_vga_signals.un1_haddress_0_cry_6 ;
    wire \this_vga_signals.un1_haddress_0_cry_7_i ;
    wire \this_vga_signals.un1_haddress_0_cry_7 ;
    wire \this_vga_signals.un1_haddress_0_cry_7_c_RNIRVBSZ0Z7 ;
    wire \this_vga_signals.m8_0_1_tz_cascade_ ;
    wire \this_vga_signals.g1_cascade_ ;
    wire \this_vga_signals.g1_1_0_cascade_ ;
    wire \this_vga_signals.N_75_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_m_1_1 ;
    wire \this_vga_signals.mult1_un54_sum_m_1_1_cascade_ ;
    wire \this_vga_signals.N_75 ;
    wire \this_vga_signals.mult1_un54_sum_m_x0_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_m_x1_1 ;
    wire \this_vga_signals.M_hcounter_q_7_rep1_esr_RNIJOMZ0Z71_cascade_ ;
    wire \this_vga_signals.m8_0_2_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_i_0_3_cascade_ ;
    wire \this_vga_signals.g1_6_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3 ;
    wire \this_vga_signals.g0_13_N_3L3_ns ;
    wire \this_vga_signals.g0_13_N_2L1_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axb2_0_0 ;
    wire \this_vga_signals.mult1_un75_sum_axb2_0_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5 ;
    wire \this_vga_signals.if_m2_0 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5_cascade_ ;
    wire \this_vga_signals.g0_10_3_0_a2_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_1 ;
    wire \this_vga_signals.g1_0 ;
    wire \this_vga_signals.g0_10_3_0_a2_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axb2_x0 ;
    wire \this_vga_signals.mult1_un75_sum_axb2_x1 ;
    wire \this_vga_signals.mult1_un75_sum_axb2_i_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_3_0_1_x1 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_3_0_1_x0_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_ac0_1 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_3_0_1_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axb2_i ;
    wire \this_vga_signals.mult1_un75_sum_axbxc2 ;
    wire \this_vga_signals.N_510_i ;
    wire \this_vga_signals.mult1_un61_sum_c3 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axb1 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1_i_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_ac0_3_0_0_cascade_ ;
    wire \this_vga_signals.new_pixel_1_axb_1_N_4L5_xZ0Z1_cascade_ ;
    wire \this_vga_signals.M_hcounter_q_RNIPIQRNRZ0Z_2 ;
    wire \this_vga_signals.M_hcounter_q_RNI5HOBQCZ0Z_1 ;
    wire \this_vga_signals.M_hcounter_q_RNI8TTVN32Z0Z_2_cascade_ ;
    wire \this_vga_signals.new_pixel_1_axb_1 ;
    wire \this_vga_signals.N_510_cascade_ ;
    wire \this_vga_signals.un1_haddress_0_axb_6 ;
    wire \this_vga_signals.un1_haddress_0 ;
    wire \this_vga_signals.mult1_un89_sum_axbxc3_0_cascade_ ;
    wire \this_vga_signals.un1_haddress_0_cry_1_c_RNOZ0 ;
    wire \this_vga_signals.m8_0_1_tz ;
    wire \this_vga_signals.ANC2_4_1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2_cascade_ ;
    wire \this_vga_signals.M_hcounter_q_7_repZ0Z1 ;
    wire \this_vga_signals.M_hcounter_q_5_repZ0Z1 ;
    wire \this_vga_signals.M_hcounter_q_fastZ0Z_9 ;
    wire \this_vga_signals.M_hcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.M_hcounter_q_6_repZ0Z1 ;
    wire \this_vga_signals.M_hcounter_q_9_repZ0Z1 ;
    wire \this_vga_signals.M_hcounter_q_fast_esr_RNIHH441Z0Z_5_cascade_ ;
    wire \this_vga_signals.M_hcounter_q_fast_esr_RNIN6RRZ0Z_7 ;
    wire \this_vga_signals.M_hcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.M_hcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.N_550_1 ;
    wire \this_vga_signals.m8_0_2 ;
    wire \this_vga_signals.g1_0_1 ;
    wire \this_vga_signals.g4_1_1_cascade_ ;
    wire \this_vga_signals.M_hcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.M_hcounter_q_fast_esr_RNI52HLZ0Z_9 ;
    wire \this_vga_signals.m8_0_1_0 ;
    wire \this_vga_signals.M_hcounter_q_8_repZ0Z1 ;
    wire \this_vga_signals.m8_0_3 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_3 ;
    wire \this_vga_signals.g1_1_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_2_0 ;
    wire \this_vga_signals.g1_0_0_cascade_ ;
    wire \this_vga_signals.g1_6_0 ;
    wire \this_vga_signals.g4_1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_1_1 ;
    wire \this_vga_signals.g0_13_N_4L5 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_1_1_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_3 ;
    wire \this_vga_signals.mult1_un68_sum_1_3 ;
    wire \this_vga_signals.mult1_un75_sum_axb2_i_1_0_0 ;
    wire \this_vga_signals.g4 ;
    wire \this_vga_signals.g0_0_2_cascade_ ;
    wire \this_vga_signals.g1_1_1_0_0 ;
    wire \this_vga_signals.N_4_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_0_3_cascade_ ;
    wire \this_vga_signals.g1_0_a2_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3 ;
    wire \this_vga_signals.N_19 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_3_0_1 ;
    wire \this_vga_signals.mult1_un75_sum_axb2_i_0_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_ac0_1_0 ;
    wire \this_vga_signals.g0_i_x2_0_0_a2_3_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_c3_0_0 ;
    wire \this_vga_signals.if_i4_mux_0_cascade_ ;
    wire \this_vga_signals.g1_0_a2 ;
    wire \this_vga_signals.g0_i_x2_0_0_a2_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0 ;
    wire \this_vga_signals.g1_1 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_0 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_0_3 ;
    wire \this_vga_signals.g0_0_a2_4 ;
    wire \this_vga_signals.mult1_un89_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un89_sum_c3 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3 ;
    wire M_this_vga_signals_address_0;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un82_sum_axb2_i ;
    wire \this_vga_signals.mult1_un82_sum_ac0_1 ;
    wire \this_vga_signals.mult1_un82_sum_ac0_3_0_0 ;
    wire M_this_vga_signals_address_1;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1_i ;
    wire \this_vga_signals.mult1_un75_sum_c3 ;
    wire M_this_vga_signals_address_2;
    wire \this_vga_signals.mult1_un61_sum_ac0_1 ;
    wire \this_vga_signals.mult1_un54_sum_i_0_3 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c ;
    wire \this_vga_signals.mult1_un54_sum_m_ns_1 ;
    wire M_this_vga_signals_address_4;
    wire \this_vga_signals.new_pixel_1 ;
    wire bfn_12_20_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.N_583_g ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRDZ0 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_12_21_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire \this_vga_signals.g0_4_0 ;
    wire debug_c_1;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.g0_0_a2_1 ;
    wire \this_delay_clk.M_pipe_qZ0Z_1 ;
    wire \this_delay_clk.M_pipe_qZ0Z_2 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_1_2 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_1_2_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c2 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_0_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_ac0_4 ;
    wire \this_vga_signals.un2_vsynclt8 ;
    wire this_vga_signals_vsync_1_i;
    wire M_this_vga_signals_address_6;
    wire \this_vga_signals.if_N_9 ;
    wire \this_vga_signals.if_N_10_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c2_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c2_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb1_i ;
    wire \this_vga_signals.SUM_2 ;
    wire \this_vga_signals.mult1_un47_sum_c2 ;
    wire \this_vga_signals.mult1_un47_sum_axb2_0_3 ;
    wire \this_vga_signals.mult1_un47_sum_c2_cascade_ ;
    wire \this_vga_signals.vaddress_6 ;
    wire \this_vga_signals.mult1_un47_sum_axb2_3_tz ;
    wire \this_vga_signals.vaddress_7 ;
    wire \this_vga_signals.M_vcounter_d7lt8_0_cascade_ ;
    wire \this_vga_signals.M_vcounter_d7lt9_cascade_ ;
    wire \this_vga_signals.M_vcounter_d7lto8_1 ;
    wire \this_vga_signals.un6_vvisibilitylt9_0_cascade_ ;
    wire \this_vga_signals.vaddress_c5_i ;
    wire \this_vga_signals.vvisibility ;
    wire \this_vga_signals.vsync_1_0_cascade_ ;
    wire \this_vga_signals.vsync_1_4 ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_ns_1 ;
    wire \this_vga_signals.mult1_un75_sum_c2 ;
    wire \this_vga_signals.mult1_un82_sum_c3_cascade_ ;
    wire M_this_vga_signals_address_7;
    wire \this_vga_signals.mult1_un68_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un75_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_i_1_3 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3 ;
    wire M_this_vga_signals_address_10;
    wire \this_vga_signals.mult1_un82_sum_c3_0_bm ;
    wire \this_vga_signals.mult1_un61_sum_axb2 ;
    wire \this_vga_signals.mult1_un61_sum_c2 ;
    wire \this_vga_signals.if_N_10 ;
    wire M_this_vga_signals_address_9;
    wire \this_vga_signals.mult1_un68_sum_axbxc2_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc2 ;
    wire \this_vga_signals.mult1_un75_sum_c3_0 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc2_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0_0 ;
    wire M_this_vga_signals_address_8;
    wire \this_vga_signals.mult1_un40_sum_c3 ;
    wire \this_vga_signals.mult1_un40_sum_c3_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_x0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_ns_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_axb2_0_3_1_1 ;
    wire \this_vga_signals.M_hcounter_d6_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire bfn_15_20_0_;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_2 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7 ;
    wire \this_vga_signals.GZ0Z_296 ;
    wire bfn_15_21_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_0_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_1_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_2_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_3_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_4_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_5_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_6_THRU_CO ;
    wire bfn_15_22_0_;
    wire \this_vga_signals.M_vcounter_qZ0Z_9 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un54_sum_c2 ;
    wire \this_vga_signals.mult1_un47_sum_i_3 ;
    wire \this_vga_signals.vaddress_8 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_8 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_7 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a2_x1 ;
    wire port_dmab_c_i;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire bfn_16_23_0_;
    wire un1_M_this_data_count_q_cry_0;
    wire un1_M_this_data_count_q_cry_1;
    wire un1_M_this_data_count_q_cry_2;
    wire un1_M_this_data_count_q_cry_3;
    wire un1_M_this_data_count_q_cry_4;
    wire un1_M_this_data_count_q_cry_5;
    wire un1_M_this_data_count_q_cry_6;
    wire un1_M_this_data_count_q_cry_7;
    wire bfn_16_24_0_;
    wire un1_M_this_data_count_q_cry_8;
    wire un1_M_this_data_count_q_cry_9;
    wire un1_M_this_data_count_q_cry_10;
    wire un1_M_this_data_count_q_cry_11;
    wire un1_M_this_data_count_q_cry_12;
    wire un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO;
    wire GNDG0;
    wire un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO;
    wire un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO;
    wire bfn_16_25_0_;
    wire \this_vga_signals.mult1_un54_sum_1_c2_1_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_2Z0Z_9 ;
    wire \this_vga_signals.mult1_un54_sum_1_c2_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_signals.mult1_un54_sum1_i_1_3 ;
    wire M_this_vga_signals_address_5;
    wire \this_vga_signals.vaddress_c2 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_1 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_3 ;
    wire \this_vga_signals.N_550_2 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_6 ;
    wire \this_vga_signals.N_550_0 ;
    wire \this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9 ;
    wire \this_start_data_delay.M_this_state_q_srsts_i_1_2_cascade_ ;
    wire \this_start_data_delay.N_389_1 ;
    wire port_dmab_c;
    wire port_dmab_c_cascade_;
    wire \this_start_data_delay.N_385_cascade_ ;
    wire M_this_data_count_qZ0Z_3;
    wire M_this_data_count_qZ0Z_1;
    wire M_this_data_count_qZ0Z_12;
    wire M_this_data_count_qZ0Z_2;
    wire M_this_data_count_qZ0Z_13;
    wire M_this_data_count_qZ0Z_0;
    wire \this_start_data_delay.M_this_state_q_srsts_i_a2_1_9Z0Z_1 ;
    wire \this_start_data_delay.M_this_state_q_srsts_i_a2_1_6Z0Z_1_cascade_ ;
    wire \this_start_data_delay.N_413 ;
    wire M_this_data_count_qZ0Z_6;
    wire M_this_data_count_qZ0Z_5;
    wire M_this_data_count_qZ0Z_7;
    wire M_this_data_count_qZ0Z_4;
    wire \this_start_data_delay.M_this_state_q_srsts_i_a2_1_8Z0Z_1 ;
    wire M_this_data_count_qZ0Z_10;
    wire M_this_data_count_qZ0Z_8;
    wire M_this_data_count_qZ0Z_11;
    wire M_this_data_count_qZ0Z_9;
    wire \this_start_data_delay.M_this_state_q_srsts_i_a2_1_7Z0Z_1 ;
    wire M_this_state_q_RNI20CEZ0Z_0;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire M_this_state_q_nss_0;
    wire \this_delay_clk.M_pipe_qZ0Z_3 ;
    wire \this_start_data_delay.N_353_0 ;
    wire M_this_start_data_delay_out_0_cascade_;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_11 ;
    wire port_rw_in;
    wire \this_start_data_delay.M_this_state_q_srsts_0_a2_1_4 ;
    wire \this_start_data_delay.N_352_0_cascade_ ;
    wire \this_start_data_delay.M_this_state_q_srsts_0_0_4 ;
    wire port_enb_c;
    wire M_this_delay_clk_out_0;
    wire \this_start_data_delay.M_last_qZ0 ;
    wire \this_start_data_delay.N_352_0 ;
    wire \this_start_data_delay.N_407_cascade_ ;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_1 ;
    wire M_this_state_qZ0Z_6;
    wire M_this_state_qZ0Z_1;
    wire M_this_state_qZ0Z_4;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_4 ;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_9 ;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_2 ;
    wire \this_start_data_delay.N_407 ;
    wire \this_start_data_delay.N_398 ;
    wire \this_start_data_delay.M_this_state_dZ0Z29 ;
    wire \this_start_data_delay.N_396 ;
    wire \this_start_data_delay.M_this_state_dZ0Z27 ;
    wire port_address_in_0;
    wire port_address_in_1;
    wire \this_start_data_delay.M_this_state_dZ0Z28 ;
    wire M_this_vga_signals_address_13;
    wire M_this_vga_signals_address_12;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_5 ;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_3 ;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_7 ;
    wire N_346_0;
    wire M_this_internal_address_q_RNI6EA12Z0Z_0;
    wire bfn_20_21_0_;
    wire M_this_internal_address_qZ0Z_1;
    wire un1_M_this_internal_address_q_cry_0_c_RNI4MQIZ0;
    wire un1_M_this_internal_address_q_cry_0;
    wire M_this_internal_address_qZ0Z_2;
    wire un1_M_this_internal_address_q_cry_1_c_RNI6PRIZ0;
    wire un1_M_this_internal_address_q_cry_1;
    wire M_this_internal_address_qZ0Z_3;
    wire un1_M_this_internal_address_q_cry_2_c_RNI8SSIZ0;
    wire un1_M_this_internal_address_q_cry_2;
    wire M_this_internal_address_qZ0Z_4;
    wire un1_M_this_internal_address_q_cry_3_c_RNIAVTIZ0;
    wire un1_M_this_internal_address_q_cry_3;
    wire M_this_internal_address_qZ0Z_5;
    wire un1_M_this_internal_address_q_cry_4_c_RNIC2VIZ0;
    wire un1_M_this_internal_address_q_cry_4;
    wire un1_M_this_internal_address_q_cry_5;
    wire M_this_internal_address_qZ0Z_7;
    wire un1_M_this_internal_address_q_cry_6_c_RNIG81JZ0;
    wire un1_M_this_internal_address_q_cry_6;
    wire un1_M_this_internal_address_q_cry_7;
    wire bfn_20_22_0_;
    wire M_this_internal_address_qZ0Z_9;
    wire un1_M_this_internal_address_q_cry_8_c_RNIKE3JZ0;
    wire un1_M_this_internal_address_q_cry_8;
    wire un1_M_this_internal_address_q_cry_9;
    wire un1_M_this_internal_address_q_cry_10_c_RNI6I0DZ0;
    wire un1_M_this_internal_address_q_cry_10;
    wire un1_M_this_internal_address_q_cry_11;
    wire un1_M_this_internal_address_q_cry_12;
    wire M_this_internal_address_qZ0Z_0;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_0 ;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_10 ;
    wire un1_M_this_internal_address_q_cry_9_c_RNITQCIZ0;
    wire M_this_internal_address_qZ0Z_10;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_12 ;
    wire un1_M_this_internal_address_q_cry_11_c_RNI8L1DZ0;
    wire un1_M_this_internal_address_q_cry_5_c_RNIE50JZ0;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_13 ;
    wire un1_M_this_internal_address_q_cry_12_c_RNIAO2DZ0;
    wire un1_M_this_internal_address_q_cry_7_c_RNIIB2JZ0;
    wire M_this_internal_address_q_3_sm0_0;
    wire \this_vram.mem_out_bus4_1 ;
    wire \this_vram.mem_out_bus0_1 ;
    wire \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0_cascade_ ;
    wire M_this_vga_signals_address_11;
    wire \this_vram.mem_DOUT_7_i_m2_ns_1_1 ;
    wire M_this_vram_read_data_1;
    wire M_this_internal_address_qZ0Z_6;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_6 ;
    wire M_this_state_qZ0Z_5;
    wire M_this_internal_address_qZ0Z_8;
    wire \this_vram.M_this_internal_address_q_3_ns_1Z0Z_8 ;
    wire port_address_in_3;
    wire port_address_in_2;
    wire \this_start_data_delay.M_this_state_d27Z0Z_2 ;
    wire \this_vram.mem_WE_14 ;
    wire \this_vram.mem_out_bus6_1 ;
    wire \this_vram.mem_out_bus2_1 ;
    wire \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0 ;
    wire \this_vram.mem_out_bus7_1 ;
    wire \this_vram.mem_out_bus3_1 ;
    wire \this_vram.mem_mem_3_0_RNI05P11Z0Z_0 ;
    wire M_this_vram_read_data_3;
    wire \this_vram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ;
    wire M_this_vram_read_data_2;
    wire \this_vram.mem_radregZ0Z_11 ;
    wire \this_vram.mem_DOUT_7_i_m2_ns_1_0 ;
    wire M_this_vram_read_data_0;
    wire port_data_c_1;
    wire port_data_c_5;
    wire M_this_vram_write_data_0_i_1;
    wire M_this_state_qZ0Z_7;
    wire M_this_state_qZ0Z_2;
    wire port_data_c_0;
    wire port_data_c_4;
    wire M_this_vram_write_data_0_sqmuxa_cascade_;
    wire M_this_vram_write_data_0_i_0;
    wire M_this_start_data_delay_out_0;
    wire \this_start_data_delay.N_351_0 ;
    wire \this_vram.mem_WE_8 ;
    wire \this_vram.mem_WE_12 ;
    wire \this_vram.mem_WE_10 ;
    wire \this_vram.mem_out_bus4_2 ;
    wire \this_vram.mem_out_bus0_2 ;
    wire \this_vram.mem_mem_0_1_RNISOIZ0Z11 ;
    wire \this_vram.mem_out_bus5_3 ;
    wire \this_vram.mem_out_bus1_3 ;
    wire \this_vram.mem_out_bus3_3 ;
    wire \this_vram.mem_out_bus7_3 ;
    wire \this_vram.mem_DOUT_6_i_m2_ns_1_3_cascade_ ;
    wire \this_vram.mem_N_102 ;
    wire \this_vram.mem_out_bus4_3 ;
    wire \this_vram.mem_out_bus0_3 ;
    wire \this_vram.mem_out_bus6_3 ;
    wire \this_vram.mem_out_bus2_3 ;
    wire \this_vram.mem_DOUT_3_i_m2_ns_1_3_cascade_ ;
    wire \this_vram.mem_radregZ0Z_12 ;
    wire \this_vram.mem_N_105 ;
    wire \this_vram.mem_out_bus0_0 ;
    wire \this_vram.mem_out_bus4_0 ;
    wire \this_vram.mem_mem_0_0_RNIQOIZ0Z11 ;
    wire \this_vram.mem_out_bus6_0 ;
    wire \this_vram.mem_out_bus2_0 ;
    wire \this_vram.mem_mem_2_0_RNIU0NZ0Z11 ;
    wire \this_vram.mem_WE_6 ;
    wire \this_vram.mem_out_bus1_1 ;
    wire \this_vram.mem_out_bus5_1 ;
    wire \this_vram.mem_mem_1_0_RNISSK11Z0Z_0 ;
    wire \this_vram.mem_out_bus5_2 ;
    wire \this_vram.mem_out_bus1_2 ;
    wire \this_vram.mem_mem_1_1_RNIUSKZ0Z11 ;
    wire \this_vram.mem_out_bus7_2 ;
    wire \this_vram.mem_out_bus3_2 ;
    wire \this_vram.mem_mem_3_1_RNI25PZ0Z11 ;
    wire \this_vram.mem_out_bus7_0 ;
    wire \this_vram.mem_out_bus3_0 ;
    wire \this_vram.mem_mem_3_0_RNI05PZ0Z11 ;
    wire \this_vram.mem_out_bus2_2 ;
    wire \this_vram.mem_out_bus6_2 ;
    wire \this_vram.mem_mem_2_1_RNI01NZ0Z11 ;
    wire \this_vram.mem_radregZ0Z_13 ;
    wire \this_vram.mem_out_bus5_0 ;
    wire \this_vram.mem_out_bus1_0 ;
    wire \this_vram.mem_mem_1_0_RNISSKZ0Z11 ;
    wire port_data_c_3;
    wire port_data_c_7;
    wire M_this_vram_write_data_0_i_3;
    wire \this_vram.mem_WE_4 ;
    wire port_data_c_2;
    wire port_data_c_6;
    wire M_this_vram_write_data_0_sqmuxa;
    wire \this_start_data_delay.un1_M_this_state_q_0 ;
    wire M_this_vram_write_data_0_i_2;
    wire \this_vram.mem_WE_0 ;
    wire M_this_internal_address_qZ0Z_12;
    wire M_this_internal_address_qZ0Z_11;
    wire M_this_internal_address_qZ0Z_13;
    wire M_this_vram_write_en_0_0;
    wire \this_vram.mem_WE_2 ;
    wire CONSTANT_ONE_NET;
    wire M_this_state_qZ0Z_3;
    wire M_this_external_address_qZ0Z_0;
    wire bfn_30_23_0_;
    wire M_this_external_address_qZ0Z_1;
    wire un1_M_this_external_address_q_cry_0;
    wire M_this_external_address_qZ0Z_2;
    wire un1_M_this_external_address_q_cry_1;
    wire M_this_external_address_qZ0Z_3;
    wire un1_M_this_external_address_q_cry_2;
    wire M_this_external_address_qZ0Z_4;
    wire un1_M_this_external_address_q_cry_3;
    wire M_this_external_address_qZ0Z_5;
    wire un1_M_this_external_address_q_cry_4;
    wire M_this_external_address_qZ0Z_6;
    wire un1_M_this_external_address_q_cry_5;
    wire M_this_external_address_qZ0Z_7;
    wire un1_M_this_external_address_q_cry_6;
    wire un1_M_this_external_address_q_cry_7;
    wire M_this_external_address_qZ0Z_8;
    wire bfn_30_24_0_;
    wire M_this_external_address_qZ0Z_9;
    wire un1_M_this_external_address_q_cry_8;
    wire M_this_external_address_qZ0Z_10;
    wire un1_M_this_external_address_q_cry_9;
    wire M_this_external_address_qZ0Z_11;
    wire un1_M_this_external_address_q_cry_10;
    wire M_this_external_address_qZ0Z_12;
    wire un1_M_this_external_address_q_cry_11;
    wire M_this_external_address_qZ0Z_13;
    wire un1_M_this_external_address_q_cry_12;
    wire M_this_external_address_qZ0Z_14;
    wire un1_M_this_external_address_q_cry_13;
    wire M_this_state_qZ0Z_0;
    wire un1_M_this_external_address_q_cry_14;
    wire M_this_external_address_qZ0Z_15;
    wire clk_0_c_g;
    wire M_this_state_q_nss_g_0;
    wire port_address_in_5;
    wire port_address_in_6;
    wire port_address_in_7;
    wire port_address_in_4;
    wire \this_start_data_delay.M_this_state_d27Z0Z_6 ;
    wire _gnd_net_;

    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,\this_vram.mem_out_bus0_1 ,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,\this_vram.mem_out_bus0_0 ,dangling_wire_11,dangling_wire_12,dangling_wire_13}),
            .RADDR({N__12467,N__12311,N__12131,N__12647,N__11732,N__13955,N__9974,N__8198,N__10370,N__10562,N__10784}),
            .WADDR({N__17300,N__16601,N__17642,N__16733,N__17879,N__16868,N__17000,N__17132,N__16256,N__16400,N__17450}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,N__18184,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__18887,dangling_wire_41,dangling_wire_42,dangling_wire_43}),
            .RCLKE(),
            .RCLK(N__21570),
            .RE(N__20438),
            .WCLKE(N__18574),
            .WCLK(N__21571),
            .WE(N__20436));
    defparam \this_vram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,\this_vram.mem_out_bus0_3 ,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,\this_vram.mem_out_bus0_2 ,dangling_wire_55,dangling_wire_56,dangling_wire_57}),
            .RADDR({N__12461,N__12305,N__12125,N__12641,N__11726,N__13949,N__9968,N__8192,N__10364,N__10556,N__10778}),
            .WADDR({N__17294,N__16595,N__17636,N__16727,N__17873,N__16862,N__16994,N__17126,N__16250,N__16394,N__17444}),
            .MASK({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .WDATA({dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,N__19442,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,N__20855,dangling_wire_85,dangling_wire_86,dangling_wire_87}),
            .RCLKE(),
            .RCLK(N__21572),
            .RE(N__20437),
            .WCLKE(N__18575),
            .WCLK(N__21573),
            .WE(N__20435));
    defparam \this_vram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,\this_vram.mem_out_bus1_1 ,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,\this_vram.mem_out_bus1_0 ,dangling_wire_99,dangling_wire_100,dangling_wire_101}),
            .RADDR({N__12455,N__12299,N__12119,N__12635,N__11720,N__13943,N__9962,N__8186,N__10358,N__10550,N__10772}),
            .WADDR({N__17288,N__16589,N__17630,N__16721,N__17867,N__16856,N__16988,N__17120,N__16244,N__16388,N__17438}),
            .MASK({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .WDATA({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__18180,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,N__18883,dangling_wire_129,dangling_wire_130,dangling_wire_131}),
            .RCLKE(),
            .RCLK(N__21574),
            .RE(N__20420),
            .WCLKE(N__18650),
            .WCLK(N__21575),
            .WE(N__20427));
    defparam \this_vram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,\this_vram.mem_out_bus1_3 ,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,\this_vram.mem_out_bus1_2 ,dangling_wire_143,dangling_wire_144,dangling_wire_145}),
            .RADDR({N__12449,N__12293,N__12113,N__12629,N__11714,N__13937,N__9956,N__8180,N__10352,N__10544,N__10766}),
            .WADDR({N__17282,N__16583,N__17624,N__16715,N__17861,N__16850,N__16982,N__17114,N__16238,N__16382,N__17432}),
            .MASK({dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161}),
            .WDATA({dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,N__19438,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,N__20851,dangling_wire_173,dangling_wire_174,dangling_wire_175}),
            .RCLKE(),
            .RCLK(N__21576),
            .RE(N__20419),
            .WCLKE(N__18646),
            .WCLK(N__21577),
            .WE(N__20434));
    defparam \this_vram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,\this_vram.mem_out_bus2_1 ,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,\this_vram.mem_out_bus2_0 ,dangling_wire_187,dangling_wire_188,dangling_wire_189}),
            .RADDR({N__12443,N__12287,N__12107,N__12623,N__11708,N__13931,N__9950,N__8174,N__10346,N__10538,N__10760}),
            .WADDR({N__17276,N__16577,N__17618,N__16709,N__17855,N__16844,N__16976,N__17108,N__16232,N__16376,N__17426}),
            .MASK({dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205}),
            .WDATA({dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,N__18164,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,N__18876,dangling_wire_217,dangling_wire_218,dangling_wire_219}),
            .RCLKE(),
            .RCLK(N__21581),
            .RE(N__20394),
            .WCLKE(N__18623),
            .WCLK(N__21580),
            .WE(N__20415));
    defparam \this_vram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,\this_vram.mem_out_bus2_3 ,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,\this_vram.mem_out_bus2_2 ,dangling_wire_231,dangling_wire_232,dangling_wire_233}),
            .RADDR({N__12437,N__12281,N__12101,N__12617,N__11702,N__13925,N__9944,N__8168,N__10340,N__10532,N__10754}),
            .WADDR({N__17270,N__16571,N__17612,N__16703,N__17849,N__16838,N__16970,N__17102,N__16226,N__16370,N__17420}),
            .MASK({dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249}),
            .WDATA({dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,N__19431,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,N__20844,dangling_wire_261,dangling_wire_262,dangling_wire_263}),
            .RCLKE(),
            .RCLK(N__21585),
            .RE(N__20393),
            .WCLKE(N__18622),
            .WCLK(N__21586),
            .WE(N__20414));
    defparam \this_vram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,\this_vram.mem_out_bus3_1 ,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,\this_vram.mem_out_bus3_0 ,dangling_wire_275,dangling_wire_276,dangling_wire_277}),
            .RADDR({N__12431,N__12275,N__12095,N__12611,N__11696,N__13919,N__9938,N__8162,N__10334,N__10526,N__10748}),
            .WADDR({N__17264,N__16565,N__17606,N__16697,N__17843,N__16832,N__16964,N__17096,N__16220,N__16364,N__17414}),
            .MASK({dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293}),
            .WDATA({dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,N__18185,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,N__18866,dangling_wire_305,dangling_wire_306,dangling_wire_307}),
            .RCLKE(),
            .RCLK(N__21593),
            .RE(N__20362),
            .WCLKE(N__18668),
            .WCLK(N__21594),
            .WE(N__20382));
    defparam \this_vram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,\this_vram.mem_out_bus3_3 ,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,\this_vram.mem_out_bus3_2 ,dangling_wire_319,dangling_wire_320,dangling_wire_321}),
            .RADDR({N__12425,N__12269,N__12089,N__12605,N__11690,N__13913,N__9932,N__8156,N__10328,N__10520,N__10742}),
            .WADDR({N__17258,N__16559,N__17600,N__16691,N__17837,N__16826,N__16958,N__17090,N__16214,N__16358,N__17408}),
            .MASK({dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337}),
            .WDATA({dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,N__19421,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,N__20834,dangling_wire_349,dangling_wire_350,dangling_wire_351}),
            .RCLKE(),
            .RCLK(N__21611),
            .RE(N__20361),
            .WCLKE(N__18661),
            .WCLK(N__21612),
            .WE(N__20381));
    defparam \this_vram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,\this_vram.mem_out_bus4_1 ,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,\this_vram.mem_out_bus4_0 ,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .RADDR({N__12419,N__12263,N__12083,N__12599,N__11684,N__13907,N__9926,N__8150,N__10322,N__10514,N__10736}),
            .WADDR({N__17252,N__16553,N__17594,N__16685,N__17831,N__16820,N__16952,N__17084,N__16208,N__16352,N__17402}),
            .MASK({dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381}),
            .WDATA({dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,N__18171,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,N__18853,dangling_wire_393,dangling_wire_394,dangling_wire_395}),
            .RCLKE(),
            .RCLK(N__21621),
            .RE(N__20324),
            .WCLKE(N__19087),
            .WCLK(N__21622),
            .WE(N__20344));
    defparam \this_vram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,\this_vram.mem_out_bus4_3 ,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,\this_vram.mem_out_bus4_2 ,dangling_wire_407,dangling_wire_408,dangling_wire_409}),
            .RADDR({N__12413,N__12257,N__12077,N__12593,N__11678,N__13901,N__9920,N__8144,N__10316,N__10508,N__10730}),
            .WADDR({N__17246,N__16547,N__17588,N__16679,N__17825,N__16814,N__16946,N__17078,N__16202,N__16346,N__17396}),
            .MASK({dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425}),
            .WDATA({dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,N__19388,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,N__20801,dangling_wire_437,dangling_wire_438,dangling_wire_439}),
            .RCLKE(),
            .RCLK(N__21630),
            .RE(N__20323),
            .WCLKE(N__19091),
            .WCLK(N__21631),
            .WE(N__20343));
    defparam \this_vram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,\this_vram.mem_out_bus5_1 ,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,\this_vram.mem_out_bus5_0 ,dangling_wire_451,dangling_wire_452,dangling_wire_453}),
            .RADDR({N__12407,N__12251,N__12071,N__12587,N__11672,N__13895,N__9914,N__8138,N__10310,N__10502,N__10724}),
            .WADDR({N__17240,N__16541,N__17582,N__16673,N__17819,N__16808,N__16940,N__17072,N__16196,N__16340,N__17390}),
            .MASK({dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469}),
            .WDATA({dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,N__18131,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,N__18831,dangling_wire_481,dangling_wire_482,dangling_wire_483}),
            .RCLKE(),
            .RCLK(N__21635),
            .RE(N__20271),
            .WCLKE(N__19369),
            .WCLK(N__21636),
            .WE(N__20294));
    defparam \this_vram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,\this_vram.mem_out_bus5_3 ,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,\this_vram.mem_out_bus5_2 ,dangling_wire_495,dangling_wire_496,dangling_wire_497}),
            .RADDR({N__12401,N__12245,N__12065,N__12581,N__11666,N__13889,N__9908,N__8132,N__10304,N__10496,N__10718}),
            .WADDR({N__17234,N__16535,N__17576,N__16667,N__17813,N__16802,N__16934,N__17066,N__16190,N__16334,N__17384}),
            .MASK({dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513}),
            .WDATA({dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,N__19402,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,N__20815,dangling_wire_525,dangling_wire_526,dangling_wire_527}),
            .RCLKE(),
            .RCLK(N__21640),
            .RE(N__20188),
            .WCLKE(N__19370),
            .WCLK(N__21641),
            .WE(N__20149));
    defparam \this_vram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,\this_vram.mem_out_bus6_1 ,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,\this_vram.mem_out_bus6_0 ,dangling_wire_539,dangling_wire_540,dangling_wire_541}),
            .RADDR({N__12395,N__12239,N__12059,N__12575,N__11660,N__13883,N__9902,N__8126,N__10298,N__10490,N__10712}),
            .WADDR({N__17228,N__16529,N__17570,N__16661,N__17807,N__16796,N__16928,N__17060,N__16184,N__16328,N__17378}),
            .MASK({dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557}),
            .WDATA({dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,N__18175,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,N__18849,dangling_wire_569,dangling_wire_570,dangling_wire_571}),
            .RCLKE(),
            .RCLK(N__21644),
            .RE(N__20180),
            .WCLKE(N__20455),
            .WCLK(N__21645),
            .WE(N__20207));
    defparam \this_vram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,\this_vram.mem_out_bus6_3 ,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,\this_vram.mem_out_bus6_2 ,dangling_wire_583,dangling_wire_584,dangling_wire_585}),
            .RADDR({N__12389,N__12233,N__12053,N__12569,N__11654,N__13877,N__9896,N__8120,N__10292,N__10484,N__10706}),
            .WADDR({N__17222,N__16523,N__17564,N__16655,N__17801,N__16790,N__16922,N__17054,N__16178,N__16322,N__17372}),
            .MASK({dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601}),
            .WDATA({dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,N__19417,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,N__20830,dangling_wire_613,dangling_wire_614,dangling_wire_615}),
            .RCLKE(),
            .RCLK(N__21646),
            .RE(N__20322),
            .WCLKE(N__20459),
            .WCLK(N__21647),
            .WE(N__20234));
    defparam \this_vram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,\this_vram.mem_out_bus7_1 ,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,\this_vram.mem_out_bus7_0 ,dangling_wire_627,dangling_wire_628,dangling_wire_629}),
            .RADDR({N__12383,N__12227,N__12047,N__12563,N__11648,N__13871,N__9890,N__8114,N__10286,N__10478,N__10700}),
            .WADDR({N__17216,N__16517,N__17558,N__16649,N__17795,N__16784,N__16916,N__17048,N__16172,N__16316,N__17366}),
            .MASK({dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645}),
            .WDATA({dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,N__18176,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,N__18865,dangling_wire_657,dangling_wire_658,dangling_wire_659}),
            .RCLKE(),
            .RCLK(N__21649),
            .RE(N__20305),
            .WCLKE(N__20782),
            .WCLK(N__21650),
            .WE(N__20307));
    defparam \this_vram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,\this_vram.mem_out_bus7_3 ,dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,\this_vram.mem_out_bus7_2 ,dangling_wire_671,dangling_wire_672,dangling_wire_673}),
            .RADDR({N__12377,N__12221,N__12041,N__12557,N__11642,N__13865,N__9884,N__8108,N__10280,N__10472,N__10694}),
            .WADDR({N__17210,N__16511,N__17552,N__16643,N__17789,N__16778,N__16910,N__17042,N__16166,N__16310,N__17360}),
            .MASK({dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689}),
            .WDATA({dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,N__19430,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,N__20843,dangling_wire_701,dangling_wire_702,dangling_wire_703}),
            .RCLKE(),
            .RCLK(N__21652),
            .RE(N__20306),
            .WCLKE(N__20783),
            .WCLK(N__21653),
            .WE(N__20308));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__22314),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__22316),
            .DIN(N__22315),
            .DOUT(N__22314),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__22316),
            .PADOUT(N__22315),
            .PADIN(N__22314),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_0_iopad (
            .OE(N__22305),
            .DIN(N__22304),
            .DOUT(N__22303),
            .PACKAGEPIN(debug[0]));
    defparam debug_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_0_preio (
            .PADOEN(N__22305),
            .PADOUT(N__22304),
            .PADIN(N__22303),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7793),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_1_iopad (
            .OE(N__22296),
            .DIN(N__22295),
            .DOUT(N__22294),
            .PACKAGEPIN(debug[1]));
    defparam debug_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_1_preio (
            .PADOEN(N__22296),
            .PADOUT(N__22295),
            .PADIN(N__22294),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11609),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__22287),
            .DIN(N__22286),
            .DOUT(N__22285),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__22287),
            .PADOUT(N__22286),
            .PADIN(N__22285),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7937),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__22278),
            .DIN(N__22277),
            .DOUT(N__22276),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__22278),
            .PADOUT(N__22277),
            .PADIN(N__22276),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7814),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_iobuf_0_iopad (
            .OE(N__22269),
            .DIN(N__22268),
            .DOUT(N__22267),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_0_preio (
            .PADOEN(N__22269),
            .PADOUT(N__22268),
            .PADIN(N__22267),
            .CLOCKENABLE(),
            .DIN0(port_address_in_0),
            .DIN1(),
            .DOUT0(N__19901),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13580));
    IO_PAD port_address_iobuf_1_iopad (
            .OE(N__22260),
            .DIN(N__22259),
            .DOUT(N__22258),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_1_preio (
            .PADOEN(N__22260),
            .PADOUT(N__22259),
            .PADIN(N__22258),
            .CLOCKENABLE(),
            .DIN0(port_address_in_1),
            .DIN1(),
            .DOUT0(N__19877),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13636));
    IO_PAD port_address_iobuf_2_iopad (
            .OE(N__22251),
            .DIN(N__22250),
            .DOUT(N__22249),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_2_preio (
            .PADOEN(N__22251),
            .PADOUT(N__22250),
            .PADIN(N__22249),
            .CLOCKENABLE(),
            .DIN0(port_address_in_2),
            .DIN1(),
            .DOUT0(N__19853),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13616));
    IO_PAD port_address_iobuf_3_iopad (
            .OE(N__22242),
            .DIN(N__22241),
            .DOUT(N__22240),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_3_preio (
            .PADOEN(N__22242),
            .PADOUT(N__22241),
            .PADIN(N__22240),
            .CLOCKENABLE(),
            .DIN0(port_address_in_3),
            .DIN1(),
            .DOUT0(N__19823),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13640));
    IO_PAD port_address_iobuf_4_iopad (
            .OE(N__22233),
            .DIN(N__22232),
            .DOUT(N__22231),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_4_preio (
            .PADOEN(N__22233),
            .PADOUT(N__22232),
            .PADIN(N__22231),
            .CLOCKENABLE(),
            .DIN0(port_address_in_4),
            .DIN1(),
            .DOUT0(N__19799),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13624));
    IO_PAD port_address_iobuf_5_iopad (
            .OE(N__22224),
            .DIN(N__22223),
            .DOUT(N__22222),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_5_preio (
            .PADOEN(N__22224),
            .PADOUT(N__22223),
            .PADIN(N__22222),
            .CLOCKENABLE(),
            .DIN0(port_address_in_5),
            .DIN1(),
            .DOUT0(N__21173),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13593));
    IO_PAD port_address_iobuf_6_iopad (
            .OE(N__22215),
            .DIN(N__22214),
            .DOUT(N__22213),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_6_preio (
            .PADOEN(N__22215),
            .PADOUT(N__22214),
            .PADIN(N__22213),
            .CLOCKENABLE(),
            .DIN0(port_address_in_6),
            .DIN1(),
            .DOUT0(N__21152),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13623));
    IO_PAD port_address_iobuf_7_iopad (
            .OE(N__22206),
            .DIN(N__22205),
            .DOUT(N__22204),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_7_preio (
            .PADOEN(N__22206),
            .PADOUT(N__22205),
            .PADIN(N__22204),
            .CLOCKENABLE(),
            .DIN0(port_address_in_7),
            .DIN1(),
            .DOUT0(N__21131),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13658));
    IO_PAD port_address_obuft_10_iopad (
            .OE(N__22197),
            .DIN(N__22196),
            .DOUT(N__22195),
            .PACKAGEPIN(port_address[10]));
    defparam port_address_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_10_preio (
            .PADOEN(N__22197),
            .PADOUT(N__22196),
            .PADIN(N__22195),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21050),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13615));
    IO_PAD port_address_obuft_11_iopad (
            .OE(N__22188),
            .DIN(N__22187),
            .DOUT(N__22186),
            .PACKAGEPIN(port_address[11]));
    defparam port_address_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_11_preio (
            .PADOEN(N__22188),
            .PADOUT(N__22187),
            .PADIN(N__22186),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21020),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13647));
    IO_PAD port_address_obuft_12_iopad (
            .OE(N__22179),
            .DIN(N__22178),
            .DOUT(N__22177),
            .PACKAGEPIN(port_address[12]));
    defparam port_address_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_12_preio (
            .PADOEN(N__22179),
            .PADOUT(N__22178),
            .PADIN(N__22177),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21002),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13625));
    IO_PAD port_address_obuft_13_iopad (
            .OE(N__22170),
            .DIN(N__22169),
            .DOUT(N__22168),
            .PACKAGEPIN(port_address[13]));
    defparam port_address_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_13_preio (
            .PADOEN(N__22170),
            .PADOUT(N__22169),
            .PADIN(N__22168),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21908),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13594));
    IO_PAD port_address_obuft_14_iopad (
            .OE(N__22161),
            .DIN(N__22160),
            .DOUT(N__22159),
            .PACKAGEPIN(port_address[14]));
    defparam port_address_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_14_preio (
            .PADOEN(N__22161),
            .PADOUT(N__22160),
            .PADIN(N__22159),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21884),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13641));
    IO_PAD port_address_obuft_15_iopad (
            .OE(N__22152),
            .DIN(N__22151),
            .DOUT(N__22150),
            .PACKAGEPIN(port_address[15]));
    defparam port_address_obuft_15_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_15_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_15_preio (
            .PADOEN(N__22152),
            .PADOUT(N__22151),
            .PADIN(N__22150),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21677),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13654));
    IO_PAD port_address_obuft_8_iopad (
            .OE(N__22143),
            .DIN(N__22142),
            .DOUT(N__22141),
            .PACKAGEPIN(port_address[8]));
    defparam port_address_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_8_preio (
            .PADOEN(N__22143),
            .PADOUT(N__22142),
            .PADIN(N__22141),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21104),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13497));
    IO_PAD port_address_obuft_9_iopad (
            .OE(N__22134),
            .DIN(N__22133),
            .DOUT(N__22132),
            .PACKAGEPIN(port_address[9]));
    defparam port_address_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_9_preio (
            .PADOEN(N__22134),
            .PADOUT(N__22133),
            .PADIN(N__22132),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21071),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13635));
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__22125),
            .DIN(N__22124),
            .DOUT(N__22123),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__22125),
            .PADOUT(N__22124),
            .PADIN(N__22123),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__22116),
            .DIN(N__22115),
            .DOUT(N__22114),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__22116),
            .PADOUT(N__22115),
            .PADIN(N__22114),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__22107),
            .DIN(N__22106),
            .DOUT(N__22105),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__22107),
            .PADOUT(N__22106),
            .PADIN(N__22105),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__22098),
            .DIN(N__22097),
            .DOUT(N__22096),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__22098),
            .PADOUT(N__22097),
            .PADIN(N__22096),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__22089),
            .DIN(N__22088),
            .DOUT(N__22087),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__22089),
            .PADOUT(N__22088),
            .PADIN(N__22087),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__22080),
            .DIN(N__22079),
            .DOUT(N__22078),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__22080),
            .PADOUT(N__22079),
            .PADIN(N__22078),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__22071),
            .DIN(N__22070),
            .DOUT(N__22069),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__22071),
            .PADOUT(N__22070),
            .PADIN(N__22069),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__22062),
            .DIN(N__22061),
            .DOUT(N__22060),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__22062),
            .PADOUT(N__22061),
            .PADIN(N__22060),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_7_iopad (
            .OE(N__22053),
            .DIN(N__22052),
            .DOUT(N__22051),
            .PACKAGEPIN(port_data[7]));
    defparam port_data_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_7_preio (
            .PADOEN(N__22053),
            .PADOUT(N__22052),
            .PADIN(N__22051),
            .CLOCKENABLE(),
            .DIN0(port_data_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__22044),
            .DIN(N__22043),
            .DOUT(N__22042),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__22044),
            .PADOUT(N__22043),
            .PADIN(N__22042),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7430),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__22035),
            .DIN(N__22034),
            .DOUT(N__22033),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__22035),
            .PADOUT(N__22034),
            .PADIN(N__22033),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__14888),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__22026),
            .DIN(N__22025),
            .DOUT(N__22024),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__22026),
            .PADOUT(N__22025),
            .PADIN(N__22024),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__22017),
            .DIN(N__22016),
            .DOUT(N__22015),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__22017),
            .PADOUT(N__22016),
            .PADIN(N__22015),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7553),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_iobuf_iopad (
            .OE(N__22008),
            .DIN(N__22007),
            .DOUT(N__22006),
            .PACKAGEPIN(port_rw));
    defparam port_rw_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO port_rw_iobuf_preio (
            .PADOEN(N__22008),
            .PADOUT(N__22007),
            .PADIN(N__22006),
            .CLOCKENABLE(),
            .DIN0(port_rw_in),
            .DIN1(),
            .DOUT0(N__20392),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__13592));
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__21999),
            .DIN(N__21998),
            .DOUT(N__21997),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__21999),
            .PADOUT(N__21998),
            .PADIN(N__21997),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7526),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__21990),
            .DIN(N__21989),
            .DOUT(N__21988),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__21990),
            .PADOUT(N__21989),
            .PADIN(N__21988),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7493),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__21981),
            .DIN(N__21980),
            .DOUT(N__21979),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__21981),
            .PADOUT(N__21980),
            .PADIN(N__21979),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7745),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__21972),
            .DIN(N__21971),
            .DOUT(N__21970),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__21972),
            .PADOUT(N__21971),
            .PADIN(N__21970),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7646),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__21963),
            .DIN(N__21962),
            .DOUT(N__21961),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__21963),
            .PADOUT(N__21962),
            .PADIN(N__21961),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7616),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__21954),
            .DIN(N__21953),
            .DOUT(N__21952),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__21954),
            .PADOUT(N__21953),
            .PADIN(N__21952),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7460),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__21945),
            .DIN(N__21944),
            .DOUT(N__21943),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__21945),
            .PADOUT(N__21944),
            .PADIN(N__21943),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__21936),
            .DIN(N__21935),
            .DOUT(N__21934),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__21936),
            .PADOUT(N__21935),
            .PADIN(N__21934),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7577),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__21927),
            .DIN(N__21926),
            .DOUT(N__21925),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__21927),
            .PADOUT(N__21926),
            .PADIN(N__21925),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11750),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IoInMux I__5365 (
            .O(N__21908),
            .I(N__21905));
    LocalMux I__5364 (
            .O(N__21905),
            .I(N__21902));
    IoSpan4Mux I__5363 (
            .O(N__21902),
            .I(N__21899));
    Sp12to4 I__5362 (
            .O(N__21899),
            .I(N__21895));
    InMux I__5361 (
            .O(N__21898),
            .I(N__21892));
    Odrv12 I__5360 (
            .O(N__21895),
            .I(M_this_external_address_qZ0Z_13));
    LocalMux I__5359 (
            .O(N__21892),
            .I(M_this_external_address_qZ0Z_13));
    InMux I__5358 (
            .O(N__21887),
            .I(un1_M_this_external_address_q_cry_12));
    IoInMux I__5357 (
            .O(N__21884),
            .I(N__21881));
    LocalMux I__5356 (
            .O(N__21881),
            .I(N__21878));
    Span4Mux_s2_h I__5355 (
            .O(N__21878),
            .I(N__21875));
    Sp12to4 I__5354 (
            .O(N__21875),
            .I(N__21871));
    InMux I__5353 (
            .O(N__21874),
            .I(N__21868));
    Odrv12 I__5352 (
            .O(N__21871),
            .I(M_this_external_address_qZ0Z_14));
    LocalMux I__5351 (
            .O(N__21868),
            .I(M_this_external_address_qZ0Z_14));
    InMux I__5350 (
            .O(N__21863),
            .I(un1_M_this_external_address_q_cry_13));
    InMux I__5349 (
            .O(N__21860),
            .I(N__21830));
    InMux I__5348 (
            .O(N__21859),
            .I(N__21830));
    InMux I__5347 (
            .O(N__21858),
            .I(N__21821));
    InMux I__5346 (
            .O(N__21857),
            .I(N__21821));
    InMux I__5345 (
            .O(N__21856),
            .I(N__21821));
    InMux I__5344 (
            .O(N__21855),
            .I(N__21821));
    InMux I__5343 (
            .O(N__21854),
            .I(N__21810));
    InMux I__5342 (
            .O(N__21853),
            .I(N__21810));
    InMux I__5341 (
            .O(N__21852),
            .I(N__21810));
    InMux I__5340 (
            .O(N__21851),
            .I(N__21810));
    InMux I__5339 (
            .O(N__21850),
            .I(N__21801));
    InMux I__5338 (
            .O(N__21849),
            .I(N__21801));
    InMux I__5337 (
            .O(N__21848),
            .I(N__21801));
    InMux I__5336 (
            .O(N__21847),
            .I(N__21801));
    InMux I__5335 (
            .O(N__21846),
            .I(N__21792));
    InMux I__5334 (
            .O(N__21845),
            .I(N__21792));
    InMux I__5333 (
            .O(N__21844),
            .I(N__21792));
    InMux I__5332 (
            .O(N__21843),
            .I(N__21792));
    InMux I__5331 (
            .O(N__21842),
            .I(N__21783));
    InMux I__5330 (
            .O(N__21841),
            .I(N__21783));
    InMux I__5329 (
            .O(N__21840),
            .I(N__21783));
    InMux I__5328 (
            .O(N__21839),
            .I(N__21783));
    InMux I__5327 (
            .O(N__21838),
            .I(N__21775));
    InMux I__5326 (
            .O(N__21837),
            .I(N__21775));
    InMux I__5325 (
            .O(N__21836),
            .I(N__21775));
    InMux I__5324 (
            .O(N__21835),
            .I(N__21772));
    LocalMux I__5323 (
            .O(N__21830),
            .I(N__21767));
    LocalMux I__5322 (
            .O(N__21821),
            .I(N__21767));
    InMux I__5321 (
            .O(N__21820),
            .I(N__21762));
    InMux I__5320 (
            .O(N__21819),
            .I(N__21762));
    LocalMux I__5319 (
            .O(N__21810),
            .I(N__21758));
    LocalMux I__5318 (
            .O(N__21801),
            .I(N__21751));
    LocalMux I__5317 (
            .O(N__21792),
            .I(N__21751));
    LocalMux I__5316 (
            .O(N__21783),
            .I(N__21751));
    InMux I__5315 (
            .O(N__21782),
            .I(N__21748));
    LocalMux I__5314 (
            .O(N__21775),
            .I(N__21743));
    LocalMux I__5313 (
            .O(N__21772),
            .I(N__21736));
    Span4Mux_v I__5312 (
            .O(N__21767),
            .I(N__21736));
    LocalMux I__5311 (
            .O(N__21762),
            .I(N__21736));
    InMux I__5310 (
            .O(N__21761),
            .I(N__21733));
    Span4Mux_v I__5309 (
            .O(N__21758),
            .I(N__21728));
    Span4Mux_v I__5308 (
            .O(N__21751),
            .I(N__21728));
    LocalMux I__5307 (
            .O(N__21748),
            .I(N__21724));
    InMux I__5306 (
            .O(N__21747),
            .I(N__21719));
    InMux I__5305 (
            .O(N__21746),
            .I(N__21719));
    Span4Mux_v I__5304 (
            .O(N__21743),
            .I(N__21714));
    Span4Mux_v I__5303 (
            .O(N__21736),
            .I(N__21711));
    LocalMux I__5302 (
            .O(N__21733),
            .I(N__21706));
    Sp12to4 I__5301 (
            .O(N__21728),
            .I(N__21706));
    InMux I__5300 (
            .O(N__21727),
            .I(N__21703));
    Span4Mux_h I__5299 (
            .O(N__21724),
            .I(N__21698));
    LocalMux I__5298 (
            .O(N__21719),
            .I(N__21698));
    InMux I__5297 (
            .O(N__21718),
            .I(N__21693));
    InMux I__5296 (
            .O(N__21717),
            .I(N__21693));
    Odrv4 I__5295 (
            .O(N__21714),
            .I(M_this_state_qZ0Z_0));
    Odrv4 I__5294 (
            .O(N__21711),
            .I(M_this_state_qZ0Z_0));
    Odrv12 I__5293 (
            .O(N__21706),
            .I(M_this_state_qZ0Z_0));
    LocalMux I__5292 (
            .O(N__21703),
            .I(M_this_state_qZ0Z_0));
    Odrv4 I__5291 (
            .O(N__21698),
            .I(M_this_state_qZ0Z_0));
    LocalMux I__5290 (
            .O(N__21693),
            .I(M_this_state_qZ0Z_0));
    InMux I__5289 (
            .O(N__21680),
            .I(un1_M_this_external_address_q_cry_14));
    IoInMux I__5288 (
            .O(N__21677),
            .I(N__21674));
    LocalMux I__5287 (
            .O(N__21674),
            .I(N__21671));
    Span4Mux_s2_h I__5286 (
            .O(N__21671),
            .I(N__21668));
    Sp12to4 I__5285 (
            .O(N__21668),
            .I(N__21665));
    Span12Mux_v I__5284 (
            .O(N__21665),
            .I(N__21661));
    InMux I__5283 (
            .O(N__21664),
            .I(N__21658));
    Odrv12 I__5282 (
            .O(N__21661),
            .I(M_this_external_address_qZ0Z_15));
    LocalMux I__5281 (
            .O(N__21658),
            .I(M_this_external_address_qZ0Z_15));
    ClkMux I__5280 (
            .O(N__21653),
            .I(N__21401));
    ClkMux I__5279 (
            .O(N__21652),
            .I(N__21401));
    ClkMux I__5278 (
            .O(N__21651),
            .I(N__21401));
    ClkMux I__5277 (
            .O(N__21650),
            .I(N__21401));
    ClkMux I__5276 (
            .O(N__21649),
            .I(N__21401));
    ClkMux I__5275 (
            .O(N__21648),
            .I(N__21401));
    ClkMux I__5274 (
            .O(N__21647),
            .I(N__21401));
    ClkMux I__5273 (
            .O(N__21646),
            .I(N__21401));
    ClkMux I__5272 (
            .O(N__21645),
            .I(N__21401));
    ClkMux I__5271 (
            .O(N__21644),
            .I(N__21401));
    ClkMux I__5270 (
            .O(N__21643),
            .I(N__21401));
    ClkMux I__5269 (
            .O(N__21642),
            .I(N__21401));
    ClkMux I__5268 (
            .O(N__21641),
            .I(N__21401));
    ClkMux I__5267 (
            .O(N__21640),
            .I(N__21401));
    ClkMux I__5266 (
            .O(N__21639),
            .I(N__21401));
    ClkMux I__5265 (
            .O(N__21638),
            .I(N__21401));
    ClkMux I__5264 (
            .O(N__21637),
            .I(N__21401));
    ClkMux I__5263 (
            .O(N__21636),
            .I(N__21401));
    ClkMux I__5262 (
            .O(N__21635),
            .I(N__21401));
    ClkMux I__5261 (
            .O(N__21634),
            .I(N__21401));
    ClkMux I__5260 (
            .O(N__21633),
            .I(N__21401));
    ClkMux I__5259 (
            .O(N__21632),
            .I(N__21401));
    ClkMux I__5258 (
            .O(N__21631),
            .I(N__21401));
    ClkMux I__5257 (
            .O(N__21630),
            .I(N__21401));
    ClkMux I__5256 (
            .O(N__21629),
            .I(N__21401));
    ClkMux I__5255 (
            .O(N__21628),
            .I(N__21401));
    ClkMux I__5254 (
            .O(N__21627),
            .I(N__21401));
    ClkMux I__5253 (
            .O(N__21626),
            .I(N__21401));
    ClkMux I__5252 (
            .O(N__21625),
            .I(N__21401));
    ClkMux I__5251 (
            .O(N__21624),
            .I(N__21401));
    ClkMux I__5250 (
            .O(N__21623),
            .I(N__21401));
    ClkMux I__5249 (
            .O(N__21622),
            .I(N__21401));
    ClkMux I__5248 (
            .O(N__21621),
            .I(N__21401));
    ClkMux I__5247 (
            .O(N__21620),
            .I(N__21401));
    ClkMux I__5246 (
            .O(N__21619),
            .I(N__21401));
    ClkMux I__5245 (
            .O(N__21618),
            .I(N__21401));
    ClkMux I__5244 (
            .O(N__21617),
            .I(N__21401));
    ClkMux I__5243 (
            .O(N__21616),
            .I(N__21401));
    ClkMux I__5242 (
            .O(N__21615),
            .I(N__21401));
    ClkMux I__5241 (
            .O(N__21614),
            .I(N__21401));
    ClkMux I__5240 (
            .O(N__21613),
            .I(N__21401));
    ClkMux I__5239 (
            .O(N__21612),
            .I(N__21401));
    ClkMux I__5238 (
            .O(N__21611),
            .I(N__21401));
    ClkMux I__5237 (
            .O(N__21610),
            .I(N__21401));
    ClkMux I__5236 (
            .O(N__21609),
            .I(N__21401));
    ClkMux I__5235 (
            .O(N__21608),
            .I(N__21401));
    ClkMux I__5234 (
            .O(N__21607),
            .I(N__21401));
    ClkMux I__5233 (
            .O(N__21606),
            .I(N__21401));
    ClkMux I__5232 (
            .O(N__21605),
            .I(N__21401));
    ClkMux I__5231 (
            .O(N__21604),
            .I(N__21401));
    ClkMux I__5230 (
            .O(N__21603),
            .I(N__21401));
    ClkMux I__5229 (
            .O(N__21602),
            .I(N__21401));
    ClkMux I__5228 (
            .O(N__21601),
            .I(N__21401));
    ClkMux I__5227 (
            .O(N__21600),
            .I(N__21401));
    ClkMux I__5226 (
            .O(N__21599),
            .I(N__21401));
    ClkMux I__5225 (
            .O(N__21598),
            .I(N__21401));
    ClkMux I__5224 (
            .O(N__21597),
            .I(N__21401));
    ClkMux I__5223 (
            .O(N__21596),
            .I(N__21401));
    ClkMux I__5222 (
            .O(N__21595),
            .I(N__21401));
    ClkMux I__5221 (
            .O(N__21594),
            .I(N__21401));
    ClkMux I__5220 (
            .O(N__21593),
            .I(N__21401));
    ClkMux I__5219 (
            .O(N__21592),
            .I(N__21401));
    ClkMux I__5218 (
            .O(N__21591),
            .I(N__21401));
    ClkMux I__5217 (
            .O(N__21590),
            .I(N__21401));
    ClkMux I__5216 (
            .O(N__21589),
            .I(N__21401));
    ClkMux I__5215 (
            .O(N__21588),
            .I(N__21401));
    ClkMux I__5214 (
            .O(N__21587),
            .I(N__21401));
    ClkMux I__5213 (
            .O(N__21586),
            .I(N__21401));
    ClkMux I__5212 (
            .O(N__21585),
            .I(N__21401));
    ClkMux I__5211 (
            .O(N__21584),
            .I(N__21401));
    ClkMux I__5210 (
            .O(N__21583),
            .I(N__21401));
    ClkMux I__5209 (
            .O(N__21582),
            .I(N__21401));
    ClkMux I__5208 (
            .O(N__21581),
            .I(N__21401));
    ClkMux I__5207 (
            .O(N__21580),
            .I(N__21401));
    ClkMux I__5206 (
            .O(N__21579),
            .I(N__21401));
    ClkMux I__5205 (
            .O(N__21578),
            .I(N__21401));
    ClkMux I__5204 (
            .O(N__21577),
            .I(N__21401));
    ClkMux I__5203 (
            .O(N__21576),
            .I(N__21401));
    ClkMux I__5202 (
            .O(N__21575),
            .I(N__21401));
    ClkMux I__5201 (
            .O(N__21574),
            .I(N__21401));
    ClkMux I__5200 (
            .O(N__21573),
            .I(N__21401));
    ClkMux I__5199 (
            .O(N__21572),
            .I(N__21401));
    ClkMux I__5198 (
            .O(N__21571),
            .I(N__21401));
    ClkMux I__5197 (
            .O(N__21570),
            .I(N__21401));
    GlobalMux I__5196 (
            .O(N__21401),
            .I(N__21398));
    gio2CtrlBuf I__5195 (
            .O(N__21398),
            .I(clk_0_c_g));
    InMux I__5194 (
            .O(N__21395),
            .I(N__21381));
    InMux I__5193 (
            .O(N__21394),
            .I(N__21378));
    InMux I__5192 (
            .O(N__21393),
            .I(N__21375));
    InMux I__5191 (
            .O(N__21392),
            .I(N__21372));
    InMux I__5190 (
            .O(N__21391),
            .I(N__21369));
    InMux I__5189 (
            .O(N__21390),
            .I(N__21366));
    InMux I__5188 (
            .O(N__21389),
            .I(N__21359));
    InMux I__5187 (
            .O(N__21388),
            .I(N__21359));
    InMux I__5186 (
            .O(N__21387),
            .I(N__21359));
    InMux I__5185 (
            .O(N__21386),
            .I(N__21354));
    InMux I__5184 (
            .O(N__21385),
            .I(N__21354));
    InMux I__5183 (
            .O(N__21384),
            .I(N__21351));
    LocalMux I__5182 (
            .O(N__21381),
            .I(N__21337));
    LocalMux I__5181 (
            .O(N__21378),
            .I(N__21334));
    LocalMux I__5180 (
            .O(N__21375),
            .I(N__21331));
    LocalMux I__5179 (
            .O(N__21372),
            .I(N__21328));
    LocalMux I__5178 (
            .O(N__21369),
            .I(N__21325));
    LocalMux I__5177 (
            .O(N__21366),
            .I(N__21322));
    LocalMux I__5176 (
            .O(N__21359),
            .I(N__21319));
    LocalMux I__5175 (
            .O(N__21354),
            .I(N__21316));
    LocalMux I__5174 (
            .O(N__21351),
            .I(N__21313));
    SRMux I__5173 (
            .O(N__21350),
            .I(N__21272));
    SRMux I__5172 (
            .O(N__21349),
            .I(N__21272));
    SRMux I__5171 (
            .O(N__21348),
            .I(N__21272));
    SRMux I__5170 (
            .O(N__21347),
            .I(N__21272));
    SRMux I__5169 (
            .O(N__21346),
            .I(N__21272));
    SRMux I__5168 (
            .O(N__21345),
            .I(N__21272));
    SRMux I__5167 (
            .O(N__21344),
            .I(N__21272));
    SRMux I__5166 (
            .O(N__21343),
            .I(N__21272));
    SRMux I__5165 (
            .O(N__21342),
            .I(N__21272));
    SRMux I__5164 (
            .O(N__21341),
            .I(N__21272));
    SRMux I__5163 (
            .O(N__21340),
            .I(N__21272));
    Glb2LocalMux I__5162 (
            .O(N__21337),
            .I(N__21272));
    Glb2LocalMux I__5161 (
            .O(N__21334),
            .I(N__21272));
    Glb2LocalMux I__5160 (
            .O(N__21331),
            .I(N__21272));
    Glb2LocalMux I__5159 (
            .O(N__21328),
            .I(N__21272));
    Glb2LocalMux I__5158 (
            .O(N__21325),
            .I(N__21272));
    Glb2LocalMux I__5157 (
            .O(N__21322),
            .I(N__21272));
    Glb2LocalMux I__5156 (
            .O(N__21319),
            .I(N__21272));
    Glb2LocalMux I__5155 (
            .O(N__21316),
            .I(N__21272));
    Glb2LocalMux I__5154 (
            .O(N__21313),
            .I(N__21272));
    GlobalMux I__5153 (
            .O(N__21272),
            .I(N__21269));
    gio2CtrlBuf I__5152 (
            .O(N__21269),
            .I(M_this_state_q_nss_g_0));
    InMux I__5151 (
            .O(N__21266),
            .I(N__21263));
    LocalMux I__5150 (
            .O(N__21263),
            .I(N__21260));
    Span4Mux_v I__5149 (
            .O(N__21260),
            .I(N__21257));
    Odrv4 I__5148 (
            .O(N__21257),
            .I(port_address_in_5));
    InMux I__5147 (
            .O(N__21254),
            .I(N__21251));
    LocalMux I__5146 (
            .O(N__21251),
            .I(N__21248));
    Span12Mux_v I__5145 (
            .O(N__21248),
            .I(N__21245));
    Odrv12 I__5144 (
            .O(N__21245),
            .I(port_address_in_6));
    CascadeMux I__5143 (
            .O(N__21242),
            .I(N__21239));
    InMux I__5142 (
            .O(N__21239),
            .I(N__21236));
    LocalMux I__5141 (
            .O(N__21236),
            .I(N__21233));
    Span4Mux_v I__5140 (
            .O(N__21233),
            .I(N__21230));
    Span4Mux_v I__5139 (
            .O(N__21230),
            .I(N__21227));
    Span4Mux_v I__5138 (
            .O(N__21227),
            .I(N__21224));
    Span4Mux_v I__5137 (
            .O(N__21224),
            .I(N__21221));
    Odrv4 I__5136 (
            .O(N__21221),
            .I(port_address_in_7));
    InMux I__5135 (
            .O(N__21218),
            .I(N__21215));
    LocalMux I__5134 (
            .O(N__21215),
            .I(N__21212));
    IoSpan4Mux I__5133 (
            .O(N__21212),
            .I(N__21209));
    Odrv4 I__5132 (
            .O(N__21209),
            .I(port_address_in_4));
    CascadeMux I__5131 (
            .O(N__21206),
            .I(N__21202));
    CascadeMux I__5130 (
            .O(N__21205),
            .I(N__21198));
    InMux I__5129 (
            .O(N__21202),
            .I(N__21188));
    InMux I__5128 (
            .O(N__21201),
            .I(N__21188));
    InMux I__5127 (
            .O(N__21198),
            .I(N__21188));
    InMux I__5126 (
            .O(N__21197),
            .I(N__21188));
    LocalMux I__5125 (
            .O(N__21188),
            .I(N__21185));
    Span12Mux_v I__5124 (
            .O(N__21185),
            .I(N__21182));
    Span12Mux_h I__5123 (
            .O(N__21182),
            .I(N__21179));
    Odrv12 I__5122 (
            .O(N__21179),
            .I(\this_start_data_delay.M_this_state_d27Z0Z_6 ));
    InMux I__5121 (
            .O(N__21176),
            .I(un1_M_this_external_address_q_cry_3));
    IoInMux I__5120 (
            .O(N__21173),
            .I(N__21170));
    LocalMux I__5119 (
            .O(N__21170),
            .I(N__21167));
    Span4Mux_s2_h I__5118 (
            .O(N__21167),
            .I(N__21163));
    InMux I__5117 (
            .O(N__21166),
            .I(N__21160));
    Odrv4 I__5116 (
            .O(N__21163),
            .I(M_this_external_address_qZ0Z_5));
    LocalMux I__5115 (
            .O(N__21160),
            .I(M_this_external_address_qZ0Z_5));
    InMux I__5114 (
            .O(N__21155),
            .I(un1_M_this_external_address_q_cry_4));
    IoInMux I__5113 (
            .O(N__21152),
            .I(N__21149));
    LocalMux I__5112 (
            .O(N__21149),
            .I(N__21146));
    Span12Mux_s2_h I__5111 (
            .O(N__21146),
            .I(N__21142));
    InMux I__5110 (
            .O(N__21145),
            .I(N__21139));
    Odrv12 I__5109 (
            .O(N__21142),
            .I(M_this_external_address_qZ0Z_6));
    LocalMux I__5108 (
            .O(N__21139),
            .I(M_this_external_address_qZ0Z_6));
    InMux I__5107 (
            .O(N__21134),
            .I(un1_M_this_external_address_q_cry_5));
    IoInMux I__5106 (
            .O(N__21131),
            .I(N__21128));
    LocalMux I__5105 (
            .O(N__21128),
            .I(N__21125));
    Span4Mux_s2_h I__5104 (
            .O(N__21125),
            .I(N__21122));
    Sp12to4 I__5103 (
            .O(N__21122),
            .I(N__21119));
    Span12Mux_v I__5102 (
            .O(N__21119),
            .I(N__21115));
    InMux I__5101 (
            .O(N__21118),
            .I(N__21112));
    Odrv12 I__5100 (
            .O(N__21115),
            .I(M_this_external_address_qZ0Z_7));
    LocalMux I__5099 (
            .O(N__21112),
            .I(M_this_external_address_qZ0Z_7));
    InMux I__5098 (
            .O(N__21107),
            .I(un1_M_this_external_address_q_cry_6));
    IoInMux I__5097 (
            .O(N__21104),
            .I(N__21101));
    LocalMux I__5096 (
            .O(N__21101),
            .I(N__21098));
    IoSpan4Mux I__5095 (
            .O(N__21098),
            .I(N__21095));
    Span4Mux_s2_v I__5094 (
            .O(N__21095),
            .I(N__21092));
    Sp12to4 I__5093 (
            .O(N__21092),
            .I(N__21089));
    Span12Mux_s8_v I__5092 (
            .O(N__21089),
            .I(N__21086));
    Span12Mux_h I__5091 (
            .O(N__21086),
            .I(N__21082));
    InMux I__5090 (
            .O(N__21085),
            .I(N__21079));
    Odrv12 I__5089 (
            .O(N__21082),
            .I(M_this_external_address_qZ0Z_8));
    LocalMux I__5088 (
            .O(N__21079),
            .I(M_this_external_address_qZ0Z_8));
    InMux I__5087 (
            .O(N__21074),
            .I(bfn_30_24_0_));
    IoInMux I__5086 (
            .O(N__21071),
            .I(N__21068));
    LocalMux I__5085 (
            .O(N__21068),
            .I(N__21065));
    Span12Mux_s8_v I__5084 (
            .O(N__21065),
            .I(N__21061));
    InMux I__5083 (
            .O(N__21064),
            .I(N__21058));
    Odrv12 I__5082 (
            .O(N__21061),
            .I(M_this_external_address_qZ0Z_9));
    LocalMux I__5081 (
            .O(N__21058),
            .I(M_this_external_address_qZ0Z_9));
    InMux I__5080 (
            .O(N__21053),
            .I(un1_M_this_external_address_q_cry_8));
    IoInMux I__5079 (
            .O(N__21050),
            .I(N__21047));
    LocalMux I__5078 (
            .O(N__21047),
            .I(N__21044));
    Span4Mux_s2_v I__5077 (
            .O(N__21044),
            .I(N__21041));
    Span4Mux_h I__5076 (
            .O(N__21041),
            .I(N__21038));
    Sp12to4 I__5075 (
            .O(N__21038),
            .I(N__21035));
    Span12Mux_s8_v I__5074 (
            .O(N__21035),
            .I(N__21031));
    InMux I__5073 (
            .O(N__21034),
            .I(N__21028));
    Odrv12 I__5072 (
            .O(N__21031),
            .I(M_this_external_address_qZ0Z_10));
    LocalMux I__5071 (
            .O(N__21028),
            .I(M_this_external_address_qZ0Z_10));
    InMux I__5070 (
            .O(N__21023),
            .I(un1_M_this_external_address_q_cry_9));
    IoInMux I__5069 (
            .O(N__21020),
            .I(N__21017));
    LocalMux I__5068 (
            .O(N__21017),
            .I(N__21013));
    InMux I__5067 (
            .O(N__21016),
            .I(N__21010));
    Odrv12 I__5066 (
            .O(N__21013),
            .I(M_this_external_address_qZ0Z_11));
    LocalMux I__5065 (
            .O(N__21010),
            .I(M_this_external_address_qZ0Z_11));
    InMux I__5064 (
            .O(N__21005),
            .I(un1_M_this_external_address_q_cry_10));
    IoInMux I__5063 (
            .O(N__21002),
            .I(N__20999));
    LocalMux I__5062 (
            .O(N__20999),
            .I(N__20995));
    InMux I__5061 (
            .O(N__20998),
            .I(N__20992));
    Odrv4 I__5060 (
            .O(N__20995),
            .I(M_this_external_address_qZ0Z_12));
    LocalMux I__5059 (
            .O(N__20992),
            .I(M_this_external_address_qZ0Z_12));
    InMux I__5058 (
            .O(N__20987),
            .I(un1_M_this_external_address_q_cry_11));
    CascadeMux I__5057 (
            .O(N__20984),
            .I(N__20981));
    InMux I__5056 (
            .O(N__20981),
            .I(N__20978));
    LocalMux I__5055 (
            .O(N__20978),
            .I(N__20974));
    CascadeMux I__5054 (
            .O(N__20977),
            .I(N__20971));
    Span4Mux_h I__5053 (
            .O(N__20974),
            .I(N__20967));
    InMux I__5052 (
            .O(N__20971),
            .I(N__20964));
    InMux I__5051 (
            .O(N__20970),
            .I(N__20961));
    Span4Mux_h I__5050 (
            .O(N__20967),
            .I(N__20958));
    LocalMux I__5049 (
            .O(N__20964),
            .I(N__20953));
    LocalMux I__5048 (
            .O(N__20961),
            .I(N__20953));
    Sp12to4 I__5047 (
            .O(N__20958),
            .I(N__20950));
    Span12Mux_h I__5046 (
            .O(N__20953),
            .I(N__20947));
    Odrv12 I__5045 (
            .O(N__20950),
            .I(port_data_c_2));
    Odrv12 I__5044 (
            .O(N__20947),
            .I(port_data_c_2));
    CascadeMux I__5043 (
            .O(N__20942),
            .I(N__20939));
    InMux I__5042 (
            .O(N__20939),
            .I(N__20935));
    CascadeMux I__5041 (
            .O(N__20938),
            .I(N__20932));
    LocalMux I__5040 (
            .O(N__20935),
            .I(N__20929));
    InMux I__5039 (
            .O(N__20932),
            .I(N__20926));
    Span4Mux_h I__5038 (
            .O(N__20929),
            .I(N__20921));
    LocalMux I__5037 (
            .O(N__20926),
            .I(N__20921));
    Span4Mux_h I__5036 (
            .O(N__20921),
            .I(N__20917));
    InMux I__5035 (
            .O(N__20920),
            .I(N__20914));
    Sp12to4 I__5034 (
            .O(N__20917),
            .I(N__20909));
    LocalMux I__5033 (
            .O(N__20914),
            .I(N__20909));
    Span12Mux_v I__5032 (
            .O(N__20909),
            .I(N__20906));
    Odrv12 I__5031 (
            .O(N__20906),
            .I(port_data_c_6));
    CascadeMux I__5030 (
            .O(N__20903),
            .I(N__20898));
    InMux I__5029 (
            .O(N__20902),
            .I(N__20895));
    InMux I__5028 (
            .O(N__20901),
            .I(N__20892));
    InMux I__5027 (
            .O(N__20898),
            .I(N__20889));
    LocalMux I__5026 (
            .O(N__20895),
            .I(N__20886));
    LocalMux I__5025 (
            .O(N__20892),
            .I(M_this_vram_write_data_0_sqmuxa));
    LocalMux I__5024 (
            .O(N__20889),
            .I(M_this_vram_write_data_0_sqmuxa));
    Odrv4 I__5023 (
            .O(N__20886),
            .I(M_this_vram_write_data_0_sqmuxa));
    InMux I__5022 (
            .O(N__20879),
            .I(N__20873));
    InMux I__5021 (
            .O(N__20878),
            .I(N__20870));
    InMux I__5020 (
            .O(N__20877),
            .I(N__20867));
    InMux I__5019 (
            .O(N__20876),
            .I(N__20864));
    LocalMux I__5018 (
            .O(N__20873),
            .I(\this_start_data_delay.un1_M_this_state_q_0 ));
    LocalMux I__5017 (
            .O(N__20870),
            .I(\this_start_data_delay.un1_M_this_state_q_0 ));
    LocalMux I__5016 (
            .O(N__20867),
            .I(\this_start_data_delay.un1_M_this_state_q_0 ));
    LocalMux I__5015 (
            .O(N__20864),
            .I(\this_start_data_delay.un1_M_this_state_q_0 ));
    InMux I__5014 (
            .O(N__20855),
            .I(N__20852));
    LocalMux I__5013 (
            .O(N__20852),
            .I(N__20848));
    InMux I__5012 (
            .O(N__20851),
            .I(N__20845));
    Span4Mux_v I__5011 (
            .O(N__20848),
            .I(N__20838));
    LocalMux I__5010 (
            .O(N__20845),
            .I(N__20838));
    InMux I__5009 (
            .O(N__20844),
            .I(N__20835));
    InMux I__5008 (
            .O(N__20843),
            .I(N__20831));
    Span4Mux_v I__5007 (
            .O(N__20838),
            .I(N__20825));
    LocalMux I__5006 (
            .O(N__20835),
            .I(N__20825));
    InMux I__5005 (
            .O(N__20834),
            .I(N__20822));
    LocalMux I__5004 (
            .O(N__20831),
            .I(N__20819));
    InMux I__5003 (
            .O(N__20830),
            .I(N__20816));
    Span4Mux_v I__5002 (
            .O(N__20825),
            .I(N__20810));
    LocalMux I__5001 (
            .O(N__20822),
            .I(N__20810));
    Span4Mux_v I__5000 (
            .O(N__20819),
            .I(N__20805));
    LocalMux I__4999 (
            .O(N__20816),
            .I(N__20805));
    InMux I__4998 (
            .O(N__20815),
            .I(N__20802));
    Span4Mux_v I__4997 (
            .O(N__20810),
            .I(N__20798));
    Span4Mux_v I__4996 (
            .O(N__20805),
            .I(N__20793));
    LocalMux I__4995 (
            .O(N__20802),
            .I(N__20793));
    InMux I__4994 (
            .O(N__20801),
            .I(N__20790));
    Odrv4 I__4993 (
            .O(N__20798),
            .I(M_this_vram_write_data_0_i_2));
    Odrv4 I__4992 (
            .O(N__20793),
            .I(M_this_vram_write_data_0_i_2));
    LocalMux I__4991 (
            .O(N__20790),
            .I(M_this_vram_write_data_0_i_2));
    CEMux I__4990 (
            .O(N__20783),
            .I(N__20779));
    CEMux I__4989 (
            .O(N__20782),
            .I(N__20776));
    LocalMux I__4988 (
            .O(N__20779),
            .I(N__20771));
    LocalMux I__4987 (
            .O(N__20776),
            .I(N__20771));
    Span4Mux_s3_v I__4986 (
            .O(N__20771),
            .I(N__20768));
    Span4Mux_v I__4985 (
            .O(N__20768),
            .I(N__20765));
    Odrv4 I__4984 (
            .O(N__20765),
            .I(\this_vram.mem_WE_0 ));
    InMux I__4983 (
            .O(N__20762),
            .I(N__20752));
    InMux I__4982 (
            .O(N__20761),
            .I(N__20752));
    InMux I__4981 (
            .O(N__20760),
            .I(N__20752));
    InMux I__4980 (
            .O(N__20759),
            .I(N__20746));
    LocalMux I__4979 (
            .O(N__20752),
            .I(N__20743));
    InMux I__4978 (
            .O(N__20751),
            .I(N__20740));
    InMux I__4977 (
            .O(N__20750),
            .I(N__20735));
    InMux I__4976 (
            .O(N__20749),
            .I(N__20735));
    LocalMux I__4975 (
            .O(N__20746),
            .I(N__20731));
    Span4Mux_v I__4974 (
            .O(N__20743),
            .I(N__20725));
    LocalMux I__4973 (
            .O(N__20740),
            .I(N__20725));
    LocalMux I__4972 (
            .O(N__20735),
            .I(N__20722));
    InMux I__4971 (
            .O(N__20734),
            .I(N__20719));
    Span4Mux_v I__4970 (
            .O(N__20731),
            .I(N__20716));
    InMux I__4969 (
            .O(N__20730),
            .I(N__20713));
    Span4Mux_h I__4968 (
            .O(N__20725),
            .I(N__20707));
    Span4Mux_h I__4967 (
            .O(N__20722),
            .I(N__20707));
    LocalMux I__4966 (
            .O(N__20719),
            .I(N__20704));
    Span4Mux_v I__4965 (
            .O(N__20716),
            .I(N__20699));
    LocalMux I__4964 (
            .O(N__20713),
            .I(N__20699));
    InMux I__4963 (
            .O(N__20712),
            .I(N__20696));
    Odrv4 I__4962 (
            .O(N__20707),
            .I(M_this_internal_address_qZ0Z_12));
    Odrv4 I__4961 (
            .O(N__20704),
            .I(M_this_internal_address_qZ0Z_12));
    Odrv4 I__4960 (
            .O(N__20699),
            .I(M_this_internal_address_qZ0Z_12));
    LocalMux I__4959 (
            .O(N__20696),
            .I(M_this_internal_address_qZ0Z_12));
    CascadeMux I__4958 (
            .O(N__20687),
            .I(N__20682));
    CascadeMux I__4957 (
            .O(N__20686),
            .I(N__20676));
    InMux I__4956 (
            .O(N__20685),
            .I(N__20672));
    InMux I__4955 (
            .O(N__20682),
            .I(N__20665));
    InMux I__4954 (
            .O(N__20681),
            .I(N__20665));
    InMux I__4953 (
            .O(N__20680),
            .I(N__20665));
    InMux I__4952 (
            .O(N__20679),
            .I(N__20660));
    InMux I__4951 (
            .O(N__20676),
            .I(N__20655));
    InMux I__4950 (
            .O(N__20675),
            .I(N__20655));
    LocalMux I__4949 (
            .O(N__20672),
            .I(N__20650));
    LocalMux I__4948 (
            .O(N__20665),
            .I(N__20650));
    CascadeMux I__4947 (
            .O(N__20664),
            .I(N__20647));
    InMux I__4946 (
            .O(N__20663),
            .I(N__20644));
    LocalMux I__4945 (
            .O(N__20660),
            .I(N__20641));
    LocalMux I__4944 (
            .O(N__20655),
            .I(N__20638));
    Span4Mux_h I__4943 (
            .O(N__20650),
            .I(N__20635));
    InMux I__4942 (
            .O(N__20647),
            .I(N__20631));
    LocalMux I__4941 (
            .O(N__20644),
            .I(N__20628));
    Span4Mux_v I__4940 (
            .O(N__20641),
            .I(N__20623));
    Span4Mux_v I__4939 (
            .O(N__20638),
            .I(N__20623));
    Span4Mux_v I__4938 (
            .O(N__20635),
            .I(N__20620));
    InMux I__4937 (
            .O(N__20634),
            .I(N__20617));
    LocalMux I__4936 (
            .O(N__20631),
            .I(N__20614));
    Span4Mux_v I__4935 (
            .O(N__20628),
            .I(N__20609));
    Span4Mux_h I__4934 (
            .O(N__20623),
            .I(N__20609));
    Span4Mux_h I__4933 (
            .O(N__20620),
            .I(N__20606));
    LocalMux I__4932 (
            .O(N__20617),
            .I(M_this_internal_address_qZ0Z_11));
    Odrv12 I__4931 (
            .O(N__20614),
            .I(M_this_internal_address_qZ0Z_11));
    Odrv4 I__4930 (
            .O(N__20609),
            .I(M_this_internal_address_qZ0Z_11));
    Odrv4 I__4929 (
            .O(N__20606),
            .I(M_this_internal_address_qZ0Z_11));
    CascadeMux I__4928 (
            .O(N__20597),
            .I(N__20591));
    CascadeMux I__4927 (
            .O(N__20596),
            .I(N__20587));
    CascadeMux I__4926 (
            .O(N__20595),
            .I(N__20584));
    CascadeMux I__4925 (
            .O(N__20594),
            .I(N__20581));
    InMux I__4924 (
            .O(N__20591),
            .I(N__20574));
    InMux I__4923 (
            .O(N__20590),
            .I(N__20574));
    InMux I__4922 (
            .O(N__20587),
            .I(N__20574));
    InMux I__4921 (
            .O(N__20584),
            .I(N__20571));
    InMux I__4920 (
            .O(N__20581),
            .I(N__20568));
    LocalMux I__4919 (
            .O(N__20574),
            .I(N__20561));
    LocalMux I__4918 (
            .O(N__20571),
            .I(N__20561));
    LocalMux I__4917 (
            .O(N__20568),
            .I(N__20558));
    InMux I__4916 (
            .O(N__20567),
            .I(N__20555));
    CascadeMux I__4915 (
            .O(N__20566),
            .I(N__20551));
    Span4Mux_v I__4914 (
            .O(N__20561),
            .I(N__20543));
    Span4Mux_h I__4913 (
            .O(N__20558),
            .I(N__20543));
    LocalMux I__4912 (
            .O(N__20555),
            .I(N__20543));
    InMux I__4911 (
            .O(N__20554),
            .I(N__20538));
    InMux I__4910 (
            .O(N__20551),
            .I(N__20538));
    InMux I__4909 (
            .O(N__20550),
            .I(N__20535));
    Span4Mux_v I__4908 (
            .O(N__20543),
            .I(N__20530));
    LocalMux I__4907 (
            .O(N__20538),
            .I(N__20530));
    LocalMux I__4906 (
            .O(N__20535),
            .I(N__20527));
    Span4Mux_h I__4905 (
            .O(N__20530),
            .I(N__20521));
    Span4Mux_v I__4904 (
            .O(N__20527),
            .I(N__20521));
    InMux I__4903 (
            .O(N__20526),
            .I(N__20518));
    Odrv4 I__4902 (
            .O(N__20521),
            .I(M_this_internal_address_qZ0Z_13));
    LocalMux I__4901 (
            .O(N__20518),
            .I(M_this_internal_address_qZ0Z_13));
    InMux I__4900 (
            .O(N__20513),
            .I(N__20503));
    InMux I__4899 (
            .O(N__20512),
            .I(N__20503));
    InMux I__4898 (
            .O(N__20511),
            .I(N__20503));
    InMux I__4897 (
            .O(N__20510),
            .I(N__20499));
    LocalMux I__4896 (
            .O(N__20503),
            .I(N__20496));
    InMux I__4895 (
            .O(N__20502),
            .I(N__20493));
    LocalMux I__4894 (
            .O(N__20499),
            .I(N__20490));
    Span4Mux_v I__4893 (
            .O(N__20496),
            .I(N__20484));
    LocalMux I__4892 (
            .O(N__20493),
            .I(N__20481));
    Span4Mux_h I__4891 (
            .O(N__20490),
            .I(N__20478));
    InMux I__4890 (
            .O(N__20489),
            .I(N__20475));
    InMux I__4889 (
            .O(N__20488),
            .I(N__20470));
    InMux I__4888 (
            .O(N__20487),
            .I(N__20470));
    Odrv4 I__4887 (
            .O(N__20484),
            .I(M_this_vram_write_en_0_0));
    Odrv12 I__4886 (
            .O(N__20481),
            .I(M_this_vram_write_en_0_0));
    Odrv4 I__4885 (
            .O(N__20478),
            .I(M_this_vram_write_en_0_0));
    LocalMux I__4884 (
            .O(N__20475),
            .I(M_this_vram_write_en_0_0));
    LocalMux I__4883 (
            .O(N__20470),
            .I(M_this_vram_write_en_0_0));
    CEMux I__4882 (
            .O(N__20459),
            .I(N__20456));
    LocalMux I__4881 (
            .O(N__20456),
            .I(N__20452));
    CEMux I__4880 (
            .O(N__20455),
            .I(N__20449));
    Span4Mux_v I__4879 (
            .O(N__20452),
            .I(N__20444));
    LocalMux I__4878 (
            .O(N__20449),
            .I(N__20444));
    Span4Mux_v I__4877 (
            .O(N__20444),
            .I(N__20441));
    Odrv4 I__4876 (
            .O(N__20441),
            .I(\this_vram.mem_WE_2 ));
    SRMux I__4875 (
            .O(N__20438),
            .I(N__20431));
    SRMux I__4874 (
            .O(N__20437),
            .I(N__20428));
    SRMux I__4873 (
            .O(N__20436),
            .I(N__20424));
    SRMux I__4872 (
            .O(N__20435),
            .I(N__20421));
    SRMux I__4871 (
            .O(N__20434),
            .I(N__20416));
    LocalMux I__4870 (
            .O(N__20431),
            .I(N__20409));
    LocalMux I__4869 (
            .O(N__20428),
            .I(N__20409));
    SRMux I__4868 (
            .O(N__20427),
            .I(N__20406));
    LocalMux I__4867 (
            .O(N__20424),
            .I(N__20401));
    LocalMux I__4866 (
            .O(N__20421),
            .I(N__20401));
    SRMux I__4865 (
            .O(N__20420),
            .I(N__20398));
    SRMux I__4864 (
            .O(N__20419),
            .I(N__20395));
    LocalMux I__4863 (
            .O(N__20416),
            .I(N__20389));
    SRMux I__4862 (
            .O(N__20415),
            .I(N__20386));
    SRMux I__4861 (
            .O(N__20414),
            .I(N__20383));
    Span4Mux_s3_v I__4860 (
            .O(N__20409),
            .I(N__20376));
    LocalMux I__4859 (
            .O(N__20406),
            .I(N__20376));
    Span4Mux_s3_v I__4858 (
            .O(N__20401),
            .I(N__20369));
    LocalMux I__4857 (
            .O(N__20398),
            .I(N__20369));
    LocalMux I__4856 (
            .O(N__20395),
            .I(N__20369));
    SRMux I__4855 (
            .O(N__20394),
            .I(N__20366));
    SRMux I__4854 (
            .O(N__20393),
            .I(N__20363));
    IoInMux I__4853 (
            .O(N__20392),
            .I(N__20357));
    Span4Mux_h I__4852 (
            .O(N__20389),
            .I(N__20351));
    LocalMux I__4851 (
            .O(N__20386),
            .I(N__20351));
    LocalMux I__4850 (
            .O(N__20383),
            .I(N__20348));
    SRMux I__4849 (
            .O(N__20382),
            .I(N__20345));
    SRMux I__4848 (
            .O(N__20381),
            .I(N__20340));
    Span4Mux_v I__4847 (
            .O(N__20376),
            .I(N__20331));
    Span4Mux_v I__4846 (
            .O(N__20369),
            .I(N__20331));
    LocalMux I__4845 (
            .O(N__20366),
            .I(N__20331));
    LocalMux I__4844 (
            .O(N__20363),
            .I(N__20331));
    SRMux I__4843 (
            .O(N__20362),
            .I(N__20328));
    SRMux I__4842 (
            .O(N__20361),
            .I(N__20325));
    InMux I__4841 (
            .O(N__20360),
            .I(N__20319));
    LocalMux I__4840 (
            .O(N__20357),
            .I(N__20313));
    CascadeMux I__4839 (
            .O(N__20356),
            .I(N__20309));
    Span4Mux_v I__4838 (
            .O(N__20351),
            .I(N__20298));
    Span4Mux_h I__4837 (
            .O(N__20348),
            .I(N__20298));
    LocalMux I__4836 (
            .O(N__20345),
            .I(N__20298));
    SRMux I__4835 (
            .O(N__20344),
            .I(N__20295));
    SRMux I__4834 (
            .O(N__20343),
            .I(N__20291));
    LocalMux I__4833 (
            .O(N__20340),
            .I(N__20288));
    Span4Mux_v I__4832 (
            .O(N__20331),
            .I(N__20281));
    LocalMux I__4831 (
            .O(N__20328),
            .I(N__20281));
    LocalMux I__4830 (
            .O(N__20325),
            .I(N__20281));
    SRMux I__4829 (
            .O(N__20324),
            .I(N__20278));
    SRMux I__4828 (
            .O(N__20323),
            .I(N__20275));
    SRMux I__4827 (
            .O(N__20322),
            .I(N__20272));
    LocalMux I__4826 (
            .O(N__20319),
            .I(N__20268));
    CascadeMux I__4825 (
            .O(N__20318),
            .I(N__20264));
    CascadeMux I__4824 (
            .O(N__20317),
            .I(N__20260));
    CascadeMux I__4823 (
            .O(N__20316),
            .I(N__20256));
    IoSpan4Mux I__4822 (
            .O(N__20313),
            .I(N__20252));
    InMux I__4821 (
            .O(N__20312),
            .I(N__20247));
    InMux I__4820 (
            .O(N__20309),
            .I(N__20247));
    SRMux I__4819 (
            .O(N__20308),
            .I(N__20244));
    SRMux I__4818 (
            .O(N__20307),
            .I(N__20241));
    SRMux I__4817 (
            .O(N__20306),
            .I(N__20238));
    SRMux I__4816 (
            .O(N__20305),
            .I(N__20235));
    Span4Mux_v I__4815 (
            .O(N__20298),
            .I(N__20229));
    LocalMux I__4814 (
            .O(N__20295),
            .I(N__20229));
    SRMux I__4813 (
            .O(N__20294),
            .I(N__20226));
    LocalMux I__4812 (
            .O(N__20291),
            .I(N__20223));
    Span4Mux_h I__4811 (
            .O(N__20288),
            .I(N__20214));
    Span4Mux_v I__4810 (
            .O(N__20281),
            .I(N__20214));
    LocalMux I__4809 (
            .O(N__20278),
            .I(N__20214));
    LocalMux I__4808 (
            .O(N__20275),
            .I(N__20214));
    LocalMux I__4807 (
            .O(N__20272),
            .I(N__20211));
    SRMux I__4806 (
            .O(N__20271),
            .I(N__20208));
    Span4Mux_h I__4805 (
            .O(N__20268),
            .I(N__20204));
    InMux I__4804 (
            .O(N__20267),
            .I(N__20189));
    InMux I__4803 (
            .O(N__20264),
            .I(N__20189));
    InMux I__4802 (
            .O(N__20263),
            .I(N__20189));
    InMux I__4801 (
            .O(N__20260),
            .I(N__20189));
    InMux I__4800 (
            .O(N__20259),
            .I(N__20189));
    InMux I__4799 (
            .O(N__20256),
            .I(N__20189));
    InMux I__4798 (
            .O(N__20255),
            .I(N__20189));
    Span4Mux_s2_h I__4797 (
            .O(N__20252),
            .I(N__20185));
    LocalMux I__4796 (
            .O(N__20247),
            .I(N__20182));
    LocalMux I__4795 (
            .O(N__20244),
            .I(N__20175));
    LocalMux I__4794 (
            .O(N__20241),
            .I(N__20175));
    LocalMux I__4793 (
            .O(N__20238),
            .I(N__20170));
    LocalMux I__4792 (
            .O(N__20235),
            .I(N__20170));
    SRMux I__4791 (
            .O(N__20234),
            .I(N__20167));
    Span4Mux_v I__4790 (
            .O(N__20229),
            .I(N__20162));
    LocalMux I__4789 (
            .O(N__20226),
            .I(N__20162));
    Span4Mux_h I__4788 (
            .O(N__20223),
            .I(N__20153));
    Span4Mux_v I__4787 (
            .O(N__20214),
            .I(N__20153));
    Span4Mux_v I__4786 (
            .O(N__20211),
            .I(N__20153));
    LocalMux I__4785 (
            .O(N__20208),
            .I(N__20153));
    SRMux I__4784 (
            .O(N__20207),
            .I(N__20150));
    Span4Mux_h I__4783 (
            .O(N__20204),
            .I(N__20144));
    LocalMux I__4782 (
            .O(N__20189),
            .I(N__20144));
    SRMux I__4781 (
            .O(N__20188),
            .I(N__20141));
    Span4Mux_h I__4780 (
            .O(N__20185),
            .I(N__20136));
    Span4Mux_v I__4779 (
            .O(N__20182),
            .I(N__20136));
    CascadeMux I__4778 (
            .O(N__20181),
            .I(N__20132));
    SRMux I__4777 (
            .O(N__20180),
            .I(N__20128));
    Span4Mux_v I__4776 (
            .O(N__20175),
            .I(N__20115));
    Span4Mux_v I__4775 (
            .O(N__20170),
            .I(N__20115));
    LocalMux I__4774 (
            .O(N__20167),
            .I(N__20115));
    Span4Mux_v I__4773 (
            .O(N__20162),
            .I(N__20115));
    Span4Mux_v I__4772 (
            .O(N__20153),
            .I(N__20115));
    LocalMux I__4771 (
            .O(N__20150),
            .I(N__20115));
    SRMux I__4770 (
            .O(N__20149),
            .I(N__20112));
    Span4Mux_v I__4769 (
            .O(N__20144),
            .I(N__20109));
    LocalMux I__4768 (
            .O(N__20141),
            .I(N__20106));
    Sp12to4 I__4767 (
            .O(N__20136),
            .I(N__20103));
    InMux I__4766 (
            .O(N__20135),
            .I(N__20096));
    InMux I__4765 (
            .O(N__20132),
            .I(N__20096));
    InMux I__4764 (
            .O(N__20131),
            .I(N__20096));
    LocalMux I__4763 (
            .O(N__20128),
            .I(N__20093));
    Span4Mux_v I__4762 (
            .O(N__20115),
            .I(N__20088));
    LocalMux I__4761 (
            .O(N__20112),
            .I(N__20088));
    Span4Mux_h I__4760 (
            .O(N__20109),
            .I(N__20083));
    Span4Mux_h I__4759 (
            .O(N__20106),
            .I(N__20083));
    Span12Mux_h I__4758 (
            .O(N__20103),
            .I(N__20078));
    LocalMux I__4757 (
            .O(N__20096),
            .I(N__20078));
    Span4Mux_h I__4756 (
            .O(N__20093),
            .I(N__20075));
    Sp12to4 I__4755 (
            .O(N__20088),
            .I(N__20072));
    Span4Mux_h I__4754 (
            .O(N__20083),
            .I(N__20069));
    Odrv12 I__4753 (
            .O(N__20078),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4752 (
            .O(N__20075),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4751 (
            .O(N__20072),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4750 (
            .O(N__20069),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__4749 (
            .O(N__20060),
            .I(N__20056));
    InMux I__4748 (
            .O(N__20059),
            .I(N__20044));
    InMux I__4747 (
            .O(N__20056),
            .I(N__20041));
    CascadeMux I__4746 (
            .O(N__20055),
            .I(N__20036));
    CascadeMux I__4745 (
            .O(N__20054),
            .I(N__20033));
    CascadeMux I__4744 (
            .O(N__20053),
            .I(N__20030));
    CascadeMux I__4743 (
            .O(N__20052),
            .I(N__20027));
    CascadeMux I__4742 (
            .O(N__20051),
            .I(N__20024));
    CascadeMux I__4741 (
            .O(N__20050),
            .I(N__20020));
    CascadeMux I__4740 (
            .O(N__20049),
            .I(N__20016));
    CascadeMux I__4739 (
            .O(N__20048),
            .I(N__20012));
    CascadeMux I__4738 (
            .O(N__20047),
            .I(N__20008));
    LocalMux I__4737 (
            .O(N__20044),
            .I(N__20003));
    LocalMux I__4736 (
            .O(N__20041),
            .I(N__20003));
    InMux I__4735 (
            .O(N__20040),
            .I(N__20000));
    CascadeMux I__4734 (
            .O(N__20039),
            .I(N__19997));
    InMux I__4733 (
            .O(N__20036),
            .I(N__19990));
    InMux I__4732 (
            .O(N__20033),
            .I(N__19990));
    InMux I__4731 (
            .O(N__20030),
            .I(N__19983));
    InMux I__4730 (
            .O(N__20027),
            .I(N__19983));
    InMux I__4729 (
            .O(N__20024),
            .I(N__19983));
    InMux I__4728 (
            .O(N__20023),
            .I(N__19966));
    InMux I__4727 (
            .O(N__20020),
            .I(N__19966));
    InMux I__4726 (
            .O(N__20019),
            .I(N__19966));
    InMux I__4725 (
            .O(N__20016),
            .I(N__19966));
    InMux I__4724 (
            .O(N__20015),
            .I(N__19966));
    InMux I__4723 (
            .O(N__20012),
            .I(N__19966));
    InMux I__4722 (
            .O(N__20011),
            .I(N__19966));
    InMux I__4721 (
            .O(N__20008),
            .I(N__19966));
    Span4Mux_s2_h I__4720 (
            .O(N__20003),
            .I(N__19962));
    LocalMux I__4719 (
            .O(N__20000),
            .I(N__19959));
    InMux I__4718 (
            .O(N__19997),
            .I(N__19956));
    InMux I__4717 (
            .O(N__19996),
            .I(N__19951));
    InMux I__4716 (
            .O(N__19995),
            .I(N__19951));
    LocalMux I__4715 (
            .O(N__19990),
            .I(N__19944));
    LocalMux I__4714 (
            .O(N__19983),
            .I(N__19944));
    LocalMux I__4713 (
            .O(N__19966),
            .I(N__19944));
    InMux I__4712 (
            .O(N__19965),
            .I(N__19940));
    Span4Mux_h I__4711 (
            .O(N__19962),
            .I(N__19937));
    Span4Mux_v I__4710 (
            .O(N__19959),
            .I(N__19932));
    LocalMux I__4709 (
            .O(N__19956),
            .I(N__19932));
    LocalMux I__4708 (
            .O(N__19951),
            .I(N__19927));
    Span4Mux_v I__4707 (
            .O(N__19944),
            .I(N__19927));
    InMux I__4706 (
            .O(N__19943),
            .I(N__19924));
    LocalMux I__4705 (
            .O(N__19940),
            .I(N__19921));
    Span4Mux_h I__4704 (
            .O(N__19937),
            .I(N__19918));
    Span4Mux_h I__4703 (
            .O(N__19932),
            .I(N__19911));
    Span4Mux_h I__4702 (
            .O(N__19927),
            .I(N__19911));
    LocalMux I__4701 (
            .O(N__19924),
            .I(N__19911));
    Span4Mux_h I__4700 (
            .O(N__19921),
            .I(N__19908));
    Odrv4 I__4699 (
            .O(N__19918),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__4698 (
            .O(N__19911),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__4697 (
            .O(N__19908),
            .I(M_this_state_qZ0Z_3));
    IoInMux I__4696 (
            .O(N__19901),
            .I(N__19898));
    LocalMux I__4695 (
            .O(N__19898),
            .I(N__19895));
    Span4Mux_s1_v I__4694 (
            .O(N__19895),
            .I(N__19892));
    Sp12to4 I__4693 (
            .O(N__19892),
            .I(N__19889));
    Span12Mux_h I__4692 (
            .O(N__19889),
            .I(N__19885));
    InMux I__4691 (
            .O(N__19888),
            .I(N__19882));
    Odrv12 I__4690 (
            .O(N__19885),
            .I(M_this_external_address_qZ0Z_0));
    LocalMux I__4689 (
            .O(N__19882),
            .I(M_this_external_address_qZ0Z_0));
    IoInMux I__4688 (
            .O(N__19877),
            .I(N__19874));
    LocalMux I__4687 (
            .O(N__19874),
            .I(N__19871));
    IoSpan4Mux I__4686 (
            .O(N__19871),
            .I(N__19868));
    Sp12to4 I__4685 (
            .O(N__19868),
            .I(N__19864));
    InMux I__4684 (
            .O(N__19867),
            .I(N__19861));
    Odrv12 I__4683 (
            .O(N__19864),
            .I(M_this_external_address_qZ0Z_1));
    LocalMux I__4682 (
            .O(N__19861),
            .I(M_this_external_address_qZ0Z_1));
    InMux I__4681 (
            .O(N__19856),
            .I(un1_M_this_external_address_q_cry_0));
    IoInMux I__4680 (
            .O(N__19853),
            .I(N__19850));
    LocalMux I__4679 (
            .O(N__19850),
            .I(N__19847));
    IoSpan4Mux I__4678 (
            .O(N__19847),
            .I(N__19844));
    IoSpan4Mux I__4677 (
            .O(N__19844),
            .I(N__19841));
    Span4Mux_s2_v I__4676 (
            .O(N__19841),
            .I(N__19838));
    Span4Mux_v I__4675 (
            .O(N__19838),
            .I(N__19834));
    InMux I__4674 (
            .O(N__19837),
            .I(N__19831));
    Odrv4 I__4673 (
            .O(N__19834),
            .I(M_this_external_address_qZ0Z_2));
    LocalMux I__4672 (
            .O(N__19831),
            .I(M_this_external_address_qZ0Z_2));
    InMux I__4671 (
            .O(N__19826),
            .I(un1_M_this_external_address_q_cry_1));
    IoInMux I__4670 (
            .O(N__19823),
            .I(N__19820));
    LocalMux I__4669 (
            .O(N__19820),
            .I(N__19817));
    Span4Mux_s2_h I__4668 (
            .O(N__19817),
            .I(N__19814));
    Span4Mux_v I__4667 (
            .O(N__19814),
            .I(N__19810));
    InMux I__4666 (
            .O(N__19813),
            .I(N__19807));
    Odrv4 I__4665 (
            .O(N__19810),
            .I(M_this_external_address_qZ0Z_3));
    LocalMux I__4664 (
            .O(N__19807),
            .I(M_this_external_address_qZ0Z_3));
    InMux I__4663 (
            .O(N__19802),
            .I(un1_M_this_external_address_q_cry_2));
    IoInMux I__4662 (
            .O(N__19799),
            .I(N__19796));
    LocalMux I__4661 (
            .O(N__19796),
            .I(N__19792));
    InMux I__4660 (
            .O(N__19795),
            .I(N__19789));
    Odrv4 I__4659 (
            .O(N__19792),
            .I(M_this_external_address_qZ0Z_4));
    LocalMux I__4658 (
            .O(N__19789),
            .I(M_this_external_address_qZ0Z_4));
    InMux I__4657 (
            .O(N__19784),
            .I(N__19781));
    LocalMux I__4656 (
            .O(N__19781),
            .I(N__19778));
    Odrv4 I__4655 (
            .O(N__19778),
            .I(\this_vram.mem_out_bus5_1 ));
    InMux I__4654 (
            .O(N__19775),
            .I(N__19772));
    LocalMux I__4653 (
            .O(N__19772),
            .I(N__19769));
    Odrv4 I__4652 (
            .O(N__19769),
            .I(\this_vram.mem_mem_1_0_RNISSK11Z0Z_0 ));
    InMux I__4651 (
            .O(N__19766),
            .I(N__19763));
    LocalMux I__4650 (
            .O(N__19763),
            .I(N__19760));
    Span4Mux_v I__4649 (
            .O(N__19760),
            .I(N__19757));
    Odrv4 I__4648 (
            .O(N__19757),
            .I(\this_vram.mem_out_bus5_2 ));
    InMux I__4647 (
            .O(N__19754),
            .I(N__19751));
    LocalMux I__4646 (
            .O(N__19751),
            .I(N__19748));
    Span4Mux_v I__4645 (
            .O(N__19748),
            .I(N__19745));
    Span4Mux_v I__4644 (
            .O(N__19745),
            .I(N__19742));
    Odrv4 I__4643 (
            .O(N__19742),
            .I(\this_vram.mem_out_bus1_2 ));
    InMux I__4642 (
            .O(N__19739),
            .I(N__19736));
    LocalMux I__4641 (
            .O(N__19736),
            .I(\this_vram.mem_mem_1_1_RNIUSKZ0Z11 ));
    InMux I__4640 (
            .O(N__19733),
            .I(N__19730));
    LocalMux I__4639 (
            .O(N__19730),
            .I(N__19727));
    Span4Mux_v I__4638 (
            .O(N__19727),
            .I(N__19724));
    Sp12to4 I__4637 (
            .O(N__19724),
            .I(N__19721));
    Odrv12 I__4636 (
            .O(N__19721),
            .I(\this_vram.mem_out_bus7_2 ));
    InMux I__4635 (
            .O(N__19718),
            .I(N__19715));
    LocalMux I__4634 (
            .O(N__19715),
            .I(N__19712));
    Span4Mux_h I__4633 (
            .O(N__19712),
            .I(N__19709));
    Odrv4 I__4632 (
            .O(N__19709),
            .I(\this_vram.mem_out_bus3_2 ));
    InMux I__4631 (
            .O(N__19706),
            .I(N__19703));
    LocalMux I__4630 (
            .O(N__19703),
            .I(\this_vram.mem_mem_3_1_RNI25PZ0Z11 ));
    InMux I__4629 (
            .O(N__19700),
            .I(N__19697));
    LocalMux I__4628 (
            .O(N__19697),
            .I(N__19694));
    Span4Mux_v I__4627 (
            .O(N__19694),
            .I(N__19691));
    Span4Mux_v I__4626 (
            .O(N__19691),
            .I(N__19688));
    Odrv4 I__4625 (
            .O(N__19688),
            .I(\this_vram.mem_out_bus7_0 ));
    InMux I__4624 (
            .O(N__19685),
            .I(N__19682));
    LocalMux I__4623 (
            .O(N__19682),
            .I(N__19679));
    Span4Mux_v I__4622 (
            .O(N__19679),
            .I(N__19676));
    Span4Mux_v I__4621 (
            .O(N__19676),
            .I(N__19673));
    Odrv4 I__4620 (
            .O(N__19673),
            .I(\this_vram.mem_out_bus3_0 ));
    InMux I__4619 (
            .O(N__19670),
            .I(N__19667));
    LocalMux I__4618 (
            .O(N__19667),
            .I(\this_vram.mem_mem_3_0_RNI05PZ0Z11 ));
    InMux I__4617 (
            .O(N__19664),
            .I(N__19661));
    LocalMux I__4616 (
            .O(N__19661),
            .I(N__19658));
    Span4Mux_v I__4615 (
            .O(N__19658),
            .I(N__19655));
    Odrv4 I__4614 (
            .O(N__19655),
            .I(\this_vram.mem_out_bus2_2 ));
    CascadeMux I__4613 (
            .O(N__19652),
            .I(N__19649));
    InMux I__4612 (
            .O(N__19649),
            .I(N__19646));
    LocalMux I__4611 (
            .O(N__19646),
            .I(N__19643));
    Sp12to4 I__4610 (
            .O(N__19643),
            .I(N__19640));
    Odrv12 I__4609 (
            .O(N__19640),
            .I(\this_vram.mem_out_bus6_2 ));
    CascadeMux I__4608 (
            .O(N__19637),
            .I(N__19634));
    InMux I__4607 (
            .O(N__19634),
            .I(N__19631));
    LocalMux I__4606 (
            .O(N__19631),
            .I(\this_vram.mem_mem_2_1_RNI01NZ0Z11 ));
    InMux I__4605 (
            .O(N__19628),
            .I(N__19612));
    InMux I__4604 (
            .O(N__19627),
            .I(N__19601));
    InMux I__4603 (
            .O(N__19626),
            .I(N__19601));
    InMux I__4602 (
            .O(N__19625),
            .I(N__19601));
    InMux I__4601 (
            .O(N__19624),
            .I(N__19601));
    InMux I__4600 (
            .O(N__19623),
            .I(N__19601));
    InMux I__4599 (
            .O(N__19622),
            .I(N__19598));
    InMux I__4598 (
            .O(N__19621),
            .I(N__19593));
    InMux I__4597 (
            .O(N__19620),
            .I(N__19593));
    InMux I__4596 (
            .O(N__19619),
            .I(N__19590));
    InMux I__4595 (
            .O(N__19618),
            .I(N__19587));
    InMux I__4594 (
            .O(N__19617),
            .I(N__19580));
    InMux I__4593 (
            .O(N__19616),
            .I(N__19580));
    InMux I__4592 (
            .O(N__19615),
            .I(N__19580));
    LocalMux I__4591 (
            .O(N__19612),
            .I(N__19571));
    LocalMux I__4590 (
            .O(N__19601),
            .I(N__19571));
    LocalMux I__4589 (
            .O(N__19598),
            .I(N__19571));
    LocalMux I__4588 (
            .O(N__19593),
            .I(N__19571));
    LocalMux I__4587 (
            .O(N__19590),
            .I(N__19564));
    LocalMux I__4586 (
            .O(N__19587),
            .I(N__19564));
    LocalMux I__4585 (
            .O(N__19580),
            .I(N__19564));
    Span4Mux_v I__4584 (
            .O(N__19571),
            .I(N__19561));
    Span4Mux_h I__4583 (
            .O(N__19564),
            .I(N__19558));
    Odrv4 I__4582 (
            .O(N__19561),
            .I(\this_vram.mem_radregZ0Z_13 ));
    Odrv4 I__4581 (
            .O(N__19558),
            .I(\this_vram.mem_radregZ0Z_13 ));
    InMux I__4580 (
            .O(N__19553),
            .I(N__19550));
    LocalMux I__4579 (
            .O(N__19550),
            .I(N__19547));
    Odrv4 I__4578 (
            .O(N__19547),
            .I(\this_vram.mem_out_bus5_0 ));
    InMux I__4577 (
            .O(N__19544),
            .I(N__19541));
    LocalMux I__4576 (
            .O(N__19541),
            .I(N__19538));
    Span4Mux_v I__4575 (
            .O(N__19538),
            .I(N__19535));
    Span4Mux_v I__4574 (
            .O(N__19535),
            .I(N__19532));
    Span4Mux_v I__4573 (
            .O(N__19532),
            .I(N__19529));
    Odrv4 I__4572 (
            .O(N__19529),
            .I(\this_vram.mem_out_bus1_0 ));
    InMux I__4571 (
            .O(N__19526),
            .I(N__19523));
    LocalMux I__4570 (
            .O(N__19523),
            .I(\this_vram.mem_mem_1_0_RNISSKZ0Z11 ));
    CascadeMux I__4569 (
            .O(N__19520),
            .I(N__19516));
    CascadeMux I__4568 (
            .O(N__19519),
            .I(N__19513));
    InMux I__4567 (
            .O(N__19516),
            .I(N__19510));
    InMux I__4566 (
            .O(N__19513),
            .I(N__19507));
    LocalMux I__4565 (
            .O(N__19510),
            .I(N__19503));
    LocalMux I__4564 (
            .O(N__19507),
            .I(N__19500));
    InMux I__4563 (
            .O(N__19506),
            .I(N__19497));
    Span4Mux_v I__4562 (
            .O(N__19503),
            .I(N__19494));
    Span4Mux_h I__4561 (
            .O(N__19500),
            .I(N__19491));
    LocalMux I__4560 (
            .O(N__19497),
            .I(N__19488));
    Sp12to4 I__4559 (
            .O(N__19494),
            .I(N__19485));
    Span4Mux_h I__4558 (
            .O(N__19491),
            .I(N__19480));
    Span4Mux_v I__4557 (
            .O(N__19488),
            .I(N__19480));
    Span12Mux_h I__4556 (
            .O(N__19485),
            .I(N__19477));
    Span4Mux_h I__4555 (
            .O(N__19480),
            .I(N__19474));
    Span12Mux_v I__4554 (
            .O(N__19477),
            .I(N__19471));
    Sp12to4 I__4553 (
            .O(N__19474),
            .I(N__19468));
    Odrv12 I__4552 (
            .O(N__19471),
            .I(port_data_c_3));
    Odrv12 I__4551 (
            .O(N__19468),
            .I(port_data_c_3));
    CascadeMux I__4550 (
            .O(N__19463),
            .I(N__19460));
    InMux I__4549 (
            .O(N__19460),
            .I(N__19457));
    LocalMux I__4548 (
            .O(N__19457),
            .I(N__19454));
    Span4Mux_h I__4547 (
            .O(N__19454),
            .I(N__19451));
    Sp12to4 I__4546 (
            .O(N__19451),
            .I(N__19448));
    Span12Mux_v I__4545 (
            .O(N__19448),
            .I(N__19445));
    Odrv12 I__4544 (
            .O(N__19445),
            .I(port_data_c_7));
    InMux I__4543 (
            .O(N__19442),
            .I(N__19439));
    LocalMux I__4542 (
            .O(N__19439),
            .I(N__19435));
    InMux I__4541 (
            .O(N__19438),
            .I(N__19432));
    Span4Mux_v I__4540 (
            .O(N__19435),
            .I(N__19425));
    LocalMux I__4539 (
            .O(N__19432),
            .I(N__19425));
    InMux I__4538 (
            .O(N__19431),
            .I(N__19422));
    InMux I__4537 (
            .O(N__19430),
            .I(N__19418));
    Span4Mux_v I__4536 (
            .O(N__19425),
            .I(N__19412));
    LocalMux I__4535 (
            .O(N__19422),
            .I(N__19412));
    InMux I__4534 (
            .O(N__19421),
            .I(N__19409));
    LocalMux I__4533 (
            .O(N__19418),
            .I(N__19406));
    InMux I__4532 (
            .O(N__19417),
            .I(N__19403));
    Span4Mux_v I__4531 (
            .O(N__19412),
            .I(N__19397));
    LocalMux I__4530 (
            .O(N__19409),
            .I(N__19397));
    Span4Mux_v I__4529 (
            .O(N__19406),
            .I(N__19392));
    LocalMux I__4528 (
            .O(N__19403),
            .I(N__19392));
    InMux I__4527 (
            .O(N__19402),
            .I(N__19389));
    Span4Mux_v I__4526 (
            .O(N__19397),
            .I(N__19385));
    Span4Mux_v I__4525 (
            .O(N__19392),
            .I(N__19380));
    LocalMux I__4524 (
            .O(N__19389),
            .I(N__19380));
    InMux I__4523 (
            .O(N__19388),
            .I(N__19377));
    Odrv4 I__4522 (
            .O(N__19385),
            .I(M_this_vram_write_data_0_i_3));
    Odrv4 I__4521 (
            .O(N__19380),
            .I(M_this_vram_write_data_0_i_3));
    LocalMux I__4520 (
            .O(N__19377),
            .I(M_this_vram_write_data_0_i_3));
    CEMux I__4519 (
            .O(N__19370),
            .I(N__19366));
    CEMux I__4518 (
            .O(N__19369),
            .I(N__19363));
    LocalMux I__4517 (
            .O(N__19366),
            .I(N__19360));
    LocalMux I__4516 (
            .O(N__19363),
            .I(N__19357));
    Span4Mux_v I__4515 (
            .O(N__19360),
            .I(N__19354));
    Span4Mux_h I__4514 (
            .O(N__19357),
            .I(N__19351));
    Span4Mux_h I__4513 (
            .O(N__19354),
            .I(N__19348));
    Span4Mux_h I__4512 (
            .O(N__19351),
            .I(N__19345));
    Odrv4 I__4511 (
            .O(N__19348),
            .I(\this_vram.mem_WE_4 ));
    Odrv4 I__4510 (
            .O(N__19345),
            .I(\this_vram.mem_WE_4 ));
    InMux I__4509 (
            .O(N__19340),
            .I(N__19337));
    LocalMux I__4508 (
            .O(N__19337),
            .I(N__19334));
    Odrv4 I__4507 (
            .O(N__19334),
            .I(\this_vram.mem_mem_0_1_RNISOIZ0Z11 ));
    InMux I__4506 (
            .O(N__19331),
            .I(N__19328));
    LocalMux I__4505 (
            .O(N__19328),
            .I(N__19325));
    Span4Mux_v I__4504 (
            .O(N__19325),
            .I(N__19322));
    Odrv4 I__4503 (
            .O(N__19322),
            .I(\this_vram.mem_out_bus5_3 ));
    InMux I__4502 (
            .O(N__19319),
            .I(N__19316));
    LocalMux I__4501 (
            .O(N__19316),
            .I(N__19313));
    Span4Mux_v I__4500 (
            .O(N__19313),
            .I(N__19310));
    Span4Mux_v I__4499 (
            .O(N__19310),
            .I(N__19307));
    Odrv4 I__4498 (
            .O(N__19307),
            .I(\this_vram.mem_out_bus1_3 ));
    InMux I__4497 (
            .O(N__19304),
            .I(N__19301));
    LocalMux I__4496 (
            .O(N__19301),
            .I(N__19298));
    Odrv4 I__4495 (
            .O(N__19298),
            .I(\this_vram.mem_out_bus3_3 ));
    InMux I__4494 (
            .O(N__19295),
            .I(N__19292));
    LocalMux I__4493 (
            .O(N__19292),
            .I(N__19289));
    Sp12to4 I__4492 (
            .O(N__19289),
            .I(N__19286));
    Span12Mux_v I__4491 (
            .O(N__19286),
            .I(N__19283));
    Odrv12 I__4490 (
            .O(N__19283),
            .I(\this_vram.mem_out_bus7_3 ));
    CascadeMux I__4489 (
            .O(N__19280),
            .I(\this_vram.mem_DOUT_6_i_m2_ns_1_3_cascade_ ));
    InMux I__4488 (
            .O(N__19277),
            .I(N__19274));
    LocalMux I__4487 (
            .O(N__19274),
            .I(\this_vram.mem_N_102 ));
    InMux I__4486 (
            .O(N__19271),
            .I(N__19268));
    LocalMux I__4485 (
            .O(N__19268),
            .I(N__19265));
    Span4Mux_h I__4484 (
            .O(N__19265),
            .I(N__19262));
    Odrv4 I__4483 (
            .O(N__19262),
            .I(\this_vram.mem_out_bus4_3 ));
    InMux I__4482 (
            .O(N__19259),
            .I(N__19256));
    LocalMux I__4481 (
            .O(N__19256),
            .I(N__19253));
    Sp12to4 I__4480 (
            .O(N__19253),
            .I(N__19250));
    Span12Mux_v I__4479 (
            .O(N__19250),
            .I(N__19247));
    Odrv12 I__4478 (
            .O(N__19247),
            .I(\this_vram.mem_out_bus0_3 ));
    InMux I__4477 (
            .O(N__19244),
            .I(N__19241));
    LocalMux I__4476 (
            .O(N__19241),
            .I(N__19238));
    Span4Mux_v I__4475 (
            .O(N__19238),
            .I(N__19235));
    Span4Mux_v I__4474 (
            .O(N__19235),
            .I(N__19232));
    Odrv4 I__4473 (
            .O(N__19232),
            .I(\this_vram.mem_out_bus6_3 ));
    InMux I__4472 (
            .O(N__19229),
            .I(N__19226));
    LocalMux I__4471 (
            .O(N__19226),
            .I(N__19223));
    Span4Mux_v I__4470 (
            .O(N__19223),
            .I(N__19220));
    Odrv4 I__4469 (
            .O(N__19220),
            .I(\this_vram.mem_out_bus2_3 ));
    CascadeMux I__4468 (
            .O(N__19217),
            .I(\this_vram.mem_DOUT_3_i_m2_ns_1_3_cascade_ ));
    CascadeMux I__4467 (
            .O(N__19214),
            .I(N__19206));
    CascadeMux I__4466 (
            .O(N__19213),
            .I(N__19203));
    InMux I__4465 (
            .O(N__19212),
            .I(N__19200));
    InMux I__4464 (
            .O(N__19211),
            .I(N__19196));
    InMux I__4463 (
            .O(N__19210),
            .I(N__19187));
    InMux I__4462 (
            .O(N__19209),
            .I(N__19187));
    InMux I__4461 (
            .O(N__19206),
            .I(N__19187));
    InMux I__4460 (
            .O(N__19203),
            .I(N__19187));
    LocalMux I__4459 (
            .O(N__19200),
            .I(N__19184));
    InMux I__4458 (
            .O(N__19199),
            .I(N__19181));
    LocalMux I__4457 (
            .O(N__19196),
            .I(N__19178));
    LocalMux I__4456 (
            .O(N__19187),
            .I(N__19175));
    Span4Mux_h I__4455 (
            .O(N__19184),
            .I(N__19172));
    LocalMux I__4454 (
            .O(N__19181),
            .I(N__19165));
    Span4Mux_v I__4453 (
            .O(N__19178),
            .I(N__19165));
    Span4Mux_v I__4452 (
            .O(N__19175),
            .I(N__19165));
    Odrv4 I__4451 (
            .O(N__19172),
            .I(\this_vram.mem_radregZ0Z_12 ));
    Odrv4 I__4450 (
            .O(N__19165),
            .I(\this_vram.mem_radregZ0Z_12 ));
    InMux I__4449 (
            .O(N__19160),
            .I(N__19157));
    LocalMux I__4448 (
            .O(N__19157),
            .I(\this_vram.mem_N_105 ));
    InMux I__4447 (
            .O(N__19154),
            .I(N__19151));
    LocalMux I__4446 (
            .O(N__19151),
            .I(N__19148));
    Sp12to4 I__4445 (
            .O(N__19148),
            .I(N__19145));
    Span12Mux_v I__4444 (
            .O(N__19145),
            .I(N__19142));
    Odrv12 I__4443 (
            .O(N__19142),
            .I(\this_vram.mem_out_bus0_0 ));
    InMux I__4442 (
            .O(N__19139),
            .I(N__19136));
    LocalMux I__4441 (
            .O(N__19136),
            .I(\this_vram.mem_out_bus4_0 ));
    CascadeMux I__4440 (
            .O(N__19133),
            .I(N__19130));
    InMux I__4439 (
            .O(N__19130),
            .I(N__19127));
    LocalMux I__4438 (
            .O(N__19127),
            .I(\this_vram.mem_mem_0_0_RNIQOIZ0Z11 ));
    InMux I__4437 (
            .O(N__19124),
            .I(N__19121));
    LocalMux I__4436 (
            .O(N__19121),
            .I(N__19118));
    Sp12to4 I__4435 (
            .O(N__19118),
            .I(N__19115));
    Odrv12 I__4434 (
            .O(N__19115),
            .I(\this_vram.mem_out_bus6_0 ));
    InMux I__4433 (
            .O(N__19112),
            .I(N__19109));
    LocalMux I__4432 (
            .O(N__19109),
            .I(N__19106));
    Span4Mux_v I__4431 (
            .O(N__19106),
            .I(N__19103));
    Span4Mux_v I__4430 (
            .O(N__19103),
            .I(N__19100));
    Odrv4 I__4429 (
            .O(N__19100),
            .I(\this_vram.mem_out_bus2_0 ));
    InMux I__4428 (
            .O(N__19097),
            .I(N__19094));
    LocalMux I__4427 (
            .O(N__19094),
            .I(\this_vram.mem_mem_2_0_RNIU0NZ0Z11 ));
    CEMux I__4426 (
            .O(N__19091),
            .I(N__19088));
    LocalMux I__4425 (
            .O(N__19088),
            .I(N__19084));
    CEMux I__4424 (
            .O(N__19087),
            .I(N__19081));
    Span4Mux_h I__4423 (
            .O(N__19084),
            .I(N__19078));
    LocalMux I__4422 (
            .O(N__19081),
            .I(N__19075));
    Odrv4 I__4421 (
            .O(N__19078),
            .I(\this_vram.mem_WE_6 ));
    Odrv12 I__4420 (
            .O(N__19075),
            .I(\this_vram.mem_WE_6 ));
    InMux I__4419 (
            .O(N__19070),
            .I(N__19067));
    LocalMux I__4418 (
            .O(N__19067),
            .I(N__19064));
    Sp12to4 I__4417 (
            .O(N__19064),
            .I(N__19061));
    Span12Mux_v I__4416 (
            .O(N__19061),
            .I(N__19058));
    Odrv12 I__4415 (
            .O(N__19058),
            .I(\this_vram.mem_out_bus1_1 ));
    InMux I__4414 (
            .O(N__19055),
            .I(N__19048));
    InMux I__4413 (
            .O(N__19054),
            .I(N__19048));
    CascadeMux I__4412 (
            .O(N__19053),
            .I(N__19045));
    LocalMux I__4411 (
            .O(N__19048),
            .I(N__19042));
    InMux I__4410 (
            .O(N__19045),
            .I(N__19039));
    Span4Mux_h I__4409 (
            .O(N__19042),
            .I(N__19036));
    LocalMux I__4408 (
            .O(N__19039),
            .I(M_this_state_qZ0Z_7));
    Odrv4 I__4407 (
            .O(N__19036),
            .I(M_this_state_qZ0Z_7));
    InMux I__4406 (
            .O(N__19031),
            .I(N__19027));
    InMux I__4405 (
            .O(N__19030),
            .I(N__19024));
    LocalMux I__4404 (
            .O(N__19027),
            .I(N__19020));
    LocalMux I__4403 (
            .O(N__19024),
            .I(N__19016));
    InMux I__4402 (
            .O(N__19023),
            .I(N__19011));
    Span4Mux_v I__4401 (
            .O(N__19020),
            .I(N__19008));
    InMux I__4400 (
            .O(N__19019),
            .I(N__19005));
    Span4Mux_v I__4399 (
            .O(N__19016),
            .I(N__19002));
    InMux I__4398 (
            .O(N__19015),
            .I(N__18999));
    InMux I__4397 (
            .O(N__19014),
            .I(N__18996));
    LocalMux I__4396 (
            .O(N__19011),
            .I(N__18989));
    Sp12to4 I__4395 (
            .O(N__19008),
            .I(N__18989));
    LocalMux I__4394 (
            .O(N__19005),
            .I(N__18989));
    Odrv4 I__4393 (
            .O(N__19002),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__4392 (
            .O(N__18999),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__4391 (
            .O(N__18996),
            .I(M_this_state_qZ0Z_2));
    Odrv12 I__4390 (
            .O(N__18989),
            .I(M_this_state_qZ0Z_2));
    CascadeMux I__4389 (
            .O(N__18980),
            .I(N__18976));
    InMux I__4388 (
            .O(N__18979),
            .I(N__18972));
    InMux I__4387 (
            .O(N__18976),
            .I(N__18969));
    InMux I__4386 (
            .O(N__18975),
            .I(N__18966));
    LocalMux I__4385 (
            .O(N__18972),
            .I(N__18963));
    LocalMux I__4384 (
            .O(N__18969),
            .I(N__18960));
    LocalMux I__4383 (
            .O(N__18966),
            .I(N__18957));
    Span4Mux_v I__4382 (
            .O(N__18963),
            .I(N__18952));
    Span4Mux_v I__4381 (
            .O(N__18960),
            .I(N__18952));
    Span4Mux_v I__4380 (
            .O(N__18957),
            .I(N__18949));
    Sp12to4 I__4379 (
            .O(N__18952),
            .I(N__18944));
    Sp12to4 I__4378 (
            .O(N__18949),
            .I(N__18944));
    Span12Mux_h I__4377 (
            .O(N__18944),
            .I(N__18941));
    Odrv12 I__4376 (
            .O(N__18941),
            .I(port_data_c_0));
    InMux I__4375 (
            .O(N__18938),
            .I(N__18934));
    CascadeMux I__4374 (
            .O(N__18937),
            .I(N__18930));
    LocalMux I__4373 (
            .O(N__18934),
            .I(N__18927));
    InMux I__4372 (
            .O(N__18933),
            .I(N__18924));
    InMux I__4371 (
            .O(N__18930),
            .I(N__18921));
    Span4Mux_v I__4370 (
            .O(N__18927),
            .I(N__18918));
    LocalMux I__4369 (
            .O(N__18924),
            .I(N__18915));
    LocalMux I__4368 (
            .O(N__18921),
            .I(N__18912));
    Span4Mux_h I__4367 (
            .O(N__18918),
            .I(N__18907));
    Span4Mux_v I__4366 (
            .O(N__18915),
            .I(N__18907));
    Span12Mux_v I__4365 (
            .O(N__18912),
            .I(N__18904));
    Span4Mux_v I__4364 (
            .O(N__18907),
            .I(N__18901));
    Span12Mux_h I__4363 (
            .O(N__18904),
            .I(N__18898));
    Sp12to4 I__4362 (
            .O(N__18901),
            .I(N__18895));
    Odrv12 I__4361 (
            .O(N__18898),
            .I(port_data_c_4));
    Odrv12 I__4360 (
            .O(N__18895),
            .I(port_data_c_4));
    CascadeMux I__4359 (
            .O(N__18890),
            .I(M_this_vram_write_data_0_sqmuxa_cascade_));
    InMux I__4358 (
            .O(N__18887),
            .I(N__18884));
    LocalMux I__4357 (
            .O(N__18884),
            .I(N__18880));
    InMux I__4356 (
            .O(N__18883),
            .I(N__18877));
    Span4Mux_h I__4355 (
            .O(N__18880),
            .I(N__18873));
    LocalMux I__4354 (
            .O(N__18877),
            .I(N__18870));
    InMux I__4353 (
            .O(N__18876),
            .I(N__18867));
    Span4Mux_v I__4352 (
            .O(N__18873),
            .I(N__18860));
    Span4Mux_h I__4351 (
            .O(N__18870),
            .I(N__18860));
    LocalMux I__4350 (
            .O(N__18867),
            .I(N__18857));
    InMux I__4349 (
            .O(N__18866),
            .I(N__18854));
    InMux I__4348 (
            .O(N__18865),
            .I(N__18850));
    Span4Mux_v I__4347 (
            .O(N__18860),
            .I(N__18844));
    Span4Mux_h I__4346 (
            .O(N__18857),
            .I(N__18844));
    LocalMux I__4345 (
            .O(N__18854),
            .I(N__18841));
    InMux I__4344 (
            .O(N__18853),
            .I(N__18838));
    LocalMux I__4343 (
            .O(N__18850),
            .I(N__18835));
    InMux I__4342 (
            .O(N__18849),
            .I(N__18832));
    Span4Mux_v I__4341 (
            .O(N__18844),
            .I(N__18826));
    Span4Mux_h I__4340 (
            .O(N__18841),
            .I(N__18826));
    LocalMux I__4339 (
            .O(N__18838),
            .I(N__18823));
    Span4Mux_v I__4338 (
            .O(N__18835),
            .I(N__18818));
    LocalMux I__4337 (
            .O(N__18832),
            .I(N__18818));
    InMux I__4336 (
            .O(N__18831),
            .I(N__18815));
    Span4Mux_v I__4335 (
            .O(N__18826),
            .I(N__18810));
    Span4Mux_h I__4334 (
            .O(N__18823),
            .I(N__18810));
    Span4Mux_v I__4333 (
            .O(N__18818),
            .I(N__18805));
    LocalMux I__4332 (
            .O(N__18815),
            .I(N__18805));
    Odrv4 I__4331 (
            .O(N__18810),
            .I(M_this_vram_write_data_0_i_0));
    Odrv4 I__4330 (
            .O(N__18805),
            .I(M_this_vram_write_data_0_i_0));
    InMux I__4329 (
            .O(N__18800),
            .I(N__18787));
    InMux I__4328 (
            .O(N__18799),
            .I(N__18784));
    InMux I__4327 (
            .O(N__18798),
            .I(N__18780));
    InMux I__4326 (
            .O(N__18797),
            .I(N__18777));
    InMux I__4325 (
            .O(N__18796),
            .I(N__18772));
    InMux I__4324 (
            .O(N__18795),
            .I(N__18772));
    InMux I__4323 (
            .O(N__18794),
            .I(N__18764));
    InMux I__4322 (
            .O(N__18793),
            .I(N__18764));
    InMux I__4321 (
            .O(N__18792),
            .I(N__18764));
    InMux I__4320 (
            .O(N__18791),
            .I(N__18756));
    InMux I__4319 (
            .O(N__18790),
            .I(N__18756));
    LocalMux I__4318 (
            .O(N__18787),
            .I(N__18751));
    LocalMux I__4317 (
            .O(N__18784),
            .I(N__18751));
    InMux I__4316 (
            .O(N__18783),
            .I(N__18748));
    LocalMux I__4315 (
            .O(N__18780),
            .I(N__18741));
    LocalMux I__4314 (
            .O(N__18777),
            .I(N__18741));
    LocalMux I__4313 (
            .O(N__18772),
            .I(N__18741));
    InMux I__4312 (
            .O(N__18771),
            .I(N__18733));
    LocalMux I__4311 (
            .O(N__18764),
            .I(N__18730));
    InMux I__4310 (
            .O(N__18763),
            .I(N__18725));
    InMux I__4309 (
            .O(N__18762),
            .I(N__18725));
    InMux I__4308 (
            .O(N__18761),
            .I(N__18722));
    LocalMux I__4307 (
            .O(N__18756),
            .I(N__18717));
    Span12Mux_h I__4306 (
            .O(N__18751),
            .I(N__18717));
    LocalMux I__4305 (
            .O(N__18748),
            .I(N__18712));
    Span4Mux_h I__4304 (
            .O(N__18741),
            .I(N__18712));
    InMux I__4303 (
            .O(N__18740),
            .I(N__18709));
    InMux I__4302 (
            .O(N__18739),
            .I(N__18700));
    InMux I__4301 (
            .O(N__18738),
            .I(N__18700));
    InMux I__4300 (
            .O(N__18737),
            .I(N__18700));
    InMux I__4299 (
            .O(N__18736),
            .I(N__18700));
    LocalMux I__4298 (
            .O(N__18733),
            .I(M_this_start_data_delay_out_0));
    Odrv4 I__4297 (
            .O(N__18730),
            .I(M_this_start_data_delay_out_0));
    LocalMux I__4296 (
            .O(N__18725),
            .I(M_this_start_data_delay_out_0));
    LocalMux I__4295 (
            .O(N__18722),
            .I(M_this_start_data_delay_out_0));
    Odrv12 I__4294 (
            .O(N__18717),
            .I(M_this_start_data_delay_out_0));
    Odrv4 I__4293 (
            .O(N__18712),
            .I(M_this_start_data_delay_out_0));
    LocalMux I__4292 (
            .O(N__18709),
            .I(M_this_start_data_delay_out_0));
    LocalMux I__4291 (
            .O(N__18700),
            .I(M_this_start_data_delay_out_0));
    InMux I__4290 (
            .O(N__18683),
            .I(N__18679));
    InMux I__4289 (
            .O(N__18682),
            .I(N__18676));
    LocalMux I__4288 (
            .O(N__18679),
            .I(N__18673));
    LocalMux I__4287 (
            .O(N__18676),
            .I(\this_start_data_delay.N_351_0 ));
    Odrv12 I__4286 (
            .O(N__18673),
            .I(\this_start_data_delay.N_351_0 ));
    CEMux I__4285 (
            .O(N__18668),
            .I(N__18665));
    LocalMux I__4284 (
            .O(N__18665),
            .I(N__18662));
    Span12Mux_s8_h I__4283 (
            .O(N__18662),
            .I(N__18658));
    CEMux I__4282 (
            .O(N__18661),
            .I(N__18655));
    Odrv12 I__4281 (
            .O(N__18658),
            .I(\this_vram.mem_WE_8 ));
    LocalMux I__4280 (
            .O(N__18655),
            .I(\this_vram.mem_WE_8 ));
    CEMux I__4279 (
            .O(N__18650),
            .I(N__18647));
    LocalMux I__4278 (
            .O(N__18647),
            .I(N__18643));
    CEMux I__4277 (
            .O(N__18646),
            .I(N__18640));
    Span4Mux_v I__4276 (
            .O(N__18643),
            .I(N__18637));
    LocalMux I__4275 (
            .O(N__18640),
            .I(N__18634));
    Span4Mux_v I__4274 (
            .O(N__18637),
            .I(N__18631));
    Span12Mux_s8_h I__4273 (
            .O(N__18634),
            .I(N__18628));
    Odrv4 I__4272 (
            .O(N__18631),
            .I(\this_vram.mem_WE_12 ));
    Odrv12 I__4271 (
            .O(N__18628),
            .I(\this_vram.mem_WE_12 ));
    CEMux I__4270 (
            .O(N__18623),
            .I(N__18619));
    CEMux I__4269 (
            .O(N__18622),
            .I(N__18616));
    LocalMux I__4268 (
            .O(N__18619),
            .I(N__18613));
    LocalMux I__4267 (
            .O(N__18616),
            .I(N__18610));
    Span4Mux_v I__4266 (
            .O(N__18613),
            .I(N__18605));
    Span4Mux_h I__4265 (
            .O(N__18610),
            .I(N__18605));
    Odrv4 I__4264 (
            .O(N__18605),
            .I(\this_vram.mem_WE_10 ));
    InMux I__4263 (
            .O(N__18602),
            .I(N__18599));
    LocalMux I__4262 (
            .O(N__18599),
            .I(N__18596));
    Span4Mux_h I__4261 (
            .O(N__18596),
            .I(N__18593));
    Odrv4 I__4260 (
            .O(N__18593),
            .I(\this_vram.mem_out_bus4_2 ));
    InMux I__4259 (
            .O(N__18590),
            .I(N__18587));
    LocalMux I__4258 (
            .O(N__18587),
            .I(N__18584));
    Sp12to4 I__4257 (
            .O(N__18584),
            .I(N__18581));
    Span12Mux_v I__4256 (
            .O(N__18581),
            .I(N__18578));
    Odrv12 I__4255 (
            .O(N__18578),
            .I(\this_vram.mem_out_bus0_2 ));
    CEMux I__4254 (
            .O(N__18575),
            .I(N__18571));
    CEMux I__4253 (
            .O(N__18574),
            .I(N__18568));
    LocalMux I__4252 (
            .O(N__18571),
            .I(N__18565));
    LocalMux I__4251 (
            .O(N__18568),
            .I(N__18562));
    Span4Mux_h I__4250 (
            .O(N__18565),
            .I(N__18559));
    Span4Mux_h I__4249 (
            .O(N__18562),
            .I(N__18556));
    Span4Mux_v I__4248 (
            .O(N__18559),
            .I(N__18553));
    Sp12to4 I__4247 (
            .O(N__18556),
            .I(N__18550));
    Span4Mux_v I__4246 (
            .O(N__18553),
            .I(N__18547));
    Odrv12 I__4245 (
            .O(N__18550),
            .I(\this_vram.mem_WE_14 ));
    Odrv4 I__4244 (
            .O(N__18547),
            .I(\this_vram.mem_WE_14 ));
    InMux I__4243 (
            .O(N__18542),
            .I(N__18539));
    LocalMux I__4242 (
            .O(N__18539),
            .I(N__18536));
    Span4Mux_h I__4241 (
            .O(N__18536),
            .I(N__18533));
    Span4Mux_v I__4240 (
            .O(N__18533),
            .I(N__18530));
    Odrv4 I__4239 (
            .O(N__18530),
            .I(\this_vram.mem_out_bus6_1 ));
    InMux I__4238 (
            .O(N__18527),
            .I(N__18524));
    LocalMux I__4237 (
            .O(N__18524),
            .I(N__18521));
    Span4Mux_v I__4236 (
            .O(N__18521),
            .I(N__18518));
    Span4Mux_v I__4235 (
            .O(N__18518),
            .I(N__18515));
    Odrv4 I__4234 (
            .O(N__18515),
            .I(\this_vram.mem_out_bus2_1 ));
    InMux I__4233 (
            .O(N__18512),
            .I(N__18509));
    LocalMux I__4232 (
            .O(N__18509),
            .I(\this_vram.mem_mem_2_0_RNIU0N11Z0Z_0 ));
    InMux I__4231 (
            .O(N__18506),
            .I(N__18503));
    LocalMux I__4230 (
            .O(N__18503),
            .I(N__18500));
    Span4Mux_v I__4229 (
            .O(N__18500),
            .I(N__18497));
    Span4Mux_v I__4228 (
            .O(N__18497),
            .I(N__18494));
    Span4Mux_v I__4227 (
            .O(N__18494),
            .I(N__18491));
    Odrv4 I__4226 (
            .O(N__18491),
            .I(\this_vram.mem_out_bus7_1 ));
    InMux I__4225 (
            .O(N__18488),
            .I(N__18485));
    LocalMux I__4224 (
            .O(N__18485),
            .I(N__18482));
    Span4Mux_v I__4223 (
            .O(N__18482),
            .I(N__18479));
    Span4Mux_v I__4222 (
            .O(N__18479),
            .I(N__18476));
    Odrv4 I__4221 (
            .O(N__18476),
            .I(\this_vram.mem_out_bus3_1 ));
    InMux I__4220 (
            .O(N__18473),
            .I(N__18470));
    LocalMux I__4219 (
            .O(N__18470),
            .I(\this_vram.mem_mem_3_0_RNI05P11Z0Z_0 ));
    CascadeMux I__4218 (
            .O(N__18467),
            .I(N__18463));
    InMux I__4217 (
            .O(N__18466),
            .I(N__18456));
    InMux I__4216 (
            .O(N__18463),
            .I(N__18451));
    InMux I__4215 (
            .O(N__18462),
            .I(N__18451));
    InMux I__4214 (
            .O(N__18461),
            .I(N__18444));
    InMux I__4213 (
            .O(N__18460),
            .I(N__18444));
    InMux I__4212 (
            .O(N__18459),
            .I(N__18444));
    LocalMux I__4211 (
            .O(N__18456),
            .I(N__18441));
    LocalMux I__4210 (
            .O(N__18451),
            .I(N__18436));
    LocalMux I__4209 (
            .O(N__18444),
            .I(N__18436));
    Span4Mux_v I__4208 (
            .O(N__18441),
            .I(N__18431));
    Span4Mux_v I__4207 (
            .O(N__18436),
            .I(N__18431));
    Sp12to4 I__4206 (
            .O(N__18431),
            .I(N__18428));
    Span12Mux_h I__4205 (
            .O(N__18428),
            .I(N__18425));
    Odrv12 I__4204 (
            .O(N__18425),
            .I(M_this_vram_read_data_3));
    CascadeMux I__4203 (
            .O(N__18422),
            .I(\this_vram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ));
    CascadeMux I__4202 (
            .O(N__18419),
            .I(N__18414));
    CascadeMux I__4201 (
            .O(N__18418),
            .I(N__18409));
    CascadeMux I__4200 (
            .O(N__18417),
            .I(N__18406));
    InMux I__4199 (
            .O(N__18414),
            .I(N__18403));
    CascadeMux I__4198 (
            .O(N__18413),
            .I(N__18400));
    InMux I__4197 (
            .O(N__18412),
            .I(N__18393));
    InMux I__4196 (
            .O(N__18409),
            .I(N__18393));
    InMux I__4195 (
            .O(N__18406),
            .I(N__18393));
    LocalMux I__4194 (
            .O(N__18403),
            .I(N__18390));
    InMux I__4193 (
            .O(N__18400),
            .I(N__18387));
    LocalMux I__4192 (
            .O(N__18393),
            .I(N__18384));
    Span12Mux_s10_h I__4191 (
            .O(N__18390),
            .I(N__18381));
    LocalMux I__4190 (
            .O(N__18387),
            .I(N__18376));
    Span12Mux_s5_h I__4189 (
            .O(N__18384),
            .I(N__18376));
    Span12Mux_h I__4188 (
            .O(N__18381),
            .I(N__18373));
    Span12Mux_h I__4187 (
            .O(N__18376),
            .I(N__18370));
    Odrv12 I__4186 (
            .O(N__18373),
            .I(M_this_vram_read_data_2));
    Odrv12 I__4185 (
            .O(N__18370),
            .I(M_this_vram_read_data_2));
    CascadeMux I__4184 (
            .O(N__18365),
            .I(N__18360));
    CascadeMux I__4183 (
            .O(N__18364),
            .I(N__18356));
    InMux I__4182 (
            .O(N__18363),
            .I(N__18352));
    InMux I__4181 (
            .O(N__18360),
            .I(N__18347));
    InMux I__4180 (
            .O(N__18359),
            .I(N__18340));
    InMux I__4179 (
            .O(N__18356),
            .I(N__18340));
    InMux I__4178 (
            .O(N__18355),
            .I(N__18340));
    LocalMux I__4177 (
            .O(N__18352),
            .I(N__18337));
    InMux I__4176 (
            .O(N__18351),
            .I(N__18332));
    InMux I__4175 (
            .O(N__18350),
            .I(N__18332));
    LocalMux I__4174 (
            .O(N__18347),
            .I(\this_vram.mem_radregZ0Z_11 ));
    LocalMux I__4173 (
            .O(N__18340),
            .I(\this_vram.mem_radregZ0Z_11 ));
    Odrv4 I__4172 (
            .O(N__18337),
            .I(\this_vram.mem_radregZ0Z_11 ));
    LocalMux I__4171 (
            .O(N__18332),
            .I(\this_vram.mem_radregZ0Z_11 ));
    InMux I__4170 (
            .O(N__18323),
            .I(N__18320));
    LocalMux I__4169 (
            .O(N__18320),
            .I(\this_vram.mem_DOUT_7_i_m2_ns_1_0 ));
    InMux I__4168 (
            .O(N__18317),
            .I(N__18314));
    LocalMux I__4167 (
            .O(N__18314),
            .I(N__18311));
    Span4Mux_v I__4166 (
            .O(N__18311),
            .I(N__18303));
    InMux I__4165 (
            .O(N__18310),
            .I(N__18296));
    InMux I__4164 (
            .O(N__18309),
            .I(N__18296));
    InMux I__4163 (
            .O(N__18308),
            .I(N__18296));
    InMux I__4162 (
            .O(N__18307),
            .I(N__18291));
    InMux I__4161 (
            .O(N__18306),
            .I(N__18291));
    Sp12to4 I__4160 (
            .O(N__18303),
            .I(N__18284));
    LocalMux I__4159 (
            .O(N__18296),
            .I(N__18284));
    LocalMux I__4158 (
            .O(N__18291),
            .I(N__18284));
    Span12Mux_s11_h I__4157 (
            .O(N__18284),
            .I(N__18281));
    Odrv12 I__4156 (
            .O(N__18281),
            .I(M_this_vram_read_data_0));
    CascadeMux I__4155 (
            .O(N__18278),
            .I(N__18275));
    InMux I__4154 (
            .O(N__18275),
            .I(N__18271));
    InMux I__4153 (
            .O(N__18274),
            .I(N__18267));
    LocalMux I__4152 (
            .O(N__18271),
            .I(N__18264));
    CascadeMux I__4151 (
            .O(N__18270),
            .I(N__18261));
    LocalMux I__4150 (
            .O(N__18267),
            .I(N__18258));
    Span4Mux_v I__4149 (
            .O(N__18264),
            .I(N__18255));
    InMux I__4148 (
            .O(N__18261),
            .I(N__18252));
    Span4Mux_v I__4147 (
            .O(N__18258),
            .I(N__18249));
    Span4Mux_h I__4146 (
            .O(N__18255),
            .I(N__18244));
    LocalMux I__4145 (
            .O(N__18252),
            .I(N__18244));
    Span4Mux_v I__4144 (
            .O(N__18249),
            .I(N__18241));
    Span4Mux_v I__4143 (
            .O(N__18244),
            .I(N__18238));
    Sp12to4 I__4142 (
            .O(N__18241),
            .I(N__18233));
    Sp12to4 I__4141 (
            .O(N__18238),
            .I(N__18233));
    Span12Mux_h I__4140 (
            .O(N__18233),
            .I(N__18230));
    Odrv12 I__4139 (
            .O(N__18230),
            .I(port_data_c_1));
    CascadeMux I__4138 (
            .O(N__18227),
            .I(N__18223));
    CascadeMux I__4137 (
            .O(N__18226),
            .I(N__18220));
    InMux I__4136 (
            .O(N__18223),
            .I(N__18216));
    InMux I__4135 (
            .O(N__18220),
            .I(N__18213));
    CascadeMux I__4134 (
            .O(N__18219),
            .I(N__18210));
    LocalMux I__4133 (
            .O(N__18216),
            .I(N__18205));
    LocalMux I__4132 (
            .O(N__18213),
            .I(N__18205));
    InMux I__4131 (
            .O(N__18210),
            .I(N__18202));
    Span4Mux_v I__4130 (
            .O(N__18205),
            .I(N__18199));
    LocalMux I__4129 (
            .O(N__18202),
            .I(N__18196));
    Span4Mux_h I__4128 (
            .O(N__18199),
            .I(N__18191));
    Span4Mux_v I__4127 (
            .O(N__18196),
            .I(N__18191));
    Sp12to4 I__4126 (
            .O(N__18191),
            .I(N__18188));
    Odrv12 I__4125 (
            .O(N__18188),
            .I(port_data_c_5));
    InMux I__4124 (
            .O(N__18185),
            .I(N__18181));
    InMux I__4123 (
            .O(N__18184),
            .I(N__18177));
    LocalMux I__4122 (
            .O(N__18181),
            .I(N__18172));
    InMux I__4121 (
            .O(N__18180),
            .I(N__18168));
    LocalMux I__4120 (
            .O(N__18177),
            .I(N__18165));
    InMux I__4119 (
            .O(N__18176),
            .I(N__18161));
    InMux I__4118 (
            .O(N__18175),
            .I(N__18158));
    Span4Mux_h I__4117 (
            .O(N__18172),
            .I(N__18155));
    InMux I__4116 (
            .O(N__18171),
            .I(N__18152));
    LocalMux I__4115 (
            .O(N__18168),
            .I(N__18149));
    Span4Mux_h I__4114 (
            .O(N__18165),
            .I(N__18146));
    InMux I__4113 (
            .O(N__18164),
            .I(N__18143));
    LocalMux I__4112 (
            .O(N__18161),
            .I(N__18140));
    LocalMux I__4111 (
            .O(N__18158),
            .I(N__18137));
    Span4Mux_v I__4110 (
            .O(N__18155),
            .I(N__18132));
    LocalMux I__4109 (
            .O(N__18152),
            .I(N__18132));
    Span12Mux_s9_h I__4108 (
            .O(N__18149),
            .I(N__18128));
    Sp12to4 I__4107 (
            .O(N__18146),
            .I(N__18125));
    LocalMux I__4106 (
            .O(N__18143),
            .I(N__18122));
    Span4Mux_v I__4105 (
            .O(N__18140),
            .I(N__18119));
    Span4Mux_h I__4104 (
            .O(N__18137),
            .I(N__18116));
    Span4Mux_h I__4103 (
            .O(N__18132),
            .I(N__18113));
    InMux I__4102 (
            .O(N__18131),
            .I(N__18110));
    Span12Mux_v I__4101 (
            .O(N__18128),
            .I(N__18107));
    Span12Mux_s8_v I__4100 (
            .O(N__18125),
            .I(N__18102));
    Span12Mux_s9_h I__4099 (
            .O(N__18122),
            .I(N__18102));
    Span4Mux_v I__4098 (
            .O(N__18119),
            .I(N__18093));
    Span4Mux_v I__4097 (
            .O(N__18116),
            .I(N__18093));
    Span4Mux_v I__4096 (
            .O(N__18113),
            .I(N__18093));
    LocalMux I__4095 (
            .O(N__18110),
            .I(N__18093));
    Odrv12 I__4094 (
            .O(N__18107),
            .I(M_this_vram_write_data_0_i_1));
    Odrv12 I__4093 (
            .O(N__18102),
            .I(M_this_vram_write_data_0_i_1));
    Odrv4 I__4092 (
            .O(N__18093),
            .I(M_this_vram_write_data_0_i_1));
    CascadeMux I__4091 (
            .O(N__18086),
            .I(N__18077));
    CascadeMux I__4090 (
            .O(N__18085),
            .I(N__18074));
    CascadeMux I__4089 (
            .O(N__18084),
            .I(N__18070));
    CascadeMux I__4088 (
            .O(N__18083),
            .I(N__18066));
    CascadeMux I__4087 (
            .O(N__18082),
            .I(N__18063));
    CascadeMux I__4086 (
            .O(N__18081),
            .I(N__18060));
    CascadeMux I__4085 (
            .O(N__18080),
            .I(N__18057));
    InMux I__4084 (
            .O(N__18077),
            .I(N__18052));
    InMux I__4083 (
            .O(N__18074),
            .I(N__18052));
    CascadeMux I__4082 (
            .O(N__18073),
            .I(N__18047));
    InMux I__4081 (
            .O(N__18070),
            .I(N__18042));
    InMux I__4080 (
            .O(N__18069),
            .I(N__18035));
    InMux I__4079 (
            .O(N__18066),
            .I(N__18035));
    InMux I__4078 (
            .O(N__18063),
            .I(N__18035));
    InMux I__4077 (
            .O(N__18060),
            .I(N__18032));
    InMux I__4076 (
            .O(N__18057),
            .I(N__18029));
    LocalMux I__4075 (
            .O(N__18052),
            .I(N__18026));
    CascadeMux I__4074 (
            .O(N__18051),
            .I(N__18023));
    InMux I__4073 (
            .O(N__18050),
            .I(N__18014));
    InMux I__4072 (
            .O(N__18047),
            .I(N__18014));
    InMux I__4071 (
            .O(N__18046),
            .I(N__18014));
    InMux I__4070 (
            .O(N__18045),
            .I(N__18014));
    LocalMux I__4069 (
            .O(N__18042),
            .I(N__18008));
    LocalMux I__4068 (
            .O(N__18035),
            .I(N__18008));
    LocalMux I__4067 (
            .O(N__18032),
            .I(N__18001));
    LocalMux I__4066 (
            .O(N__18029),
            .I(N__18001));
    Span4Mux_h I__4065 (
            .O(N__18026),
            .I(N__18001));
    InMux I__4064 (
            .O(N__18023),
            .I(N__17998));
    LocalMux I__4063 (
            .O(N__18014),
            .I(N__17995));
    InMux I__4062 (
            .O(N__18013),
            .I(N__17992));
    Span4Mux_h I__4061 (
            .O(N__18008),
            .I(N__17989));
    Span4Mux_v I__4060 (
            .O(N__18001),
            .I(N__17986));
    LocalMux I__4059 (
            .O(N__17998),
            .I(N__17981));
    Span12Mux_h I__4058 (
            .O(N__17995),
            .I(N__17981));
    LocalMux I__4057 (
            .O(N__17992),
            .I(M_this_internal_address_q_3_sm0_0));
    Odrv4 I__4056 (
            .O(N__17989),
            .I(M_this_internal_address_q_3_sm0_0));
    Odrv4 I__4055 (
            .O(N__17986),
            .I(M_this_internal_address_q_3_sm0_0));
    Odrv12 I__4054 (
            .O(N__17981),
            .I(M_this_internal_address_q_3_sm0_0));
    InMux I__4053 (
            .O(N__17972),
            .I(N__17969));
    LocalMux I__4052 (
            .O(N__17969),
            .I(N__17966));
    Odrv4 I__4051 (
            .O(N__17966),
            .I(\this_vram.mem_out_bus4_1 ));
    InMux I__4050 (
            .O(N__17963),
            .I(N__17960));
    LocalMux I__4049 (
            .O(N__17960),
            .I(N__17957));
    Span12Mux_h I__4048 (
            .O(N__17957),
            .I(N__17954));
    Span12Mux_v I__4047 (
            .O(N__17954),
            .I(N__17951));
    Odrv12 I__4046 (
            .O(N__17951),
            .I(\this_vram.mem_out_bus0_1 ));
    CascadeMux I__4045 (
            .O(N__17948),
            .I(\this_vram.mem_mem_0_0_RNIQOI11Z0Z_0_cascade_ ));
    InMux I__4044 (
            .O(N__17945),
            .I(N__17942));
    LocalMux I__4043 (
            .O(N__17942),
            .I(N__17939));
    Odrv12 I__4042 (
            .O(N__17939),
            .I(M_this_vga_signals_address_11));
    InMux I__4041 (
            .O(N__17936),
            .I(N__17933));
    LocalMux I__4040 (
            .O(N__17933),
            .I(\this_vram.mem_DOUT_7_i_m2_ns_1_1 ));
    CascadeMux I__4039 (
            .O(N__17930),
            .I(N__17927));
    InMux I__4038 (
            .O(N__17927),
            .I(N__17915));
    InMux I__4037 (
            .O(N__17926),
            .I(N__17915));
    InMux I__4036 (
            .O(N__17925),
            .I(N__17915));
    InMux I__4035 (
            .O(N__17924),
            .I(N__17912));
    InMux I__4034 (
            .O(N__17923),
            .I(N__17907));
    InMux I__4033 (
            .O(N__17922),
            .I(N__17907));
    LocalMux I__4032 (
            .O(N__17915),
            .I(N__17904));
    LocalMux I__4031 (
            .O(N__17912),
            .I(N__17899));
    LocalMux I__4030 (
            .O(N__17907),
            .I(N__17899));
    Span4Mux_v I__4029 (
            .O(N__17904),
            .I(N__17896));
    Span4Mux_v I__4028 (
            .O(N__17899),
            .I(N__17893));
    Span4Mux_h I__4027 (
            .O(N__17896),
            .I(N__17890));
    Sp12to4 I__4026 (
            .O(N__17893),
            .I(N__17885));
    Sp12to4 I__4025 (
            .O(N__17890),
            .I(N__17885));
    Span12Mux_h I__4024 (
            .O(N__17885),
            .I(N__17882));
    Odrv12 I__4023 (
            .O(N__17882),
            .I(M_this_vram_read_data_1));
    CascadeMux I__4022 (
            .O(N__17879),
            .I(N__17876));
    CascadeBuf I__4021 (
            .O(N__17876),
            .I(N__17873));
    CascadeMux I__4020 (
            .O(N__17873),
            .I(N__17870));
    CascadeBuf I__4019 (
            .O(N__17870),
            .I(N__17867));
    CascadeMux I__4018 (
            .O(N__17867),
            .I(N__17864));
    CascadeBuf I__4017 (
            .O(N__17864),
            .I(N__17861));
    CascadeMux I__4016 (
            .O(N__17861),
            .I(N__17858));
    CascadeBuf I__4015 (
            .O(N__17858),
            .I(N__17855));
    CascadeMux I__4014 (
            .O(N__17855),
            .I(N__17852));
    CascadeBuf I__4013 (
            .O(N__17852),
            .I(N__17849));
    CascadeMux I__4012 (
            .O(N__17849),
            .I(N__17846));
    CascadeBuf I__4011 (
            .O(N__17846),
            .I(N__17843));
    CascadeMux I__4010 (
            .O(N__17843),
            .I(N__17840));
    CascadeBuf I__4009 (
            .O(N__17840),
            .I(N__17837));
    CascadeMux I__4008 (
            .O(N__17837),
            .I(N__17834));
    CascadeBuf I__4007 (
            .O(N__17834),
            .I(N__17831));
    CascadeMux I__4006 (
            .O(N__17831),
            .I(N__17828));
    CascadeBuf I__4005 (
            .O(N__17828),
            .I(N__17825));
    CascadeMux I__4004 (
            .O(N__17825),
            .I(N__17822));
    CascadeBuf I__4003 (
            .O(N__17822),
            .I(N__17819));
    CascadeMux I__4002 (
            .O(N__17819),
            .I(N__17816));
    CascadeBuf I__4001 (
            .O(N__17816),
            .I(N__17813));
    CascadeMux I__4000 (
            .O(N__17813),
            .I(N__17810));
    CascadeBuf I__3999 (
            .O(N__17810),
            .I(N__17807));
    CascadeMux I__3998 (
            .O(N__17807),
            .I(N__17804));
    CascadeBuf I__3997 (
            .O(N__17804),
            .I(N__17801));
    CascadeMux I__3996 (
            .O(N__17801),
            .I(N__17798));
    CascadeBuf I__3995 (
            .O(N__17798),
            .I(N__17795));
    CascadeMux I__3994 (
            .O(N__17795),
            .I(N__17792));
    CascadeBuf I__3993 (
            .O(N__17792),
            .I(N__17789));
    CascadeMux I__3992 (
            .O(N__17789),
            .I(N__17786));
    InMux I__3991 (
            .O(N__17786),
            .I(N__17783));
    LocalMux I__3990 (
            .O(N__17783),
            .I(N__17780));
    Span4Mux_v I__3989 (
            .O(N__17780),
            .I(N__17777));
    Span4Mux_h I__3988 (
            .O(N__17777),
            .I(N__17772));
    InMux I__3987 (
            .O(N__17776),
            .I(N__17769));
    InMux I__3986 (
            .O(N__17775),
            .I(N__17766));
    Span4Mux_v I__3985 (
            .O(N__17772),
            .I(N__17763));
    LocalMux I__3984 (
            .O(N__17769),
            .I(M_this_internal_address_qZ0Z_6));
    LocalMux I__3983 (
            .O(N__17766),
            .I(M_this_internal_address_qZ0Z_6));
    Odrv4 I__3982 (
            .O(N__17763),
            .I(M_this_internal_address_qZ0Z_6));
    InMux I__3981 (
            .O(N__17756),
            .I(N__17753));
    LocalMux I__3980 (
            .O(N__17753),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_6 ));
    InMux I__3979 (
            .O(N__17750),
            .I(N__17742));
    InMux I__3978 (
            .O(N__17749),
            .I(N__17738));
    InMux I__3977 (
            .O(N__17748),
            .I(N__17727));
    InMux I__3976 (
            .O(N__17747),
            .I(N__17727));
    InMux I__3975 (
            .O(N__17746),
            .I(N__17727));
    CascadeMux I__3974 (
            .O(N__17745),
            .I(N__17723));
    LocalMux I__3973 (
            .O(N__17742),
            .I(N__17716));
    InMux I__3972 (
            .O(N__17741),
            .I(N__17713));
    LocalMux I__3971 (
            .O(N__17738),
            .I(N__17710));
    InMux I__3970 (
            .O(N__17737),
            .I(N__17707));
    InMux I__3969 (
            .O(N__17736),
            .I(N__17700));
    InMux I__3968 (
            .O(N__17735),
            .I(N__17700));
    InMux I__3967 (
            .O(N__17734),
            .I(N__17700));
    LocalMux I__3966 (
            .O(N__17727),
            .I(N__17697));
    InMux I__3965 (
            .O(N__17726),
            .I(N__17694));
    InMux I__3964 (
            .O(N__17723),
            .I(N__17691));
    InMux I__3963 (
            .O(N__17722),
            .I(N__17688));
    InMux I__3962 (
            .O(N__17721),
            .I(N__17685));
    InMux I__3961 (
            .O(N__17720),
            .I(N__17680));
    InMux I__3960 (
            .O(N__17719),
            .I(N__17680));
    Span4Mux_v I__3959 (
            .O(N__17716),
            .I(N__17677));
    LocalMux I__3958 (
            .O(N__17713),
            .I(N__17674));
    Span4Mux_h I__3957 (
            .O(N__17710),
            .I(N__17671));
    LocalMux I__3956 (
            .O(N__17707),
            .I(N__17666));
    LocalMux I__3955 (
            .O(N__17700),
            .I(N__17666));
    Span4Mux_v I__3954 (
            .O(N__17697),
            .I(N__17661));
    LocalMux I__3953 (
            .O(N__17694),
            .I(N__17661));
    LocalMux I__3952 (
            .O(N__17691),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__3951 (
            .O(N__17688),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__3950 (
            .O(N__17685),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__3949 (
            .O(N__17680),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__3948 (
            .O(N__17677),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__3947 (
            .O(N__17674),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__3946 (
            .O(N__17671),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__3945 (
            .O(N__17666),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__3944 (
            .O(N__17661),
            .I(M_this_state_qZ0Z_5));
    CascadeMux I__3943 (
            .O(N__17642),
            .I(N__17639));
    CascadeBuf I__3942 (
            .O(N__17639),
            .I(N__17636));
    CascadeMux I__3941 (
            .O(N__17636),
            .I(N__17633));
    CascadeBuf I__3940 (
            .O(N__17633),
            .I(N__17630));
    CascadeMux I__3939 (
            .O(N__17630),
            .I(N__17627));
    CascadeBuf I__3938 (
            .O(N__17627),
            .I(N__17624));
    CascadeMux I__3937 (
            .O(N__17624),
            .I(N__17621));
    CascadeBuf I__3936 (
            .O(N__17621),
            .I(N__17618));
    CascadeMux I__3935 (
            .O(N__17618),
            .I(N__17615));
    CascadeBuf I__3934 (
            .O(N__17615),
            .I(N__17612));
    CascadeMux I__3933 (
            .O(N__17612),
            .I(N__17609));
    CascadeBuf I__3932 (
            .O(N__17609),
            .I(N__17606));
    CascadeMux I__3931 (
            .O(N__17606),
            .I(N__17603));
    CascadeBuf I__3930 (
            .O(N__17603),
            .I(N__17600));
    CascadeMux I__3929 (
            .O(N__17600),
            .I(N__17597));
    CascadeBuf I__3928 (
            .O(N__17597),
            .I(N__17594));
    CascadeMux I__3927 (
            .O(N__17594),
            .I(N__17591));
    CascadeBuf I__3926 (
            .O(N__17591),
            .I(N__17588));
    CascadeMux I__3925 (
            .O(N__17588),
            .I(N__17585));
    CascadeBuf I__3924 (
            .O(N__17585),
            .I(N__17582));
    CascadeMux I__3923 (
            .O(N__17582),
            .I(N__17579));
    CascadeBuf I__3922 (
            .O(N__17579),
            .I(N__17576));
    CascadeMux I__3921 (
            .O(N__17576),
            .I(N__17573));
    CascadeBuf I__3920 (
            .O(N__17573),
            .I(N__17570));
    CascadeMux I__3919 (
            .O(N__17570),
            .I(N__17567));
    CascadeBuf I__3918 (
            .O(N__17567),
            .I(N__17564));
    CascadeMux I__3917 (
            .O(N__17564),
            .I(N__17561));
    CascadeBuf I__3916 (
            .O(N__17561),
            .I(N__17558));
    CascadeMux I__3915 (
            .O(N__17558),
            .I(N__17555));
    CascadeBuf I__3914 (
            .O(N__17555),
            .I(N__17552));
    CascadeMux I__3913 (
            .O(N__17552),
            .I(N__17549));
    InMux I__3912 (
            .O(N__17549),
            .I(N__17546));
    LocalMux I__3911 (
            .O(N__17546),
            .I(N__17543));
    Span4Mux_s2_v I__3910 (
            .O(N__17543),
            .I(N__17540));
    Span4Mux_v I__3909 (
            .O(N__17540),
            .I(N__17535));
    InMux I__3908 (
            .O(N__17539),
            .I(N__17532));
    InMux I__3907 (
            .O(N__17538),
            .I(N__17529));
    Span4Mux_v I__3906 (
            .O(N__17535),
            .I(N__17526));
    LocalMux I__3905 (
            .O(N__17532),
            .I(M_this_internal_address_qZ0Z_8));
    LocalMux I__3904 (
            .O(N__17529),
            .I(M_this_internal_address_qZ0Z_8));
    Odrv4 I__3903 (
            .O(N__17526),
            .I(M_this_internal_address_qZ0Z_8));
    InMux I__3902 (
            .O(N__17519),
            .I(N__17516));
    LocalMux I__3901 (
            .O(N__17516),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_8 ));
    InMux I__3900 (
            .O(N__17513),
            .I(N__17510));
    LocalMux I__3899 (
            .O(N__17510),
            .I(N__17507));
    Span12Mux_h I__3898 (
            .O(N__17507),
            .I(N__17504));
    Odrv12 I__3897 (
            .O(N__17504),
            .I(port_address_in_3));
    InMux I__3896 (
            .O(N__17501),
            .I(N__17498));
    LocalMux I__3895 (
            .O(N__17498),
            .I(N__17495));
    Odrv12 I__3894 (
            .O(N__17495),
            .I(port_address_in_2));
    InMux I__3893 (
            .O(N__17492),
            .I(N__17480));
    InMux I__3892 (
            .O(N__17491),
            .I(N__17480));
    InMux I__3891 (
            .O(N__17490),
            .I(N__17480));
    InMux I__3890 (
            .O(N__17489),
            .I(N__17480));
    LocalMux I__3889 (
            .O(N__17480),
            .I(N__17477));
    Span4Mux_v I__3888 (
            .O(N__17477),
            .I(N__17474));
    Odrv4 I__3887 (
            .O(N__17474),
            .I(\this_start_data_delay.M_this_state_d27Z0Z_2 ));
    InMux I__3886 (
            .O(N__17471),
            .I(N__17468));
    LocalMux I__3885 (
            .O(N__17468),
            .I(N__17465));
    Span4Mux_h I__3884 (
            .O(N__17465),
            .I(N__17462));
    Odrv4 I__3883 (
            .O(N__17462),
            .I(un1_M_this_internal_address_q_cry_10_c_RNI6I0DZ0));
    InMux I__3882 (
            .O(N__17459),
            .I(un1_M_this_internal_address_q_cry_10));
    InMux I__3881 (
            .O(N__17456),
            .I(un1_M_this_internal_address_q_cry_11));
    InMux I__3880 (
            .O(N__17453),
            .I(un1_M_this_internal_address_q_cry_12));
    CascadeMux I__3879 (
            .O(N__17450),
            .I(N__17447));
    CascadeBuf I__3878 (
            .O(N__17447),
            .I(N__17444));
    CascadeMux I__3877 (
            .O(N__17444),
            .I(N__17441));
    CascadeBuf I__3876 (
            .O(N__17441),
            .I(N__17438));
    CascadeMux I__3875 (
            .O(N__17438),
            .I(N__17435));
    CascadeBuf I__3874 (
            .O(N__17435),
            .I(N__17432));
    CascadeMux I__3873 (
            .O(N__17432),
            .I(N__17429));
    CascadeBuf I__3872 (
            .O(N__17429),
            .I(N__17426));
    CascadeMux I__3871 (
            .O(N__17426),
            .I(N__17423));
    CascadeBuf I__3870 (
            .O(N__17423),
            .I(N__17420));
    CascadeMux I__3869 (
            .O(N__17420),
            .I(N__17417));
    CascadeBuf I__3868 (
            .O(N__17417),
            .I(N__17414));
    CascadeMux I__3867 (
            .O(N__17414),
            .I(N__17411));
    CascadeBuf I__3866 (
            .O(N__17411),
            .I(N__17408));
    CascadeMux I__3865 (
            .O(N__17408),
            .I(N__17405));
    CascadeBuf I__3864 (
            .O(N__17405),
            .I(N__17402));
    CascadeMux I__3863 (
            .O(N__17402),
            .I(N__17399));
    CascadeBuf I__3862 (
            .O(N__17399),
            .I(N__17396));
    CascadeMux I__3861 (
            .O(N__17396),
            .I(N__17393));
    CascadeBuf I__3860 (
            .O(N__17393),
            .I(N__17390));
    CascadeMux I__3859 (
            .O(N__17390),
            .I(N__17387));
    CascadeBuf I__3858 (
            .O(N__17387),
            .I(N__17384));
    CascadeMux I__3857 (
            .O(N__17384),
            .I(N__17381));
    CascadeBuf I__3856 (
            .O(N__17381),
            .I(N__17378));
    CascadeMux I__3855 (
            .O(N__17378),
            .I(N__17375));
    CascadeBuf I__3854 (
            .O(N__17375),
            .I(N__17372));
    CascadeMux I__3853 (
            .O(N__17372),
            .I(N__17369));
    CascadeBuf I__3852 (
            .O(N__17369),
            .I(N__17366));
    CascadeMux I__3851 (
            .O(N__17366),
            .I(N__17363));
    CascadeBuf I__3850 (
            .O(N__17363),
            .I(N__17360));
    CascadeMux I__3849 (
            .O(N__17360),
            .I(N__17357));
    InMux I__3848 (
            .O(N__17357),
            .I(N__17353));
    CascadeMux I__3847 (
            .O(N__17356),
            .I(N__17350));
    LocalMux I__3846 (
            .O(N__17353),
            .I(N__17347));
    InMux I__3845 (
            .O(N__17350),
            .I(N__17344));
    Span12Mux_h I__3844 (
            .O(N__17347),
            .I(N__17340));
    LocalMux I__3843 (
            .O(N__17344),
            .I(N__17337));
    InMux I__3842 (
            .O(N__17343),
            .I(N__17334));
    Span12Mux_v I__3841 (
            .O(N__17340),
            .I(N__17331));
    Odrv4 I__3840 (
            .O(N__17337),
            .I(M_this_internal_address_qZ0Z_0));
    LocalMux I__3839 (
            .O(N__17334),
            .I(M_this_internal_address_qZ0Z_0));
    Odrv12 I__3838 (
            .O(N__17331),
            .I(M_this_internal_address_qZ0Z_0));
    CascadeMux I__3837 (
            .O(N__17324),
            .I(N__17321));
    InMux I__3836 (
            .O(N__17321),
            .I(N__17318));
    LocalMux I__3835 (
            .O(N__17318),
            .I(N__17315));
    Odrv4 I__3834 (
            .O(N__17315),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_0 ));
    InMux I__3833 (
            .O(N__17312),
            .I(N__17309));
    LocalMux I__3832 (
            .O(N__17309),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_10 ));
    InMux I__3831 (
            .O(N__17306),
            .I(N__17303));
    LocalMux I__3830 (
            .O(N__17303),
            .I(un1_M_this_internal_address_q_cry_9_c_RNITQCIZ0));
    CascadeMux I__3829 (
            .O(N__17300),
            .I(N__17297));
    CascadeBuf I__3828 (
            .O(N__17297),
            .I(N__17294));
    CascadeMux I__3827 (
            .O(N__17294),
            .I(N__17291));
    CascadeBuf I__3826 (
            .O(N__17291),
            .I(N__17288));
    CascadeMux I__3825 (
            .O(N__17288),
            .I(N__17285));
    CascadeBuf I__3824 (
            .O(N__17285),
            .I(N__17282));
    CascadeMux I__3823 (
            .O(N__17282),
            .I(N__17279));
    CascadeBuf I__3822 (
            .O(N__17279),
            .I(N__17276));
    CascadeMux I__3821 (
            .O(N__17276),
            .I(N__17273));
    CascadeBuf I__3820 (
            .O(N__17273),
            .I(N__17270));
    CascadeMux I__3819 (
            .O(N__17270),
            .I(N__17267));
    CascadeBuf I__3818 (
            .O(N__17267),
            .I(N__17264));
    CascadeMux I__3817 (
            .O(N__17264),
            .I(N__17261));
    CascadeBuf I__3816 (
            .O(N__17261),
            .I(N__17258));
    CascadeMux I__3815 (
            .O(N__17258),
            .I(N__17255));
    CascadeBuf I__3814 (
            .O(N__17255),
            .I(N__17252));
    CascadeMux I__3813 (
            .O(N__17252),
            .I(N__17249));
    CascadeBuf I__3812 (
            .O(N__17249),
            .I(N__17246));
    CascadeMux I__3811 (
            .O(N__17246),
            .I(N__17243));
    CascadeBuf I__3810 (
            .O(N__17243),
            .I(N__17240));
    CascadeMux I__3809 (
            .O(N__17240),
            .I(N__17237));
    CascadeBuf I__3808 (
            .O(N__17237),
            .I(N__17234));
    CascadeMux I__3807 (
            .O(N__17234),
            .I(N__17231));
    CascadeBuf I__3806 (
            .O(N__17231),
            .I(N__17228));
    CascadeMux I__3805 (
            .O(N__17228),
            .I(N__17225));
    CascadeBuf I__3804 (
            .O(N__17225),
            .I(N__17222));
    CascadeMux I__3803 (
            .O(N__17222),
            .I(N__17219));
    CascadeBuf I__3802 (
            .O(N__17219),
            .I(N__17216));
    CascadeMux I__3801 (
            .O(N__17216),
            .I(N__17213));
    CascadeBuf I__3800 (
            .O(N__17213),
            .I(N__17210));
    CascadeMux I__3799 (
            .O(N__17210),
            .I(N__17207));
    InMux I__3798 (
            .O(N__17207),
            .I(N__17204));
    LocalMux I__3797 (
            .O(N__17204),
            .I(N__17201));
    Span4Mux_s2_v I__3796 (
            .O(N__17201),
            .I(N__17198));
    Span4Mux_h I__3795 (
            .O(N__17198),
            .I(N__17193));
    InMux I__3794 (
            .O(N__17197),
            .I(N__17190));
    InMux I__3793 (
            .O(N__17196),
            .I(N__17187));
    Span4Mux_v I__3792 (
            .O(N__17193),
            .I(N__17184));
    LocalMux I__3791 (
            .O(N__17190),
            .I(M_this_internal_address_qZ0Z_10));
    LocalMux I__3790 (
            .O(N__17187),
            .I(M_this_internal_address_qZ0Z_10));
    Odrv4 I__3789 (
            .O(N__17184),
            .I(M_this_internal_address_qZ0Z_10));
    InMux I__3788 (
            .O(N__17177),
            .I(N__17174));
    LocalMux I__3787 (
            .O(N__17174),
            .I(N__17171));
    Odrv4 I__3786 (
            .O(N__17171),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_12 ));
    InMux I__3785 (
            .O(N__17168),
            .I(N__17165));
    LocalMux I__3784 (
            .O(N__17165),
            .I(un1_M_this_internal_address_q_cry_11_c_RNI8L1DZ0));
    InMux I__3783 (
            .O(N__17162),
            .I(N__17159));
    LocalMux I__3782 (
            .O(N__17159),
            .I(un1_M_this_internal_address_q_cry_5_c_RNIE50JZ0));
    InMux I__3781 (
            .O(N__17156),
            .I(N__17153));
    LocalMux I__3780 (
            .O(N__17153),
            .I(N__17150));
    Span4Mux_h I__3779 (
            .O(N__17150),
            .I(N__17147));
    Odrv4 I__3778 (
            .O(N__17147),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_13 ));
    InMux I__3777 (
            .O(N__17144),
            .I(N__17141));
    LocalMux I__3776 (
            .O(N__17141),
            .I(un1_M_this_internal_address_q_cry_12_c_RNIAO2DZ0));
    InMux I__3775 (
            .O(N__17138),
            .I(N__17135));
    LocalMux I__3774 (
            .O(N__17135),
            .I(un1_M_this_internal_address_q_cry_7_c_RNIIB2JZ0));
    CascadeMux I__3773 (
            .O(N__17132),
            .I(N__17129));
    CascadeBuf I__3772 (
            .O(N__17129),
            .I(N__17126));
    CascadeMux I__3771 (
            .O(N__17126),
            .I(N__17123));
    CascadeBuf I__3770 (
            .O(N__17123),
            .I(N__17120));
    CascadeMux I__3769 (
            .O(N__17120),
            .I(N__17117));
    CascadeBuf I__3768 (
            .O(N__17117),
            .I(N__17114));
    CascadeMux I__3767 (
            .O(N__17114),
            .I(N__17111));
    CascadeBuf I__3766 (
            .O(N__17111),
            .I(N__17108));
    CascadeMux I__3765 (
            .O(N__17108),
            .I(N__17105));
    CascadeBuf I__3764 (
            .O(N__17105),
            .I(N__17102));
    CascadeMux I__3763 (
            .O(N__17102),
            .I(N__17099));
    CascadeBuf I__3762 (
            .O(N__17099),
            .I(N__17096));
    CascadeMux I__3761 (
            .O(N__17096),
            .I(N__17093));
    CascadeBuf I__3760 (
            .O(N__17093),
            .I(N__17090));
    CascadeMux I__3759 (
            .O(N__17090),
            .I(N__17087));
    CascadeBuf I__3758 (
            .O(N__17087),
            .I(N__17084));
    CascadeMux I__3757 (
            .O(N__17084),
            .I(N__17081));
    CascadeBuf I__3756 (
            .O(N__17081),
            .I(N__17078));
    CascadeMux I__3755 (
            .O(N__17078),
            .I(N__17075));
    CascadeBuf I__3754 (
            .O(N__17075),
            .I(N__17072));
    CascadeMux I__3753 (
            .O(N__17072),
            .I(N__17069));
    CascadeBuf I__3752 (
            .O(N__17069),
            .I(N__17066));
    CascadeMux I__3751 (
            .O(N__17066),
            .I(N__17063));
    CascadeBuf I__3750 (
            .O(N__17063),
            .I(N__17060));
    CascadeMux I__3749 (
            .O(N__17060),
            .I(N__17057));
    CascadeBuf I__3748 (
            .O(N__17057),
            .I(N__17054));
    CascadeMux I__3747 (
            .O(N__17054),
            .I(N__17051));
    CascadeBuf I__3746 (
            .O(N__17051),
            .I(N__17048));
    CascadeMux I__3745 (
            .O(N__17048),
            .I(N__17045));
    CascadeBuf I__3744 (
            .O(N__17045),
            .I(N__17042));
    CascadeMux I__3743 (
            .O(N__17042),
            .I(N__17039));
    InMux I__3742 (
            .O(N__17039),
            .I(N__17036));
    LocalMux I__3741 (
            .O(N__17036),
            .I(N__17032));
    InMux I__3740 (
            .O(N__17035),
            .I(N__17028));
    Span12Mux_h I__3739 (
            .O(N__17032),
            .I(N__17025));
    InMux I__3738 (
            .O(N__17031),
            .I(N__17022));
    LocalMux I__3737 (
            .O(N__17028),
            .I(N__17017));
    Span12Mux_v I__3736 (
            .O(N__17025),
            .I(N__17017));
    LocalMux I__3735 (
            .O(N__17022),
            .I(M_this_internal_address_qZ0Z_3));
    Odrv12 I__3734 (
            .O(N__17017),
            .I(M_this_internal_address_qZ0Z_3));
    CascadeMux I__3733 (
            .O(N__17012),
            .I(N__17009));
    InMux I__3732 (
            .O(N__17009),
            .I(N__17006));
    LocalMux I__3731 (
            .O(N__17006),
            .I(un1_M_this_internal_address_q_cry_2_c_RNI8SSIZ0));
    InMux I__3730 (
            .O(N__17003),
            .I(un1_M_this_internal_address_q_cry_2));
    CascadeMux I__3729 (
            .O(N__17000),
            .I(N__16997));
    CascadeBuf I__3728 (
            .O(N__16997),
            .I(N__16994));
    CascadeMux I__3727 (
            .O(N__16994),
            .I(N__16991));
    CascadeBuf I__3726 (
            .O(N__16991),
            .I(N__16988));
    CascadeMux I__3725 (
            .O(N__16988),
            .I(N__16985));
    CascadeBuf I__3724 (
            .O(N__16985),
            .I(N__16982));
    CascadeMux I__3723 (
            .O(N__16982),
            .I(N__16979));
    CascadeBuf I__3722 (
            .O(N__16979),
            .I(N__16976));
    CascadeMux I__3721 (
            .O(N__16976),
            .I(N__16973));
    CascadeBuf I__3720 (
            .O(N__16973),
            .I(N__16970));
    CascadeMux I__3719 (
            .O(N__16970),
            .I(N__16967));
    CascadeBuf I__3718 (
            .O(N__16967),
            .I(N__16964));
    CascadeMux I__3717 (
            .O(N__16964),
            .I(N__16961));
    CascadeBuf I__3716 (
            .O(N__16961),
            .I(N__16958));
    CascadeMux I__3715 (
            .O(N__16958),
            .I(N__16955));
    CascadeBuf I__3714 (
            .O(N__16955),
            .I(N__16952));
    CascadeMux I__3713 (
            .O(N__16952),
            .I(N__16949));
    CascadeBuf I__3712 (
            .O(N__16949),
            .I(N__16946));
    CascadeMux I__3711 (
            .O(N__16946),
            .I(N__16943));
    CascadeBuf I__3710 (
            .O(N__16943),
            .I(N__16940));
    CascadeMux I__3709 (
            .O(N__16940),
            .I(N__16937));
    CascadeBuf I__3708 (
            .O(N__16937),
            .I(N__16934));
    CascadeMux I__3707 (
            .O(N__16934),
            .I(N__16931));
    CascadeBuf I__3706 (
            .O(N__16931),
            .I(N__16928));
    CascadeMux I__3705 (
            .O(N__16928),
            .I(N__16925));
    CascadeBuf I__3704 (
            .O(N__16925),
            .I(N__16922));
    CascadeMux I__3703 (
            .O(N__16922),
            .I(N__16919));
    CascadeBuf I__3702 (
            .O(N__16919),
            .I(N__16916));
    CascadeMux I__3701 (
            .O(N__16916),
            .I(N__16913));
    CascadeBuf I__3700 (
            .O(N__16913),
            .I(N__16910));
    CascadeMux I__3699 (
            .O(N__16910),
            .I(N__16907));
    InMux I__3698 (
            .O(N__16907),
            .I(N__16904));
    LocalMux I__3697 (
            .O(N__16904),
            .I(N__16901));
    Span4Mux_h I__3696 (
            .O(N__16901),
            .I(N__16898));
    Span4Mux_h I__3695 (
            .O(N__16898),
            .I(N__16893));
    InMux I__3694 (
            .O(N__16897),
            .I(N__16890));
    InMux I__3693 (
            .O(N__16896),
            .I(N__16887));
    Sp12to4 I__3692 (
            .O(N__16893),
            .I(N__16884));
    LocalMux I__3691 (
            .O(N__16890),
            .I(M_this_internal_address_qZ0Z_4));
    LocalMux I__3690 (
            .O(N__16887),
            .I(M_this_internal_address_qZ0Z_4));
    Odrv12 I__3689 (
            .O(N__16884),
            .I(M_this_internal_address_qZ0Z_4));
    InMux I__3688 (
            .O(N__16877),
            .I(N__16874));
    LocalMux I__3687 (
            .O(N__16874),
            .I(un1_M_this_internal_address_q_cry_3_c_RNIAVTIZ0));
    InMux I__3686 (
            .O(N__16871),
            .I(un1_M_this_internal_address_q_cry_3));
    CascadeMux I__3685 (
            .O(N__16868),
            .I(N__16865));
    CascadeBuf I__3684 (
            .O(N__16865),
            .I(N__16862));
    CascadeMux I__3683 (
            .O(N__16862),
            .I(N__16859));
    CascadeBuf I__3682 (
            .O(N__16859),
            .I(N__16856));
    CascadeMux I__3681 (
            .O(N__16856),
            .I(N__16853));
    CascadeBuf I__3680 (
            .O(N__16853),
            .I(N__16850));
    CascadeMux I__3679 (
            .O(N__16850),
            .I(N__16847));
    CascadeBuf I__3678 (
            .O(N__16847),
            .I(N__16844));
    CascadeMux I__3677 (
            .O(N__16844),
            .I(N__16841));
    CascadeBuf I__3676 (
            .O(N__16841),
            .I(N__16838));
    CascadeMux I__3675 (
            .O(N__16838),
            .I(N__16835));
    CascadeBuf I__3674 (
            .O(N__16835),
            .I(N__16832));
    CascadeMux I__3673 (
            .O(N__16832),
            .I(N__16829));
    CascadeBuf I__3672 (
            .O(N__16829),
            .I(N__16826));
    CascadeMux I__3671 (
            .O(N__16826),
            .I(N__16823));
    CascadeBuf I__3670 (
            .O(N__16823),
            .I(N__16820));
    CascadeMux I__3669 (
            .O(N__16820),
            .I(N__16817));
    CascadeBuf I__3668 (
            .O(N__16817),
            .I(N__16814));
    CascadeMux I__3667 (
            .O(N__16814),
            .I(N__16811));
    CascadeBuf I__3666 (
            .O(N__16811),
            .I(N__16808));
    CascadeMux I__3665 (
            .O(N__16808),
            .I(N__16805));
    CascadeBuf I__3664 (
            .O(N__16805),
            .I(N__16802));
    CascadeMux I__3663 (
            .O(N__16802),
            .I(N__16799));
    CascadeBuf I__3662 (
            .O(N__16799),
            .I(N__16796));
    CascadeMux I__3661 (
            .O(N__16796),
            .I(N__16793));
    CascadeBuf I__3660 (
            .O(N__16793),
            .I(N__16790));
    CascadeMux I__3659 (
            .O(N__16790),
            .I(N__16787));
    CascadeBuf I__3658 (
            .O(N__16787),
            .I(N__16784));
    CascadeMux I__3657 (
            .O(N__16784),
            .I(N__16781));
    CascadeBuf I__3656 (
            .O(N__16781),
            .I(N__16778));
    CascadeMux I__3655 (
            .O(N__16778),
            .I(N__16775));
    InMux I__3654 (
            .O(N__16775),
            .I(N__16772));
    LocalMux I__3653 (
            .O(N__16772),
            .I(N__16769));
    Span4Mux_s2_v I__3652 (
            .O(N__16769),
            .I(N__16766));
    Sp12to4 I__3651 (
            .O(N__16766),
            .I(N__16761));
    InMux I__3650 (
            .O(N__16765),
            .I(N__16758));
    InMux I__3649 (
            .O(N__16764),
            .I(N__16755));
    Span12Mux_h I__3648 (
            .O(N__16761),
            .I(N__16752));
    LocalMux I__3647 (
            .O(N__16758),
            .I(M_this_internal_address_qZ0Z_5));
    LocalMux I__3646 (
            .O(N__16755),
            .I(M_this_internal_address_qZ0Z_5));
    Odrv12 I__3645 (
            .O(N__16752),
            .I(M_this_internal_address_qZ0Z_5));
    InMux I__3644 (
            .O(N__16745),
            .I(N__16742));
    LocalMux I__3643 (
            .O(N__16742),
            .I(un1_M_this_internal_address_q_cry_4_c_RNIC2VIZ0));
    InMux I__3642 (
            .O(N__16739),
            .I(un1_M_this_internal_address_q_cry_4));
    InMux I__3641 (
            .O(N__16736),
            .I(un1_M_this_internal_address_q_cry_5));
    CascadeMux I__3640 (
            .O(N__16733),
            .I(N__16730));
    CascadeBuf I__3639 (
            .O(N__16730),
            .I(N__16727));
    CascadeMux I__3638 (
            .O(N__16727),
            .I(N__16724));
    CascadeBuf I__3637 (
            .O(N__16724),
            .I(N__16721));
    CascadeMux I__3636 (
            .O(N__16721),
            .I(N__16718));
    CascadeBuf I__3635 (
            .O(N__16718),
            .I(N__16715));
    CascadeMux I__3634 (
            .O(N__16715),
            .I(N__16712));
    CascadeBuf I__3633 (
            .O(N__16712),
            .I(N__16709));
    CascadeMux I__3632 (
            .O(N__16709),
            .I(N__16706));
    CascadeBuf I__3631 (
            .O(N__16706),
            .I(N__16703));
    CascadeMux I__3630 (
            .O(N__16703),
            .I(N__16700));
    CascadeBuf I__3629 (
            .O(N__16700),
            .I(N__16697));
    CascadeMux I__3628 (
            .O(N__16697),
            .I(N__16694));
    CascadeBuf I__3627 (
            .O(N__16694),
            .I(N__16691));
    CascadeMux I__3626 (
            .O(N__16691),
            .I(N__16688));
    CascadeBuf I__3625 (
            .O(N__16688),
            .I(N__16685));
    CascadeMux I__3624 (
            .O(N__16685),
            .I(N__16682));
    CascadeBuf I__3623 (
            .O(N__16682),
            .I(N__16679));
    CascadeMux I__3622 (
            .O(N__16679),
            .I(N__16676));
    CascadeBuf I__3621 (
            .O(N__16676),
            .I(N__16673));
    CascadeMux I__3620 (
            .O(N__16673),
            .I(N__16670));
    CascadeBuf I__3619 (
            .O(N__16670),
            .I(N__16667));
    CascadeMux I__3618 (
            .O(N__16667),
            .I(N__16664));
    CascadeBuf I__3617 (
            .O(N__16664),
            .I(N__16661));
    CascadeMux I__3616 (
            .O(N__16661),
            .I(N__16658));
    CascadeBuf I__3615 (
            .O(N__16658),
            .I(N__16655));
    CascadeMux I__3614 (
            .O(N__16655),
            .I(N__16652));
    CascadeBuf I__3613 (
            .O(N__16652),
            .I(N__16649));
    CascadeMux I__3612 (
            .O(N__16649),
            .I(N__16646));
    CascadeBuf I__3611 (
            .O(N__16646),
            .I(N__16643));
    CascadeMux I__3610 (
            .O(N__16643),
            .I(N__16640));
    InMux I__3609 (
            .O(N__16640),
            .I(N__16637));
    LocalMux I__3608 (
            .O(N__16637),
            .I(N__16634));
    Span12Mux_s10_h I__3607 (
            .O(N__16634),
            .I(N__16629));
    InMux I__3606 (
            .O(N__16633),
            .I(N__16626));
    InMux I__3605 (
            .O(N__16632),
            .I(N__16623));
    Span12Mux_v I__3604 (
            .O(N__16629),
            .I(N__16620));
    LocalMux I__3603 (
            .O(N__16626),
            .I(M_this_internal_address_qZ0Z_7));
    LocalMux I__3602 (
            .O(N__16623),
            .I(M_this_internal_address_qZ0Z_7));
    Odrv12 I__3601 (
            .O(N__16620),
            .I(M_this_internal_address_qZ0Z_7));
    InMux I__3600 (
            .O(N__16613),
            .I(N__16610));
    LocalMux I__3599 (
            .O(N__16610),
            .I(un1_M_this_internal_address_q_cry_6_c_RNIG81JZ0));
    InMux I__3598 (
            .O(N__16607),
            .I(un1_M_this_internal_address_q_cry_6));
    InMux I__3597 (
            .O(N__16604),
            .I(bfn_20_22_0_));
    CascadeMux I__3596 (
            .O(N__16601),
            .I(N__16598));
    CascadeBuf I__3595 (
            .O(N__16598),
            .I(N__16595));
    CascadeMux I__3594 (
            .O(N__16595),
            .I(N__16592));
    CascadeBuf I__3593 (
            .O(N__16592),
            .I(N__16589));
    CascadeMux I__3592 (
            .O(N__16589),
            .I(N__16586));
    CascadeBuf I__3591 (
            .O(N__16586),
            .I(N__16583));
    CascadeMux I__3590 (
            .O(N__16583),
            .I(N__16580));
    CascadeBuf I__3589 (
            .O(N__16580),
            .I(N__16577));
    CascadeMux I__3588 (
            .O(N__16577),
            .I(N__16574));
    CascadeBuf I__3587 (
            .O(N__16574),
            .I(N__16571));
    CascadeMux I__3586 (
            .O(N__16571),
            .I(N__16568));
    CascadeBuf I__3585 (
            .O(N__16568),
            .I(N__16565));
    CascadeMux I__3584 (
            .O(N__16565),
            .I(N__16562));
    CascadeBuf I__3583 (
            .O(N__16562),
            .I(N__16559));
    CascadeMux I__3582 (
            .O(N__16559),
            .I(N__16556));
    CascadeBuf I__3581 (
            .O(N__16556),
            .I(N__16553));
    CascadeMux I__3580 (
            .O(N__16553),
            .I(N__16550));
    CascadeBuf I__3579 (
            .O(N__16550),
            .I(N__16547));
    CascadeMux I__3578 (
            .O(N__16547),
            .I(N__16544));
    CascadeBuf I__3577 (
            .O(N__16544),
            .I(N__16541));
    CascadeMux I__3576 (
            .O(N__16541),
            .I(N__16538));
    CascadeBuf I__3575 (
            .O(N__16538),
            .I(N__16535));
    CascadeMux I__3574 (
            .O(N__16535),
            .I(N__16532));
    CascadeBuf I__3573 (
            .O(N__16532),
            .I(N__16529));
    CascadeMux I__3572 (
            .O(N__16529),
            .I(N__16526));
    CascadeBuf I__3571 (
            .O(N__16526),
            .I(N__16523));
    CascadeMux I__3570 (
            .O(N__16523),
            .I(N__16520));
    CascadeBuf I__3569 (
            .O(N__16520),
            .I(N__16517));
    CascadeMux I__3568 (
            .O(N__16517),
            .I(N__16514));
    CascadeBuf I__3567 (
            .O(N__16514),
            .I(N__16511));
    CascadeMux I__3566 (
            .O(N__16511),
            .I(N__16508));
    InMux I__3565 (
            .O(N__16508),
            .I(N__16505));
    LocalMux I__3564 (
            .O(N__16505),
            .I(N__16502));
    Span4Mux_s3_v I__3563 (
            .O(N__16502),
            .I(N__16499));
    Sp12to4 I__3562 (
            .O(N__16499),
            .I(N__16494));
    InMux I__3561 (
            .O(N__16498),
            .I(N__16491));
    InMux I__3560 (
            .O(N__16497),
            .I(N__16488));
    Span12Mux_h I__3559 (
            .O(N__16494),
            .I(N__16485));
    LocalMux I__3558 (
            .O(N__16491),
            .I(M_this_internal_address_qZ0Z_9));
    LocalMux I__3557 (
            .O(N__16488),
            .I(M_this_internal_address_qZ0Z_9));
    Odrv12 I__3556 (
            .O(N__16485),
            .I(M_this_internal_address_qZ0Z_9));
    InMux I__3555 (
            .O(N__16478),
            .I(N__16475));
    LocalMux I__3554 (
            .O(N__16475),
            .I(un1_M_this_internal_address_q_cry_8_c_RNIKE3JZ0));
    InMux I__3553 (
            .O(N__16472),
            .I(un1_M_this_internal_address_q_cry_8));
    InMux I__3552 (
            .O(N__16469),
            .I(un1_M_this_internal_address_q_cry_9));
    InMux I__3551 (
            .O(N__16466),
            .I(N__16463));
    LocalMux I__3550 (
            .O(N__16463),
            .I(N__16460));
    Odrv12 I__3549 (
            .O(N__16460),
            .I(M_this_vga_signals_address_13));
    InMux I__3548 (
            .O(N__16457),
            .I(N__16454));
    LocalMux I__3547 (
            .O(N__16454),
            .I(N__16451));
    Sp12to4 I__3546 (
            .O(N__16451),
            .I(N__16448));
    Odrv12 I__3545 (
            .O(N__16448),
            .I(M_this_vga_signals_address_12));
    InMux I__3544 (
            .O(N__16445),
            .I(N__16442));
    LocalMux I__3543 (
            .O(N__16442),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_5 ));
    InMux I__3542 (
            .O(N__16439),
            .I(N__16436));
    LocalMux I__3541 (
            .O(N__16436),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_3 ));
    CascadeMux I__3540 (
            .O(N__16433),
            .I(N__16430));
    InMux I__3539 (
            .O(N__16430),
            .I(N__16427));
    LocalMux I__3538 (
            .O(N__16427),
            .I(N__16424));
    Odrv4 I__3537 (
            .O(N__16424),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_7 ));
    CascadeMux I__3536 (
            .O(N__16421),
            .I(N__16417));
    InMux I__3535 (
            .O(N__16420),
            .I(N__16414));
    InMux I__3534 (
            .O(N__16417),
            .I(N__16411));
    LocalMux I__3533 (
            .O(N__16414),
            .I(N_346_0));
    LocalMux I__3532 (
            .O(N__16411),
            .I(N_346_0));
    InMux I__3531 (
            .O(N__16406),
            .I(N__16403));
    LocalMux I__3530 (
            .O(N__16403),
            .I(M_this_internal_address_q_RNI6EA12Z0Z_0));
    CascadeMux I__3529 (
            .O(N__16400),
            .I(N__16397));
    CascadeBuf I__3528 (
            .O(N__16397),
            .I(N__16394));
    CascadeMux I__3527 (
            .O(N__16394),
            .I(N__16391));
    CascadeBuf I__3526 (
            .O(N__16391),
            .I(N__16388));
    CascadeMux I__3525 (
            .O(N__16388),
            .I(N__16385));
    CascadeBuf I__3524 (
            .O(N__16385),
            .I(N__16382));
    CascadeMux I__3523 (
            .O(N__16382),
            .I(N__16379));
    CascadeBuf I__3522 (
            .O(N__16379),
            .I(N__16376));
    CascadeMux I__3521 (
            .O(N__16376),
            .I(N__16373));
    CascadeBuf I__3520 (
            .O(N__16373),
            .I(N__16370));
    CascadeMux I__3519 (
            .O(N__16370),
            .I(N__16367));
    CascadeBuf I__3518 (
            .O(N__16367),
            .I(N__16364));
    CascadeMux I__3517 (
            .O(N__16364),
            .I(N__16361));
    CascadeBuf I__3516 (
            .O(N__16361),
            .I(N__16358));
    CascadeMux I__3515 (
            .O(N__16358),
            .I(N__16355));
    CascadeBuf I__3514 (
            .O(N__16355),
            .I(N__16352));
    CascadeMux I__3513 (
            .O(N__16352),
            .I(N__16349));
    CascadeBuf I__3512 (
            .O(N__16349),
            .I(N__16346));
    CascadeMux I__3511 (
            .O(N__16346),
            .I(N__16343));
    CascadeBuf I__3510 (
            .O(N__16343),
            .I(N__16340));
    CascadeMux I__3509 (
            .O(N__16340),
            .I(N__16337));
    CascadeBuf I__3508 (
            .O(N__16337),
            .I(N__16334));
    CascadeMux I__3507 (
            .O(N__16334),
            .I(N__16331));
    CascadeBuf I__3506 (
            .O(N__16331),
            .I(N__16328));
    CascadeMux I__3505 (
            .O(N__16328),
            .I(N__16325));
    CascadeBuf I__3504 (
            .O(N__16325),
            .I(N__16322));
    CascadeMux I__3503 (
            .O(N__16322),
            .I(N__16319));
    CascadeBuf I__3502 (
            .O(N__16319),
            .I(N__16316));
    CascadeMux I__3501 (
            .O(N__16316),
            .I(N__16313));
    CascadeBuf I__3500 (
            .O(N__16313),
            .I(N__16310));
    CascadeMux I__3499 (
            .O(N__16310),
            .I(N__16307));
    InMux I__3498 (
            .O(N__16307),
            .I(N__16304));
    LocalMux I__3497 (
            .O(N__16304),
            .I(N__16300));
    InMux I__3496 (
            .O(N__16303),
            .I(N__16297));
    Span4Mux_s3_v I__3495 (
            .O(N__16300),
            .I(N__16294));
    LocalMux I__3494 (
            .O(N__16297),
            .I(N__16291));
    Span4Mux_h I__3493 (
            .O(N__16294),
            .I(N__16287));
    Span4Mux_h I__3492 (
            .O(N__16291),
            .I(N__16284));
    InMux I__3491 (
            .O(N__16290),
            .I(N__16281));
    Span4Mux_v I__3490 (
            .O(N__16287),
            .I(N__16278));
    Odrv4 I__3489 (
            .O(N__16284),
            .I(M_this_internal_address_qZ0Z_1));
    LocalMux I__3488 (
            .O(N__16281),
            .I(M_this_internal_address_qZ0Z_1));
    Odrv4 I__3487 (
            .O(N__16278),
            .I(M_this_internal_address_qZ0Z_1));
    InMux I__3486 (
            .O(N__16271),
            .I(N__16268));
    LocalMux I__3485 (
            .O(N__16268),
            .I(N__16265));
    Span4Mux_v I__3484 (
            .O(N__16265),
            .I(N__16262));
    Odrv4 I__3483 (
            .O(N__16262),
            .I(un1_M_this_internal_address_q_cry_0_c_RNI4MQIZ0));
    InMux I__3482 (
            .O(N__16259),
            .I(un1_M_this_internal_address_q_cry_0));
    CascadeMux I__3481 (
            .O(N__16256),
            .I(N__16253));
    CascadeBuf I__3480 (
            .O(N__16253),
            .I(N__16250));
    CascadeMux I__3479 (
            .O(N__16250),
            .I(N__16247));
    CascadeBuf I__3478 (
            .O(N__16247),
            .I(N__16244));
    CascadeMux I__3477 (
            .O(N__16244),
            .I(N__16241));
    CascadeBuf I__3476 (
            .O(N__16241),
            .I(N__16238));
    CascadeMux I__3475 (
            .O(N__16238),
            .I(N__16235));
    CascadeBuf I__3474 (
            .O(N__16235),
            .I(N__16232));
    CascadeMux I__3473 (
            .O(N__16232),
            .I(N__16229));
    CascadeBuf I__3472 (
            .O(N__16229),
            .I(N__16226));
    CascadeMux I__3471 (
            .O(N__16226),
            .I(N__16223));
    CascadeBuf I__3470 (
            .O(N__16223),
            .I(N__16220));
    CascadeMux I__3469 (
            .O(N__16220),
            .I(N__16217));
    CascadeBuf I__3468 (
            .O(N__16217),
            .I(N__16214));
    CascadeMux I__3467 (
            .O(N__16214),
            .I(N__16211));
    CascadeBuf I__3466 (
            .O(N__16211),
            .I(N__16208));
    CascadeMux I__3465 (
            .O(N__16208),
            .I(N__16205));
    CascadeBuf I__3464 (
            .O(N__16205),
            .I(N__16202));
    CascadeMux I__3463 (
            .O(N__16202),
            .I(N__16199));
    CascadeBuf I__3462 (
            .O(N__16199),
            .I(N__16196));
    CascadeMux I__3461 (
            .O(N__16196),
            .I(N__16193));
    CascadeBuf I__3460 (
            .O(N__16193),
            .I(N__16190));
    CascadeMux I__3459 (
            .O(N__16190),
            .I(N__16187));
    CascadeBuf I__3458 (
            .O(N__16187),
            .I(N__16184));
    CascadeMux I__3457 (
            .O(N__16184),
            .I(N__16181));
    CascadeBuf I__3456 (
            .O(N__16181),
            .I(N__16178));
    CascadeMux I__3455 (
            .O(N__16178),
            .I(N__16175));
    CascadeBuf I__3454 (
            .O(N__16175),
            .I(N__16172));
    CascadeMux I__3453 (
            .O(N__16172),
            .I(N__16169));
    CascadeBuf I__3452 (
            .O(N__16169),
            .I(N__16166));
    CascadeMux I__3451 (
            .O(N__16166),
            .I(N__16163));
    InMux I__3450 (
            .O(N__16163),
            .I(N__16160));
    LocalMux I__3449 (
            .O(N__16160),
            .I(N__16157));
    Span4Mux_h I__3448 (
            .O(N__16157),
            .I(N__16154));
    Sp12to4 I__3447 (
            .O(N__16154),
            .I(N__16149));
    InMux I__3446 (
            .O(N__16153),
            .I(N__16146));
    InMux I__3445 (
            .O(N__16152),
            .I(N__16143));
    Span12Mux_s10_v I__3444 (
            .O(N__16149),
            .I(N__16140));
    LocalMux I__3443 (
            .O(N__16146),
            .I(M_this_internal_address_qZ0Z_2));
    LocalMux I__3442 (
            .O(N__16143),
            .I(M_this_internal_address_qZ0Z_2));
    Odrv12 I__3441 (
            .O(N__16140),
            .I(M_this_internal_address_qZ0Z_2));
    CascadeMux I__3440 (
            .O(N__16133),
            .I(N__16130));
    InMux I__3439 (
            .O(N__16130),
            .I(N__16127));
    LocalMux I__3438 (
            .O(N__16127),
            .I(N__16124));
    Odrv4 I__3437 (
            .O(N__16124),
            .I(un1_M_this_internal_address_q_cry_1_c_RNI6PRIZ0));
    InMux I__3436 (
            .O(N__16121),
            .I(un1_M_this_internal_address_q_cry_1));
    InMux I__3435 (
            .O(N__16118),
            .I(N__16115));
    LocalMux I__3434 (
            .O(N__16115),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_9 ));
    InMux I__3433 (
            .O(N__16112),
            .I(N__16109));
    LocalMux I__3432 (
            .O(N__16109),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_2 ));
    InMux I__3431 (
            .O(N__16106),
            .I(N__16102));
    InMux I__3430 (
            .O(N__16105),
            .I(N__16099));
    LocalMux I__3429 (
            .O(N__16102),
            .I(\this_start_data_delay.N_407 ));
    LocalMux I__3428 (
            .O(N__16099),
            .I(\this_start_data_delay.N_407 ));
    InMux I__3427 (
            .O(N__16094),
            .I(N__16087));
    InMux I__3426 (
            .O(N__16093),
            .I(N__16087));
    InMux I__3425 (
            .O(N__16092),
            .I(N__16084));
    LocalMux I__3424 (
            .O(N__16087),
            .I(\this_start_data_delay.N_398 ));
    LocalMux I__3423 (
            .O(N__16084),
            .I(\this_start_data_delay.N_398 ));
    InMux I__3422 (
            .O(N__16079),
            .I(N__16076));
    LocalMux I__3421 (
            .O(N__16076),
            .I(\this_start_data_delay.M_this_state_dZ0Z29 ));
    InMux I__3420 (
            .O(N__16073),
            .I(N__16070));
    LocalMux I__3419 (
            .O(N__16070),
            .I(N__16067));
    Span4Mux_v I__3418 (
            .O(N__16067),
            .I(N__16064));
    Odrv4 I__3417 (
            .O(N__16064),
            .I(\this_start_data_delay.N_396 ));
    InMux I__3416 (
            .O(N__16061),
            .I(N__16058));
    LocalMux I__3415 (
            .O(N__16058),
            .I(\this_start_data_delay.M_this_state_dZ0Z27 ));
    CascadeMux I__3414 (
            .O(N__16055),
            .I(N__16049));
    CascadeMux I__3413 (
            .O(N__16054),
            .I(N__16046));
    InMux I__3412 (
            .O(N__16053),
            .I(N__16041));
    InMux I__3411 (
            .O(N__16052),
            .I(N__16041));
    InMux I__3410 (
            .O(N__16049),
            .I(N__16036));
    InMux I__3409 (
            .O(N__16046),
            .I(N__16036));
    LocalMux I__3408 (
            .O(N__16041),
            .I(N__16031));
    LocalMux I__3407 (
            .O(N__16036),
            .I(N__16031));
    Span12Mux_h I__3406 (
            .O(N__16031),
            .I(N__16028));
    Odrv12 I__3405 (
            .O(N__16028),
            .I(port_address_in_0));
    InMux I__3404 (
            .O(N__16025),
            .I(N__16017));
    InMux I__3403 (
            .O(N__16024),
            .I(N__16017));
    InMux I__3402 (
            .O(N__16023),
            .I(N__16012));
    InMux I__3401 (
            .O(N__16022),
            .I(N__16012));
    LocalMux I__3400 (
            .O(N__16017),
            .I(N__16007));
    LocalMux I__3399 (
            .O(N__16012),
            .I(N__16007));
    Span12Mux_h I__3398 (
            .O(N__16007),
            .I(N__16004));
    Odrv12 I__3397 (
            .O(N__16004),
            .I(port_address_in_1));
    InMux I__3396 (
            .O(N__16001),
            .I(N__15998));
    LocalMux I__3395 (
            .O(N__15998),
            .I(\this_start_data_delay.M_this_state_dZ0Z28 ));
    InMux I__3394 (
            .O(N__15995),
            .I(N__15991));
    InMux I__3393 (
            .O(N__15994),
            .I(N__15988));
    LocalMux I__3392 (
            .O(N__15991),
            .I(M_this_state_qZ0Z_6));
    LocalMux I__3391 (
            .O(N__15988),
            .I(M_this_state_qZ0Z_6));
    InMux I__3390 (
            .O(N__15983),
            .I(N__15980));
    LocalMux I__3389 (
            .O(N__15980),
            .I(N__15972));
    InMux I__3388 (
            .O(N__15979),
            .I(N__15967));
    InMux I__3387 (
            .O(N__15978),
            .I(N__15967));
    InMux I__3386 (
            .O(N__15977),
            .I(N__15964));
    InMux I__3385 (
            .O(N__15976),
            .I(N__15959));
    InMux I__3384 (
            .O(N__15975),
            .I(N__15959));
    Span4Mux_v I__3383 (
            .O(N__15972),
            .I(N__15956));
    LocalMux I__3382 (
            .O(N__15967),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__3381 (
            .O(N__15964),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__3380 (
            .O(N__15959),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__3379 (
            .O(N__15956),
            .I(M_this_state_qZ0Z_1));
    CascadeMux I__3378 (
            .O(N__15947),
            .I(N__15942));
    InMux I__3377 (
            .O(N__15946),
            .I(N__15939));
    InMux I__3376 (
            .O(N__15945),
            .I(N__15936));
    InMux I__3375 (
            .O(N__15942),
            .I(N__15933));
    LocalMux I__3374 (
            .O(N__15939),
            .I(M_this_state_qZ0Z_4));
    LocalMux I__3373 (
            .O(N__15936),
            .I(M_this_state_qZ0Z_4));
    LocalMux I__3372 (
            .O(N__15933),
            .I(M_this_state_qZ0Z_4));
    InMux I__3371 (
            .O(N__15926),
            .I(N__15923));
    LocalMux I__3370 (
            .O(N__15923),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_4 ));
    CascadeMux I__3369 (
            .O(N__15920),
            .I(N__15917));
    InMux I__3368 (
            .O(N__15917),
            .I(N__15914));
    LocalMux I__3367 (
            .O(N__15914),
            .I(N__15911));
    Span12Mux_s11_v I__3366 (
            .O(N__15911),
            .I(N__15908));
    Span12Mux_h I__3365 (
            .O(N__15908),
            .I(N__15904));
    InMux I__3364 (
            .O(N__15907),
            .I(N__15901));
    Odrv12 I__3363 (
            .O(N__15904),
            .I(port_rw_in));
    LocalMux I__3362 (
            .O(N__15901),
            .I(port_rw_in));
    InMux I__3361 (
            .O(N__15896),
            .I(N__15893));
    LocalMux I__3360 (
            .O(N__15893),
            .I(\this_start_data_delay.M_this_state_q_srsts_0_a2_1_4 ));
    CascadeMux I__3359 (
            .O(N__15890),
            .I(\this_start_data_delay.N_352_0_cascade_ ));
    InMux I__3358 (
            .O(N__15887),
            .I(N__15884));
    LocalMux I__3357 (
            .O(N__15884),
            .I(N__15881));
    Odrv4 I__3356 (
            .O(N__15881),
            .I(\this_start_data_delay.M_this_state_q_srsts_0_0_4 ));
    InMux I__3355 (
            .O(N__15878),
            .I(N__15866));
    InMux I__3354 (
            .O(N__15877),
            .I(N__15866));
    InMux I__3353 (
            .O(N__15876),
            .I(N__15866));
    InMux I__3352 (
            .O(N__15875),
            .I(N__15866));
    LocalMux I__3351 (
            .O(N__15866),
            .I(N__15863));
    Span12Mux_v I__3350 (
            .O(N__15863),
            .I(N__15860));
    Span12Mux_h I__3349 (
            .O(N__15860),
            .I(N__15857));
    Odrv12 I__3348 (
            .O(N__15857),
            .I(port_enb_c));
    InMux I__3347 (
            .O(N__15854),
            .I(N__15842));
    InMux I__3346 (
            .O(N__15853),
            .I(N__15842));
    InMux I__3345 (
            .O(N__15852),
            .I(N__15842));
    InMux I__3344 (
            .O(N__15851),
            .I(N__15842));
    LocalMux I__3343 (
            .O(N__15842),
            .I(M_this_delay_clk_out_0));
    CascadeMux I__3342 (
            .O(N__15839),
            .I(N__15836));
    InMux I__3341 (
            .O(N__15836),
            .I(N__15827));
    InMux I__3340 (
            .O(N__15835),
            .I(N__15827));
    InMux I__3339 (
            .O(N__15834),
            .I(N__15827));
    LocalMux I__3338 (
            .O(N__15827),
            .I(\this_start_data_delay.M_last_qZ0 ));
    InMux I__3337 (
            .O(N__15824),
            .I(N__15821));
    LocalMux I__3336 (
            .O(N__15821),
            .I(\this_start_data_delay.N_352_0 ));
    CascadeMux I__3335 (
            .O(N__15818),
            .I(\this_start_data_delay.N_407_cascade_ ));
    CascadeMux I__3334 (
            .O(N__15815),
            .I(N__15812));
    InMux I__3333 (
            .O(N__15812),
            .I(N__15809));
    LocalMux I__3332 (
            .O(N__15809),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_1 ));
    InMux I__3331 (
            .O(N__15806),
            .I(N__15803));
    LocalMux I__3330 (
            .O(N__15803),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    InMux I__3329 (
            .O(N__15800),
            .I(N__15788));
    InMux I__3328 (
            .O(N__15799),
            .I(N__15788));
    InMux I__3327 (
            .O(N__15798),
            .I(N__15788));
    InMux I__3326 (
            .O(N__15797),
            .I(N__15788));
    LocalMux I__3325 (
            .O(N__15788),
            .I(N__15785));
    Span12Mux_v I__3324 (
            .O(N__15785),
            .I(N__15782));
    Span12Mux_v I__3323 (
            .O(N__15782),
            .I(N__15779));
    Odrv12 I__3322 (
            .O(N__15779),
            .I(rst_n_c));
    InMux I__3321 (
            .O(N__15776),
            .I(N__15773));
    LocalMux I__3320 (
            .O(N__15773),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    IoInMux I__3319 (
            .O(N__15770),
            .I(N__15767));
    LocalMux I__3318 (
            .O(N__15767),
            .I(N__15763));
    InMux I__3317 (
            .O(N__15766),
            .I(N__15760));
    Span4Mux_s3_v I__3316 (
            .O(N__15763),
            .I(N__15757));
    LocalMux I__3315 (
            .O(N__15760),
            .I(N__15752));
    Span4Mux_v I__3314 (
            .O(N__15757),
            .I(N__15752));
    Odrv4 I__3313 (
            .O(N__15752),
            .I(M_this_state_q_nss_0));
    InMux I__3312 (
            .O(N__15749),
            .I(N__15746));
    LocalMux I__3311 (
            .O(N__15746),
            .I(N__15743));
    Odrv12 I__3310 (
            .O(N__15743),
            .I(\this_delay_clk.M_pipe_qZ0Z_3 ));
    CascadeMux I__3309 (
            .O(N__15740),
            .I(N__15736));
    InMux I__3308 (
            .O(N__15739),
            .I(N__15733));
    InMux I__3307 (
            .O(N__15736),
            .I(N__15730));
    LocalMux I__3306 (
            .O(N__15733),
            .I(\this_start_data_delay.N_353_0 ));
    LocalMux I__3305 (
            .O(N__15730),
            .I(\this_start_data_delay.N_353_0 ));
    CascadeMux I__3304 (
            .O(N__15725),
            .I(M_this_start_data_delay_out_0_cascade_));
    InMux I__3303 (
            .O(N__15722),
            .I(N__15719));
    LocalMux I__3302 (
            .O(N__15719),
            .I(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_11 ));
    CascadeMux I__3301 (
            .O(N__15716),
            .I(N__15713));
    InMux I__3300 (
            .O(N__15713),
            .I(N__15709));
    InMux I__3299 (
            .O(N__15712),
            .I(N__15706));
    LocalMux I__3298 (
            .O(N__15709),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__3297 (
            .O(N__15706),
            .I(M_this_data_count_qZ0Z_3));
    CascadeMux I__3296 (
            .O(N__15701),
            .I(N__15698));
    InMux I__3295 (
            .O(N__15698),
            .I(N__15694));
    InMux I__3294 (
            .O(N__15697),
            .I(N__15691));
    LocalMux I__3293 (
            .O(N__15694),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__3292 (
            .O(N__15691),
            .I(M_this_data_count_qZ0Z_1));
    CascadeMux I__3291 (
            .O(N__15686),
            .I(N__15682));
    InMux I__3290 (
            .O(N__15685),
            .I(N__15679));
    InMux I__3289 (
            .O(N__15682),
            .I(N__15676));
    LocalMux I__3288 (
            .O(N__15679),
            .I(M_this_data_count_qZ0Z_12));
    LocalMux I__3287 (
            .O(N__15676),
            .I(M_this_data_count_qZ0Z_12));
    InMux I__3286 (
            .O(N__15671),
            .I(N__15667));
    InMux I__3285 (
            .O(N__15670),
            .I(N__15664));
    LocalMux I__3284 (
            .O(N__15667),
            .I(M_this_data_count_qZ0Z_2));
    LocalMux I__3283 (
            .O(N__15664),
            .I(M_this_data_count_qZ0Z_2));
    CascadeMux I__3282 (
            .O(N__15659),
            .I(N__15655));
    InMux I__3281 (
            .O(N__15658),
            .I(N__15652));
    InMux I__3280 (
            .O(N__15655),
            .I(N__15649));
    LocalMux I__3279 (
            .O(N__15652),
            .I(N__15646));
    LocalMux I__3278 (
            .O(N__15649),
            .I(M_this_data_count_qZ0Z_13));
    Odrv4 I__3277 (
            .O(N__15646),
            .I(M_this_data_count_qZ0Z_13));
    InMux I__3276 (
            .O(N__15641),
            .I(N__15637));
    InMux I__3275 (
            .O(N__15640),
            .I(N__15634));
    LocalMux I__3274 (
            .O(N__15637),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__3273 (
            .O(N__15634),
            .I(M_this_data_count_qZ0Z_0));
    InMux I__3272 (
            .O(N__15629),
            .I(N__15626));
    LocalMux I__3271 (
            .O(N__15626),
            .I(\this_start_data_delay.M_this_state_q_srsts_i_a2_1_9Z0Z_1 ));
    CascadeMux I__3270 (
            .O(N__15623),
            .I(\this_start_data_delay.M_this_state_q_srsts_i_a2_1_6Z0Z_1_cascade_ ));
    InMux I__3269 (
            .O(N__15620),
            .I(N__15617));
    LocalMux I__3268 (
            .O(N__15617),
            .I(N__15612));
    InMux I__3267 (
            .O(N__15616),
            .I(N__15607));
    InMux I__3266 (
            .O(N__15615),
            .I(N__15607));
    Odrv4 I__3265 (
            .O(N__15612),
            .I(\this_start_data_delay.N_413 ));
    LocalMux I__3264 (
            .O(N__15607),
            .I(\this_start_data_delay.N_413 ));
    InMux I__3263 (
            .O(N__15602),
            .I(N__15598));
    InMux I__3262 (
            .O(N__15601),
            .I(N__15595));
    LocalMux I__3261 (
            .O(N__15598),
            .I(M_this_data_count_qZ0Z_6));
    LocalMux I__3260 (
            .O(N__15595),
            .I(M_this_data_count_qZ0Z_6));
    CascadeMux I__3259 (
            .O(N__15590),
            .I(N__15587));
    InMux I__3258 (
            .O(N__15587),
            .I(N__15583));
    InMux I__3257 (
            .O(N__15586),
            .I(N__15580));
    LocalMux I__3256 (
            .O(N__15583),
            .I(M_this_data_count_qZ0Z_5));
    LocalMux I__3255 (
            .O(N__15580),
            .I(M_this_data_count_qZ0Z_5));
    CascadeMux I__3254 (
            .O(N__15575),
            .I(N__15571));
    CascadeMux I__3253 (
            .O(N__15574),
            .I(N__15568));
    InMux I__3252 (
            .O(N__15571),
            .I(N__15565));
    InMux I__3251 (
            .O(N__15568),
            .I(N__15562));
    LocalMux I__3250 (
            .O(N__15565),
            .I(M_this_data_count_qZ0Z_7));
    LocalMux I__3249 (
            .O(N__15562),
            .I(M_this_data_count_qZ0Z_7));
    InMux I__3248 (
            .O(N__15557),
            .I(N__15553));
    InMux I__3247 (
            .O(N__15556),
            .I(N__15550));
    LocalMux I__3246 (
            .O(N__15553),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__3245 (
            .O(N__15550),
            .I(M_this_data_count_qZ0Z_4));
    InMux I__3244 (
            .O(N__15545),
            .I(N__15542));
    LocalMux I__3243 (
            .O(N__15542),
            .I(\this_start_data_delay.M_this_state_q_srsts_i_a2_1_8Z0Z_1 ));
    InMux I__3242 (
            .O(N__15539),
            .I(N__15535));
    InMux I__3241 (
            .O(N__15538),
            .I(N__15532));
    LocalMux I__3240 (
            .O(N__15535),
            .I(M_this_data_count_qZ0Z_10));
    LocalMux I__3239 (
            .O(N__15532),
            .I(M_this_data_count_qZ0Z_10));
    InMux I__3238 (
            .O(N__15527),
            .I(N__15523));
    InMux I__3237 (
            .O(N__15526),
            .I(N__15520));
    LocalMux I__3236 (
            .O(N__15523),
            .I(M_this_data_count_qZ0Z_8));
    LocalMux I__3235 (
            .O(N__15520),
            .I(M_this_data_count_qZ0Z_8));
    CascadeMux I__3234 (
            .O(N__15515),
            .I(N__15511));
    InMux I__3233 (
            .O(N__15514),
            .I(N__15508));
    InMux I__3232 (
            .O(N__15511),
            .I(N__15505));
    LocalMux I__3231 (
            .O(N__15508),
            .I(M_this_data_count_qZ0Z_11));
    LocalMux I__3230 (
            .O(N__15505),
            .I(M_this_data_count_qZ0Z_11));
    InMux I__3229 (
            .O(N__15500),
            .I(N__15496));
    InMux I__3228 (
            .O(N__15499),
            .I(N__15493));
    LocalMux I__3227 (
            .O(N__15496),
            .I(M_this_data_count_qZ0Z_9));
    LocalMux I__3226 (
            .O(N__15493),
            .I(M_this_data_count_qZ0Z_9));
    InMux I__3225 (
            .O(N__15488),
            .I(N__15485));
    LocalMux I__3224 (
            .O(N__15485),
            .I(\this_start_data_delay.M_this_state_q_srsts_i_a2_1_7Z0Z_1 ));
    SRMux I__3223 (
            .O(N__15482),
            .I(N__15479));
    LocalMux I__3222 (
            .O(N__15479),
            .I(N__15475));
    SRMux I__3221 (
            .O(N__15478),
            .I(N__15472));
    Span4Mux_h I__3220 (
            .O(N__15475),
            .I(N__15467));
    LocalMux I__3219 (
            .O(N__15472),
            .I(N__15467));
    Odrv4 I__3218 (
            .O(N__15467),
            .I(M_this_state_q_RNI20CEZ0Z_0));
    InMux I__3217 (
            .O(N__15464),
            .I(N__15461));
    LocalMux I__3216 (
            .O(N__15461),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    InMux I__3215 (
            .O(N__15458),
            .I(N__15453));
    InMux I__3214 (
            .O(N__15457),
            .I(N__15448));
    InMux I__3213 (
            .O(N__15456),
            .I(N__15448));
    LocalMux I__3212 (
            .O(N__15453),
            .I(N__15442));
    LocalMux I__3211 (
            .O(N__15448),
            .I(N__15439));
    InMux I__3210 (
            .O(N__15447),
            .I(N__15436));
    InMux I__3209 (
            .O(N__15446),
            .I(N__15432));
    InMux I__3208 (
            .O(N__15445),
            .I(N__15429));
    Span4Mux_v I__3207 (
            .O(N__15442),
            .I(N__15422));
    Span4Mux_v I__3206 (
            .O(N__15439),
            .I(N__15422));
    LocalMux I__3205 (
            .O(N__15436),
            .I(N__15422));
    InMux I__3204 (
            .O(N__15435),
            .I(N__15419));
    LocalMux I__3203 (
            .O(N__15432),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__3202 (
            .O(N__15429),
            .I(\this_vga_signals.vaddress_c2 ));
    Odrv4 I__3201 (
            .O(N__15422),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__3200 (
            .O(N__15419),
            .I(\this_vga_signals.vaddress_c2 ));
    InMux I__3199 (
            .O(N__15410),
            .I(N__15406));
    CascadeMux I__3198 (
            .O(N__15409),
            .I(N__15403));
    LocalMux I__3197 (
            .O(N__15406),
            .I(N__15400));
    InMux I__3196 (
            .O(N__15403),
            .I(N__15397));
    Odrv4 I__3195 (
            .O(N__15400),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_1 ));
    LocalMux I__3194 (
            .O(N__15397),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_1 ));
    CascadeMux I__3193 (
            .O(N__15392),
            .I(N__15388));
    InMux I__3192 (
            .O(N__15391),
            .I(N__15385));
    InMux I__3191 (
            .O(N__15388),
            .I(N__15378));
    LocalMux I__3190 (
            .O(N__15385),
            .I(N__15375));
    InMux I__3189 (
            .O(N__15384),
            .I(N__15368));
    InMux I__3188 (
            .O(N__15383),
            .I(N__15368));
    InMux I__3187 (
            .O(N__15382),
            .I(N__15368));
    CascadeMux I__3186 (
            .O(N__15381),
            .I(N__15365));
    LocalMux I__3185 (
            .O(N__15378),
            .I(N__15362));
    Span4Mux_h I__3184 (
            .O(N__15375),
            .I(N__15359));
    LocalMux I__3183 (
            .O(N__15368),
            .I(N__15356));
    InMux I__3182 (
            .O(N__15365),
            .I(N__15353));
    Odrv4 I__3181 (
            .O(N__15362),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    Odrv4 I__3180 (
            .O(N__15359),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    Odrv4 I__3179 (
            .O(N__15356),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    LocalMux I__3178 (
            .O(N__15353),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    InMux I__3177 (
            .O(N__15344),
            .I(N__15341));
    LocalMux I__3176 (
            .O(N__15341),
            .I(N__15337));
    InMux I__3175 (
            .O(N__15340),
            .I(N__15334));
    Odrv4 I__3174 (
            .O(N__15337),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_3 ));
    LocalMux I__3173 (
            .O(N__15334),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_3 ));
    CEMux I__3172 (
            .O(N__15329),
            .I(N__15324));
    CEMux I__3171 (
            .O(N__15328),
            .I(N__15321));
    CEMux I__3170 (
            .O(N__15327),
            .I(N__15318));
    LocalMux I__3169 (
            .O(N__15324),
            .I(N__15313));
    LocalMux I__3168 (
            .O(N__15321),
            .I(N__15308));
    LocalMux I__3167 (
            .O(N__15318),
            .I(N__15308));
    CEMux I__3166 (
            .O(N__15317),
            .I(N__15303));
    CEMux I__3165 (
            .O(N__15316),
            .I(N__15300));
    Span4Mux_v I__3164 (
            .O(N__15313),
            .I(N__15296));
    Span4Mux_v I__3163 (
            .O(N__15308),
            .I(N__15293));
    CEMux I__3162 (
            .O(N__15307),
            .I(N__15289));
    CEMux I__3161 (
            .O(N__15306),
            .I(N__15286));
    LocalMux I__3160 (
            .O(N__15303),
            .I(N__15283));
    LocalMux I__3159 (
            .O(N__15300),
            .I(N__15280));
    CEMux I__3158 (
            .O(N__15299),
            .I(N__15277));
    Span4Mux_v I__3157 (
            .O(N__15296),
            .I(N__15272));
    Span4Mux_h I__3156 (
            .O(N__15293),
            .I(N__15272));
    CEMux I__3155 (
            .O(N__15292),
            .I(N__15269));
    LocalMux I__3154 (
            .O(N__15289),
            .I(N__15265));
    LocalMux I__3153 (
            .O(N__15286),
            .I(N__15262));
    Span4Mux_v I__3152 (
            .O(N__15283),
            .I(N__15259));
    Span4Mux_v I__3151 (
            .O(N__15280),
            .I(N__15256));
    LocalMux I__3150 (
            .O(N__15277),
            .I(N__15253));
    Span4Mux_h I__3149 (
            .O(N__15272),
            .I(N__15248));
    LocalMux I__3148 (
            .O(N__15269),
            .I(N__15248));
    CEMux I__3147 (
            .O(N__15268),
            .I(N__15245));
    Span4Mux_h I__3146 (
            .O(N__15265),
            .I(N__15242));
    Span4Mux_h I__3145 (
            .O(N__15262),
            .I(N__15239));
    Span4Mux_h I__3144 (
            .O(N__15259),
            .I(N__15232));
    Span4Mux_h I__3143 (
            .O(N__15256),
            .I(N__15232));
    Span4Mux_v I__3142 (
            .O(N__15253),
            .I(N__15232));
    Span4Mux_v I__3141 (
            .O(N__15248),
            .I(N__15227));
    LocalMux I__3140 (
            .O(N__15245),
            .I(N__15227));
    Odrv4 I__3139 (
            .O(N__15242),
            .I(\this_vga_signals.N_550_2 ));
    Odrv4 I__3138 (
            .O(N__15239),
            .I(\this_vga_signals.N_550_2 ));
    Odrv4 I__3137 (
            .O(N__15232),
            .I(\this_vga_signals.N_550_2 ));
    Odrv4 I__3136 (
            .O(N__15227),
            .I(\this_vga_signals.N_550_2 ));
    SRMux I__3135 (
            .O(N__15218),
            .I(N__15212));
    SRMux I__3134 (
            .O(N__15217),
            .I(N__15208));
    SRMux I__3133 (
            .O(N__15216),
            .I(N__15205));
    SRMux I__3132 (
            .O(N__15215),
            .I(N__15201));
    LocalMux I__3131 (
            .O(N__15212),
            .I(N__15198));
    SRMux I__3130 (
            .O(N__15211),
            .I(N__15194));
    LocalMux I__3129 (
            .O(N__15208),
            .I(N__15190));
    LocalMux I__3128 (
            .O(N__15205),
            .I(N__15187));
    SRMux I__3127 (
            .O(N__15204),
            .I(N__15184));
    LocalMux I__3126 (
            .O(N__15201),
            .I(N__15180));
    Span4Mux_v I__3125 (
            .O(N__15198),
            .I(N__15176));
    SRMux I__3124 (
            .O(N__15197),
            .I(N__15173));
    LocalMux I__3123 (
            .O(N__15194),
            .I(N__15170));
    SRMux I__3122 (
            .O(N__15193),
            .I(N__15167));
    Span4Mux_v I__3121 (
            .O(N__15190),
            .I(N__15162));
    Span4Mux_v I__3120 (
            .O(N__15187),
            .I(N__15162));
    LocalMux I__3119 (
            .O(N__15184),
            .I(N__15159));
    SRMux I__3118 (
            .O(N__15183),
            .I(N__15156));
    Span4Mux_h I__3117 (
            .O(N__15180),
            .I(N__15153));
    SRMux I__3116 (
            .O(N__15179),
            .I(N__15150));
    Span4Mux_h I__3115 (
            .O(N__15176),
            .I(N__15147));
    LocalMux I__3114 (
            .O(N__15173),
            .I(N__15144));
    Span4Mux_h I__3113 (
            .O(N__15170),
            .I(N__15139));
    LocalMux I__3112 (
            .O(N__15167),
            .I(N__15139));
    Span4Mux_v I__3111 (
            .O(N__15162),
            .I(N__15132));
    Span4Mux_v I__3110 (
            .O(N__15159),
            .I(N__15132));
    LocalMux I__3109 (
            .O(N__15156),
            .I(N__15132));
    Span4Mux_h I__3108 (
            .O(N__15153),
            .I(N__15127));
    LocalMux I__3107 (
            .O(N__15150),
            .I(N__15127));
    Span4Mux_h I__3106 (
            .O(N__15147),
            .I(N__15123));
    Span4Mux_v I__3105 (
            .O(N__15144),
            .I(N__15120));
    Span4Mux_h I__3104 (
            .O(N__15139),
            .I(N__15115));
    Span4Mux_h I__3103 (
            .O(N__15132),
            .I(N__15115));
    Sp12to4 I__3102 (
            .O(N__15127),
            .I(N__15112));
    InMux I__3101 (
            .O(N__15126),
            .I(N__15109));
    Odrv4 I__3100 (
            .O(N__15123),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9 ));
    Odrv4 I__3099 (
            .O(N__15120),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9 ));
    Odrv4 I__3098 (
            .O(N__15115),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9 ));
    Odrv12 I__3097 (
            .O(N__15112),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9 ));
    LocalMux I__3096 (
            .O(N__15109),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9 ));
    InMux I__3095 (
            .O(N__15098),
            .I(N__15094));
    InMux I__3094 (
            .O(N__15097),
            .I(N__15091));
    LocalMux I__3093 (
            .O(N__15094),
            .I(N__15088));
    LocalMux I__3092 (
            .O(N__15091),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    Odrv4 I__3091 (
            .O(N__15088),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    CascadeMux I__3090 (
            .O(N__15083),
            .I(N__15079));
    InMux I__3089 (
            .O(N__15082),
            .I(N__15074));
    InMux I__3088 (
            .O(N__15079),
            .I(N__15074));
    LocalMux I__3087 (
            .O(N__15074),
            .I(N__15064));
    InMux I__3086 (
            .O(N__15073),
            .I(N__15061));
    InMux I__3085 (
            .O(N__15072),
            .I(N__15052));
    InMux I__3084 (
            .O(N__15071),
            .I(N__15052));
    InMux I__3083 (
            .O(N__15070),
            .I(N__15052));
    InMux I__3082 (
            .O(N__15069),
            .I(N__15052));
    CascadeMux I__3081 (
            .O(N__15068),
            .I(N__15047));
    InMux I__3080 (
            .O(N__15067),
            .I(N__15044));
    Span4Mux_v I__3079 (
            .O(N__15064),
            .I(N__15037));
    LocalMux I__3078 (
            .O(N__15061),
            .I(N__15037));
    LocalMux I__3077 (
            .O(N__15052),
            .I(N__15037));
    CascadeMux I__3076 (
            .O(N__15051),
            .I(N__15034));
    InMux I__3075 (
            .O(N__15050),
            .I(N__15029));
    InMux I__3074 (
            .O(N__15047),
            .I(N__15029));
    LocalMux I__3073 (
            .O(N__15044),
            .I(N__15024));
    Span4Mux_v I__3072 (
            .O(N__15037),
            .I(N__15024));
    InMux I__3071 (
            .O(N__15034),
            .I(N__15021));
    LocalMux I__3070 (
            .O(N__15029),
            .I(N__15018));
    Odrv4 I__3069 (
            .O(N__15024),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__3068 (
            .O(N__15021),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv12 I__3067 (
            .O(N__15018),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    CEMux I__3066 (
            .O(N__15011),
            .I(N__15008));
    LocalMux I__3065 (
            .O(N__15008),
            .I(N__15004));
    CEMux I__3064 (
            .O(N__15007),
            .I(N__15000));
    Span4Mux_v I__3063 (
            .O(N__15004),
            .I(N__14997));
    CEMux I__3062 (
            .O(N__15003),
            .I(N__14994));
    LocalMux I__3061 (
            .O(N__15000),
            .I(N__14991));
    Span4Mux_h I__3060 (
            .O(N__14997),
            .I(N__14985));
    LocalMux I__3059 (
            .O(N__14994),
            .I(N__14985));
    Span4Mux_h I__3058 (
            .O(N__14991),
            .I(N__14982));
    CEMux I__3057 (
            .O(N__14990),
            .I(N__14979));
    Span4Mux_h I__3056 (
            .O(N__14985),
            .I(N__14976));
    Sp12to4 I__3055 (
            .O(N__14982),
            .I(N__14971));
    LocalMux I__3054 (
            .O(N__14979),
            .I(N__14971));
    Odrv4 I__3053 (
            .O(N__14976),
            .I(\this_vga_signals.N_550_0 ));
    Odrv12 I__3052 (
            .O(N__14971),
            .I(\this_vga_signals.N_550_0 ));
    SRMux I__3051 (
            .O(N__14966),
            .I(N__14962));
    SRMux I__3050 (
            .O(N__14965),
            .I(N__14959));
    LocalMux I__3049 (
            .O(N__14962),
            .I(N__14954));
    LocalMux I__3048 (
            .O(N__14959),
            .I(N__14951));
    SRMux I__3047 (
            .O(N__14958),
            .I(N__14948));
    SRMux I__3046 (
            .O(N__14957),
            .I(N__14945));
    Span4Mux_v I__3045 (
            .O(N__14954),
            .I(N__14942));
    Span4Mux_v I__3044 (
            .O(N__14951),
            .I(N__14937));
    LocalMux I__3043 (
            .O(N__14948),
            .I(N__14937));
    LocalMux I__3042 (
            .O(N__14945),
            .I(N__14933));
    Span4Mux_h I__3041 (
            .O(N__14942),
            .I(N__14928));
    Span4Mux_h I__3040 (
            .O(N__14937),
            .I(N__14925));
    SRMux I__3039 (
            .O(N__14936),
            .I(N__14922));
    Span4Mux_h I__3038 (
            .O(N__14933),
            .I(N__14919));
    SRMux I__3037 (
            .O(N__14932),
            .I(N__14916));
    InMux I__3036 (
            .O(N__14931),
            .I(N__14913));
    Odrv4 I__3035 (
            .O(N__14928),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9 ));
    Odrv4 I__3034 (
            .O(N__14925),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9 ));
    LocalMux I__3033 (
            .O(N__14922),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9 ));
    Odrv4 I__3032 (
            .O(N__14919),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9 ));
    LocalMux I__3031 (
            .O(N__14916),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9 ));
    LocalMux I__3030 (
            .O(N__14913),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9 ));
    CascadeMux I__3029 (
            .O(N__14900),
            .I(\this_start_data_delay.M_this_state_q_srsts_i_1_2_cascade_ ));
    CascadeMux I__3028 (
            .O(N__14897),
            .I(N__14894));
    InMux I__3027 (
            .O(N__14894),
            .I(N__14891));
    LocalMux I__3026 (
            .O(N__14891),
            .I(\this_start_data_delay.N_389_1 ));
    IoInMux I__3025 (
            .O(N__14888),
            .I(N__14885));
    LocalMux I__3024 (
            .O(N__14885),
            .I(N__14882));
    Span4Mux_s0_h I__3023 (
            .O(N__14882),
            .I(N__14879));
    Span4Mux_h I__3022 (
            .O(N__14879),
            .I(N__14875));
    InMux I__3021 (
            .O(N__14878),
            .I(N__14871));
    Sp12to4 I__3020 (
            .O(N__14875),
            .I(N__14868));
    InMux I__3019 (
            .O(N__14874),
            .I(N__14865));
    LocalMux I__3018 (
            .O(N__14871),
            .I(N__14862));
    Span12Mux_v I__3017 (
            .O(N__14868),
            .I(N__14858));
    LocalMux I__3016 (
            .O(N__14865),
            .I(N__14855));
    Span12Mux_v I__3015 (
            .O(N__14862),
            .I(N__14852));
    InMux I__3014 (
            .O(N__14861),
            .I(N__14849));
    Span12Mux_h I__3013 (
            .O(N__14858),
            .I(N__14846));
    Span12Mux_s7_h I__3012 (
            .O(N__14855),
            .I(N__14843));
    Span12Mux_h I__3011 (
            .O(N__14852),
            .I(N__14840));
    LocalMux I__3010 (
            .O(N__14849),
            .I(N__14837));
    Odrv12 I__3009 (
            .O(N__14846),
            .I(port_dmab_c));
    Odrv12 I__3008 (
            .O(N__14843),
            .I(port_dmab_c));
    Odrv12 I__3007 (
            .O(N__14840),
            .I(port_dmab_c));
    Odrv4 I__3006 (
            .O(N__14837),
            .I(port_dmab_c));
    CascadeMux I__3005 (
            .O(N__14828),
            .I(port_dmab_c_cascade_));
    CascadeMux I__3004 (
            .O(N__14825),
            .I(\this_start_data_delay.N_385_cascade_ ));
    InMux I__3003 (
            .O(N__14822),
            .I(bfn_16_25_0_));
    CascadeMux I__3002 (
            .O(N__14819),
            .I(\this_vga_signals.mult1_un54_sum_1_c2_1_cascade_ ));
    CascadeMux I__3001 (
            .O(N__14816),
            .I(N__14809));
    CascadeMux I__3000 (
            .O(N__14815),
            .I(N__14806));
    CascadeMux I__2999 (
            .O(N__14814),
            .I(N__14803));
    CascadeMux I__2998 (
            .O(N__14813),
            .I(N__14795));
    InMux I__2997 (
            .O(N__14812),
            .I(N__14792));
    InMux I__2996 (
            .O(N__14809),
            .I(N__14786));
    InMux I__2995 (
            .O(N__14806),
            .I(N__14783));
    InMux I__2994 (
            .O(N__14803),
            .I(N__14780));
    InMux I__2993 (
            .O(N__14802),
            .I(N__14777));
    InMux I__2992 (
            .O(N__14801),
            .I(N__14774));
    InMux I__2991 (
            .O(N__14800),
            .I(N__14771));
    InMux I__2990 (
            .O(N__14799),
            .I(N__14767));
    InMux I__2989 (
            .O(N__14798),
            .I(N__14762));
    InMux I__2988 (
            .O(N__14795),
            .I(N__14762));
    LocalMux I__2987 (
            .O(N__14792),
            .I(N__14759));
    InMux I__2986 (
            .O(N__14791),
            .I(N__14755));
    InMux I__2985 (
            .O(N__14790),
            .I(N__14747));
    InMux I__2984 (
            .O(N__14789),
            .I(N__14742));
    LocalMux I__2983 (
            .O(N__14786),
            .I(N__14735));
    LocalMux I__2982 (
            .O(N__14783),
            .I(N__14735));
    LocalMux I__2981 (
            .O(N__14780),
            .I(N__14726));
    LocalMux I__2980 (
            .O(N__14777),
            .I(N__14726));
    LocalMux I__2979 (
            .O(N__14774),
            .I(N__14726));
    LocalMux I__2978 (
            .O(N__14771),
            .I(N__14726));
    InMux I__2977 (
            .O(N__14770),
            .I(N__14723));
    LocalMux I__2976 (
            .O(N__14767),
            .I(N__14718));
    LocalMux I__2975 (
            .O(N__14762),
            .I(N__14718));
    Span4Mux_v I__2974 (
            .O(N__14759),
            .I(N__14714));
    InMux I__2973 (
            .O(N__14758),
            .I(N__14711));
    LocalMux I__2972 (
            .O(N__14755),
            .I(N__14708));
    InMux I__2971 (
            .O(N__14754),
            .I(N__14705));
    InMux I__2970 (
            .O(N__14753),
            .I(N__14700));
    InMux I__2969 (
            .O(N__14752),
            .I(N__14700));
    InMux I__2968 (
            .O(N__14751),
            .I(N__14695));
    InMux I__2967 (
            .O(N__14750),
            .I(N__14695));
    LocalMux I__2966 (
            .O(N__14747),
            .I(N__14692));
    InMux I__2965 (
            .O(N__14746),
            .I(N__14689));
    InMux I__2964 (
            .O(N__14745),
            .I(N__14686));
    LocalMux I__2963 (
            .O(N__14742),
            .I(N__14683));
    InMux I__2962 (
            .O(N__14741),
            .I(N__14680));
    InMux I__2961 (
            .O(N__14740),
            .I(N__14677));
    Span4Mux_v I__2960 (
            .O(N__14735),
            .I(N__14672));
    Span4Mux_v I__2959 (
            .O(N__14726),
            .I(N__14672));
    LocalMux I__2958 (
            .O(N__14723),
            .I(N__14667));
    Span4Mux_h I__2957 (
            .O(N__14718),
            .I(N__14667));
    InMux I__2956 (
            .O(N__14717),
            .I(N__14664));
    Span4Mux_h I__2955 (
            .O(N__14714),
            .I(N__14653));
    LocalMux I__2954 (
            .O(N__14711),
            .I(N__14653));
    Span4Mux_v I__2953 (
            .O(N__14708),
            .I(N__14653));
    LocalMux I__2952 (
            .O(N__14705),
            .I(N__14653));
    LocalMux I__2951 (
            .O(N__14700),
            .I(N__14653));
    LocalMux I__2950 (
            .O(N__14695),
            .I(N__14644));
    Span4Mux_h I__2949 (
            .O(N__14692),
            .I(N__14644));
    LocalMux I__2948 (
            .O(N__14689),
            .I(N__14644));
    LocalMux I__2947 (
            .O(N__14686),
            .I(N__14644));
    Odrv4 I__2946 (
            .O(N__14683),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2945 (
            .O(N__14680),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2944 (
            .O(N__14677),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__2943 (
            .O(N__14672),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__2942 (
            .O(N__14667),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2941 (
            .O(N__14664),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__2940 (
            .O(N__14653),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__2939 (
            .O(N__14644),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    InMux I__2938 (
            .O(N__14627),
            .I(N__14624));
    LocalMux I__2937 (
            .O(N__14624),
            .I(N__14621));
    Odrv4 I__2936 (
            .O(N__14621),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIUFPQ_2Z0Z_9 ));
    CascadeMux I__2935 (
            .O(N__14618),
            .I(\this_vga_signals.mult1_un54_sum_1_c2_cascade_ ));
    CascadeMux I__2934 (
            .O(N__14615),
            .I(N__14612));
    InMux I__2933 (
            .O(N__14612),
            .I(N__14603));
    InMux I__2932 (
            .O(N__14611),
            .I(N__14595));
    InMux I__2931 (
            .O(N__14610),
            .I(N__14595));
    InMux I__2930 (
            .O(N__14609),
            .I(N__14595));
    InMux I__2929 (
            .O(N__14608),
            .I(N__14592));
    CascadeMux I__2928 (
            .O(N__14607),
            .I(N__14588));
    InMux I__2927 (
            .O(N__14606),
            .I(N__14585));
    LocalMux I__2926 (
            .O(N__14603),
            .I(N__14582));
    InMux I__2925 (
            .O(N__14602),
            .I(N__14579));
    LocalMux I__2924 (
            .O(N__14595),
            .I(N__14572));
    LocalMux I__2923 (
            .O(N__14592),
            .I(N__14572));
    InMux I__2922 (
            .O(N__14591),
            .I(N__14569));
    InMux I__2921 (
            .O(N__14588),
            .I(N__14566));
    LocalMux I__2920 (
            .O(N__14585),
            .I(N__14561));
    Span4Mux_v I__2919 (
            .O(N__14582),
            .I(N__14556));
    LocalMux I__2918 (
            .O(N__14579),
            .I(N__14556));
    InMux I__2917 (
            .O(N__14578),
            .I(N__14553));
    InMux I__2916 (
            .O(N__14577),
            .I(N__14550));
    Span4Mux_h I__2915 (
            .O(N__14572),
            .I(N__14547));
    LocalMux I__2914 (
            .O(N__14569),
            .I(N__14542));
    LocalMux I__2913 (
            .O(N__14566),
            .I(N__14542));
    InMux I__2912 (
            .O(N__14565),
            .I(N__14539));
    InMux I__2911 (
            .O(N__14564),
            .I(N__14536));
    Span4Mux_h I__2910 (
            .O(N__14561),
            .I(N__14525));
    Span4Mux_h I__2909 (
            .O(N__14556),
            .I(N__14525));
    LocalMux I__2908 (
            .O(N__14553),
            .I(N__14520));
    LocalMux I__2907 (
            .O(N__14550),
            .I(N__14520));
    Span4Mux_h I__2906 (
            .O(N__14547),
            .I(N__14511));
    Span4Mux_h I__2905 (
            .O(N__14542),
            .I(N__14511));
    LocalMux I__2904 (
            .O(N__14539),
            .I(N__14511));
    LocalMux I__2903 (
            .O(N__14536),
            .I(N__14511));
    InMux I__2902 (
            .O(N__14535),
            .I(N__14506));
    InMux I__2901 (
            .O(N__14534),
            .I(N__14506));
    InMux I__2900 (
            .O(N__14533),
            .I(N__14501));
    InMux I__2899 (
            .O(N__14532),
            .I(N__14501));
    InMux I__2898 (
            .O(N__14531),
            .I(N__14496));
    InMux I__2897 (
            .O(N__14530),
            .I(N__14496));
    Odrv4 I__2896 (
            .O(N__14525),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv12 I__2895 (
            .O(N__14520),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__2894 (
            .O(N__14511),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__2893 (
            .O(N__14506),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__2892 (
            .O(N__14501),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__2891 (
            .O(N__14496),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    CascadeMux I__2890 (
            .O(N__14483),
            .I(N__14473));
    CascadeMux I__2889 (
            .O(N__14482),
            .I(N__14467));
    CascadeMux I__2888 (
            .O(N__14481),
            .I(N__14464));
    CascadeMux I__2887 (
            .O(N__14480),
            .I(N__14459));
    CascadeMux I__2886 (
            .O(N__14479),
            .I(N__14456));
    InMux I__2885 (
            .O(N__14478),
            .I(N__14453));
    InMux I__2884 (
            .O(N__14477),
            .I(N__14450));
    InMux I__2883 (
            .O(N__14476),
            .I(N__14444));
    InMux I__2882 (
            .O(N__14473),
            .I(N__14444));
    CascadeMux I__2881 (
            .O(N__14472),
            .I(N__14441));
    CascadeMux I__2880 (
            .O(N__14471),
            .I(N__14438));
    InMux I__2879 (
            .O(N__14470),
            .I(N__14434));
    InMux I__2878 (
            .O(N__14467),
            .I(N__14431));
    InMux I__2877 (
            .O(N__14464),
            .I(N__14428));
    InMux I__2876 (
            .O(N__14463),
            .I(N__14423));
    InMux I__2875 (
            .O(N__14462),
            .I(N__14423));
    InMux I__2874 (
            .O(N__14459),
            .I(N__14418));
    InMux I__2873 (
            .O(N__14456),
            .I(N__14418));
    LocalMux I__2872 (
            .O(N__14453),
            .I(N__14415));
    LocalMux I__2871 (
            .O(N__14450),
            .I(N__14412));
    CascadeMux I__2870 (
            .O(N__14449),
            .I(N__14409));
    LocalMux I__2869 (
            .O(N__14444),
            .I(N__14405));
    InMux I__2868 (
            .O(N__14441),
            .I(N__14402));
    InMux I__2867 (
            .O(N__14438),
            .I(N__14399));
    InMux I__2866 (
            .O(N__14437),
            .I(N__14394));
    LocalMux I__2865 (
            .O(N__14434),
            .I(N__14391));
    LocalMux I__2864 (
            .O(N__14431),
            .I(N__14388));
    LocalMux I__2863 (
            .O(N__14428),
            .I(N__14385));
    LocalMux I__2862 (
            .O(N__14423),
            .I(N__14380));
    LocalMux I__2861 (
            .O(N__14418),
            .I(N__14380));
    Span4Mux_v I__2860 (
            .O(N__14415),
            .I(N__14377));
    Span4Mux_v I__2859 (
            .O(N__14412),
            .I(N__14374));
    InMux I__2858 (
            .O(N__14409),
            .I(N__14371));
    InMux I__2857 (
            .O(N__14408),
            .I(N__14368));
    Span4Mux_v I__2856 (
            .O(N__14405),
            .I(N__14365));
    LocalMux I__2855 (
            .O(N__14402),
            .I(N__14362));
    LocalMux I__2854 (
            .O(N__14399),
            .I(N__14359));
    CascadeMux I__2853 (
            .O(N__14398),
            .I(N__14356));
    CascadeMux I__2852 (
            .O(N__14397),
            .I(N__14353));
    LocalMux I__2851 (
            .O(N__14394),
            .I(N__14348));
    Span4Mux_v I__2850 (
            .O(N__14391),
            .I(N__14348));
    Span4Mux_h I__2849 (
            .O(N__14388),
            .I(N__14341));
    Span4Mux_h I__2848 (
            .O(N__14385),
            .I(N__14341));
    Span4Mux_v I__2847 (
            .O(N__14380),
            .I(N__14341));
    Span4Mux_v I__2846 (
            .O(N__14377),
            .I(N__14336));
    Span4Mux_h I__2845 (
            .O(N__14374),
            .I(N__14336));
    LocalMux I__2844 (
            .O(N__14371),
            .I(N__14331));
    LocalMux I__2843 (
            .O(N__14368),
            .I(N__14331));
    Span4Mux_h I__2842 (
            .O(N__14365),
            .I(N__14324));
    Span4Mux_v I__2841 (
            .O(N__14362),
            .I(N__14324));
    Span4Mux_v I__2840 (
            .O(N__14359),
            .I(N__14324));
    InMux I__2839 (
            .O(N__14356),
            .I(N__14319));
    InMux I__2838 (
            .O(N__14353),
            .I(N__14319));
    Span4Mux_v I__2837 (
            .O(N__14348),
            .I(N__14314));
    Span4Mux_h I__2836 (
            .O(N__14341),
            .I(N__14314));
    Odrv4 I__2835 (
            .O(N__14336),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv12 I__2834 (
            .O(N__14331),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__2833 (
            .O(N__14324),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__2832 (
            .O(N__14319),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__2831 (
            .O(N__14314),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    CascadeMux I__2830 (
            .O(N__14303),
            .I(N__14299));
    InMux I__2829 (
            .O(N__14302),
            .I(N__14293));
    InMux I__2828 (
            .O(N__14299),
            .I(N__14287));
    InMux I__2827 (
            .O(N__14298),
            .I(N__14287));
    InMux I__2826 (
            .O(N__14297),
            .I(N__14284));
    InMux I__2825 (
            .O(N__14296),
            .I(N__14280));
    LocalMux I__2824 (
            .O(N__14293),
            .I(N__14275));
    InMux I__2823 (
            .O(N__14292),
            .I(N__14272));
    LocalMux I__2822 (
            .O(N__14287),
            .I(N__14268));
    LocalMux I__2821 (
            .O(N__14284),
            .I(N__14260));
    InMux I__2820 (
            .O(N__14283),
            .I(N__14255));
    LocalMux I__2819 (
            .O(N__14280),
            .I(N__14252));
    InMux I__2818 (
            .O(N__14279),
            .I(N__14249));
    InMux I__2817 (
            .O(N__14278),
            .I(N__14246));
    Span4Mux_v I__2816 (
            .O(N__14275),
            .I(N__14243));
    LocalMux I__2815 (
            .O(N__14272),
            .I(N__14240));
    InMux I__2814 (
            .O(N__14271),
            .I(N__14237));
    Span4Mux_v I__2813 (
            .O(N__14268),
            .I(N__14234));
    InMux I__2812 (
            .O(N__14267),
            .I(N__14231));
    InMux I__2811 (
            .O(N__14266),
            .I(N__14228));
    InMux I__2810 (
            .O(N__14265),
            .I(N__14225));
    InMux I__2809 (
            .O(N__14264),
            .I(N__14220));
    InMux I__2808 (
            .O(N__14263),
            .I(N__14220));
    Span4Mux_v I__2807 (
            .O(N__14260),
            .I(N__14216));
    InMux I__2806 (
            .O(N__14259),
            .I(N__14213));
    InMux I__2805 (
            .O(N__14258),
            .I(N__14210));
    LocalMux I__2804 (
            .O(N__14255),
            .I(N__14205));
    Span4Mux_v I__2803 (
            .O(N__14252),
            .I(N__14205));
    LocalMux I__2802 (
            .O(N__14249),
            .I(N__14200));
    LocalMux I__2801 (
            .O(N__14246),
            .I(N__14200));
    Span4Mux_h I__2800 (
            .O(N__14243),
            .I(N__14191));
    Span4Mux_h I__2799 (
            .O(N__14240),
            .I(N__14191));
    LocalMux I__2798 (
            .O(N__14237),
            .I(N__14191));
    Span4Mux_h I__2797 (
            .O(N__14234),
            .I(N__14182));
    LocalMux I__2796 (
            .O(N__14231),
            .I(N__14182));
    LocalMux I__2795 (
            .O(N__14228),
            .I(N__14182));
    LocalMux I__2794 (
            .O(N__14225),
            .I(N__14182));
    LocalMux I__2793 (
            .O(N__14220),
            .I(N__14179));
    CascadeMux I__2792 (
            .O(N__14219),
            .I(N__14174));
    Sp12to4 I__2791 (
            .O(N__14216),
            .I(N__14167));
    LocalMux I__2790 (
            .O(N__14213),
            .I(N__14167));
    LocalMux I__2789 (
            .O(N__14210),
            .I(N__14167));
    Span4Mux_v I__2788 (
            .O(N__14205),
            .I(N__14162));
    Span4Mux_v I__2787 (
            .O(N__14200),
            .I(N__14162));
    InMux I__2786 (
            .O(N__14199),
            .I(N__14157));
    InMux I__2785 (
            .O(N__14198),
            .I(N__14157));
    Span4Mux_v I__2784 (
            .O(N__14191),
            .I(N__14150));
    Span4Mux_v I__2783 (
            .O(N__14182),
            .I(N__14150));
    Span4Mux_h I__2782 (
            .O(N__14179),
            .I(N__14150));
    InMux I__2781 (
            .O(N__14178),
            .I(N__14147));
    InMux I__2780 (
            .O(N__14177),
            .I(N__14144));
    InMux I__2779 (
            .O(N__14174),
            .I(N__14141));
    Odrv12 I__2778 (
            .O(N__14167),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__2777 (
            .O(N__14162),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2776 (
            .O(N__14157),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__2775 (
            .O(N__14150),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2774 (
            .O(N__14147),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2773 (
            .O(N__14144),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2772 (
            .O(N__14141),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    CascadeMux I__2771 (
            .O(N__14126),
            .I(N__14123));
    InMux I__2770 (
            .O(N__14123),
            .I(N__14120));
    LocalMux I__2769 (
            .O(N__14120),
            .I(N__14108));
    InMux I__2768 (
            .O(N__14119),
            .I(N__14103));
    InMux I__2767 (
            .O(N__14118),
            .I(N__14103));
    InMux I__2766 (
            .O(N__14117),
            .I(N__14099));
    InMux I__2765 (
            .O(N__14116),
            .I(N__14094));
    InMux I__2764 (
            .O(N__14115),
            .I(N__14087));
    InMux I__2763 (
            .O(N__14114),
            .I(N__14087));
    InMux I__2762 (
            .O(N__14113),
            .I(N__14084));
    InMux I__2761 (
            .O(N__14112),
            .I(N__14081));
    InMux I__2760 (
            .O(N__14111),
            .I(N__14078));
    Span4Mux_v I__2759 (
            .O(N__14108),
            .I(N__14071));
    LocalMux I__2758 (
            .O(N__14103),
            .I(N__14071));
    InMux I__2757 (
            .O(N__14102),
            .I(N__14068));
    LocalMux I__2756 (
            .O(N__14099),
            .I(N__14065));
    InMux I__2755 (
            .O(N__14098),
            .I(N__14062));
    InMux I__2754 (
            .O(N__14097),
            .I(N__14059));
    LocalMux I__2753 (
            .O(N__14094),
            .I(N__14056));
    InMux I__2752 (
            .O(N__14093),
            .I(N__14053));
    InMux I__2751 (
            .O(N__14092),
            .I(N__14050));
    LocalMux I__2750 (
            .O(N__14087),
            .I(N__14045));
    LocalMux I__2749 (
            .O(N__14084),
            .I(N__14045));
    LocalMux I__2748 (
            .O(N__14081),
            .I(N__14040));
    LocalMux I__2747 (
            .O(N__14078),
            .I(N__14040));
    InMux I__2746 (
            .O(N__14077),
            .I(N__14035));
    InMux I__2745 (
            .O(N__14076),
            .I(N__14032));
    Span4Mux_h I__2744 (
            .O(N__14071),
            .I(N__14027));
    LocalMux I__2743 (
            .O(N__14068),
            .I(N__14027));
    Span4Mux_v I__2742 (
            .O(N__14065),
            .I(N__14020));
    LocalMux I__2741 (
            .O(N__14062),
            .I(N__14020));
    LocalMux I__2740 (
            .O(N__14059),
            .I(N__14020));
    Span4Mux_v I__2739 (
            .O(N__14056),
            .I(N__14015));
    LocalMux I__2738 (
            .O(N__14053),
            .I(N__14015));
    LocalMux I__2737 (
            .O(N__14050),
            .I(N__14012));
    Span4Mux_v I__2736 (
            .O(N__14045),
            .I(N__14007));
    Span4Mux_v I__2735 (
            .O(N__14040),
            .I(N__14007));
    InMux I__2734 (
            .O(N__14039),
            .I(N__14002));
    InMux I__2733 (
            .O(N__14038),
            .I(N__14002));
    LocalMux I__2732 (
            .O(N__14035),
            .I(N__13994));
    LocalMux I__2731 (
            .O(N__14032),
            .I(N__13994));
    Span4Mux_h I__2730 (
            .O(N__14027),
            .I(N__13985));
    Span4Mux_v I__2729 (
            .O(N__14020),
            .I(N__13985));
    Span4Mux_v I__2728 (
            .O(N__14015),
            .I(N__13985));
    Span4Mux_v I__2727 (
            .O(N__14012),
            .I(N__13985));
    Span4Mux_h I__2726 (
            .O(N__14007),
            .I(N__13980));
    LocalMux I__2725 (
            .O(N__14002),
            .I(N__13980));
    InMux I__2724 (
            .O(N__14001),
            .I(N__13975));
    InMux I__2723 (
            .O(N__14000),
            .I(N__13975));
    InMux I__2722 (
            .O(N__13999),
            .I(N__13972));
    Odrv12 I__2721 (
            .O(N__13994),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__2720 (
            .O(N__13985),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__2719 (
            .O(N__13980),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__2718 (
            .O(N__13975),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__2717 (
            .O(N__13972),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    InMux I__2716 (
            .O(N__13961),
            .I(N__13958));
    LocalMux I__2715 (
            .O(N__13958),
            .I(\this_vga_signals.mult1_un54_sum1_i_1_3 ));
    CascadeMux I__2714 (
            .O(N__13955),
            .I(N__13952));
    CascadeBuf I__2713 (
            .O(N__13952),
            .I(N__13949));
    CascadeMux I__2712 (
            .O(N__13949),
            .I(N__13946));
    CascadeBuf I__2711 (
            .O(N__13946),
            .I(N__13943));
    CascadeMux I__2710 (
            .O(N__13943),
            .I(N__13940));
    CascadeBuf I__2709 (
            .O(N__13940),
            .I(N__13937));
    CascadeMux I__2708 (
            .O(N__13937),
            .I(N__13934));
    CascadeBuf I__2707 (
            .O(N__13934),
            .I(N__13931));
    CascadeMux I__2706 (
            .O(N__13931),
            .I(N__13928));
    CascadeBuf I__2705 (
            .O(N__13928),
            .I(N__13925));
    CascadeMux I__2704 (
            .O(N__13925),
            .I(N__13922));
    CascadeBuf I__2703 (
            .O(N__13922),
            .I(N__13919));
    CascadeMux I__2702 (
            .O(N__13919),
            .I(N__13916));
    CascadeBuf I__2701 (
            .O(N__13916),
            .I(N__13913));
    CascadeMux I__2700 (
            .O(N__13913),
            .I(N__13910));
    CascadeBuf I__2699 (
            .O(N__13910),
            .I(N__13907));
    CascadeMux I__2698 (
            .O(N__13907),
            .I(N__13904));
    CascadeBuf I__2697 (
            .O(N__13904),
            .I(N__13901));
    CascadeMux I__2696 (
            .O(N__13901),
            .I(N__13898));
    CascadeBuf I__2695 (
            .O(N__13898),
            .I(N__13895));
    CascadeMux I__2694 (
            .O(N__13895),
            .I(N__13892));
    CascadeBuf I__2693 (
            .O(N__13892),
            .I(N__13889));
    CascadeMux I__2692 (
            .O(N__13889),
            .I(N__13886));
    CascadeBuf I__2691 (
            .O(N__13886),
            .I(N__13883));
    CascadeMux I__2690 (
            .O(N__13883),
            .I(N__13880));
    CascadeBuf I__2689 (
            .O(N__13880),
            .I(N__13877));
    CascadeMux I__2688 (
            .O(N__13877),
            .I(N__13874));
    CascadeBuf I__2687 (
            .O(N__13874),
            .I(N__13871));
    CascadeMux I__2686 (
            .O(N__13871),
            .I(N__13868));
    CascadeBuf I__2685 (
            .O(N__13868),
            .I(N__13865));
    CascadeMux I__2684 (
            .O(N__13865),
            .I(N__13862));
    InMux I__2683 (
            .O(N__13862),
            .I(N__13859));
    LocalMux I__2682 (
            .O(N__13859),
            .I(N__13856));
    Span12Mux_h I__2681 (
            .O(N__13856),
            .I(N__13853));
    Span12Mux_v I__2680 (
            .O(N__13853),
            .I(N__13850));
    Odrv12 I__2679 (
            .O(N__13850),
            .I(M_this_vga_signals_address_5));
    InMux I__2678 (
            .O(N__13847),
            .I(un1_M_this_data_count_q_cry_2));
    InMux I__2677 (
            .O(N__13844),
            .I(un1_M_this_data_count_q_cry_3));
    InMux I__2676 (
            .O(N__13841),
            .I(un1_M_this_data_count_q_cry_4));
    InMux I__2675 (
            .O(N__13838),
            .I(un1_M_this_data_count_q_cry_5));
    InMux I__2674 (
            .O(N__13835),
            .I(un1_M_this_data_count_q_cry_6));
    InMux I__2673 (
            .O(N__13832),
            .I(bfn_16_24_0_));
    InMux I__2672 (
            .O(N__13829),
            .I(un1_M_this_data_count_q_cry_8));
    InMux I__2671 (
            .O(N__13826),
            .I(un1_M_this_data_count_q_cry_9));
    InMux I__2670 (
            .O(N__13823),
            .I(un1_M_this_data_count_q_cry_10));
    InMux I__2669 (
            .O(N__13820),
            .I(un1_M_this_data_count_q_cry_11));
    InMux I__2668 (
            .O(N__13817),
            .I(N__13814));
    LocalMux I__2667 (
            .O(N__13814),
            .I(N__13811));
    Odrv4 I__2666 (
            .O(N__13811),
            .I(\this_vga_signals.vaddress_8 ));
    CascadeMux I__2665 (
            .O(N__13808),
            .I(N__13800));
    InMux I__2664 (
            .O(N__13807),
            .I(N__13791));
    InMux I__2663 (
            .O(N__13806),
            .I(N__13785));
    InMux I__2662 (
            .O(N__13805),
            .I(N__13785));
    InMux I__2661 (
            .O(N__13804),
            .I(N__13776));
    InMux I__2660 (
            .O(N__13803),
            .I(N__13776));
    InMux I__2659 (
            .O(N__13800),
            .I(N__13776));
    InMux I__2658 (
            .O(N__13799),
            .I(N__13776));
    InMux I__2657 (
            .O(N__13798),
            .I(N__13773));
    InMux I__2656 (
            .O(N__13797),
            .I(N__13768));
    InMux I__2655 (
            .O(N__13796),
            .I(N__13768));
    InMux I__2654 (
            .O(N__13795),
            .I(N__13763));
    InMux I__2653 (
            .O(N__13794),
            .I(N__13763));
    LocalMux I__2652 (
            .O(N__13791),
            .I(N__13760));
    InMux I__2651 (
            .O(N__13790),
            .I(N__13757));
    LocalMux I__2650 (
            .O(N__13785),
            .I(N__13752));
    LocalMux I__2649 (
            .O(N__13776),
            .I(N__13752));
    LocalMux I__2648 (
            .O(N__13773),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2647 (
            .O(N__13768),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2646 (
            .O(N__13763),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2645 (
            .O(N__13760),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2644 (
            .O(N__13757),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2643 (
            .O(N__13752),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    InMux I__2642 (
            .O(N__13739),
            .I(N__13735));
    CascadeMux I__2641 (
            .O(N__13738),
            .I(N__13732));
    LocalMux I__2640 (
            .O(N__13735),
            .I(N__13729));
    InMux I__2639 (
            .O(N__13732),
            .I(N__13724));
    Span4Mux_v I__2638 (
            .O(N__13729),
            .I(N__13712));
    InMux I__2637 (
            .O(N__13728),
            .I(N__13709));
    InMux I__2636 (
            .O(N__13727),
            .I(N__13706));
    LocalMux I__2635 (
            .O(N__13724),
            .I(N__13703));
    InMux I__2634 (
            .O(N__13723),
            .I(N__13696));
    InMux I__2633 (
            .O(N__13722),
            .I(N__13696));
    InMux I__2632 (
            .O(N__13721),
            .I(N__13696));
    InMux I__2631 (
            .O(N__13720),
            .I(N__13693));
    InMux I__2630 (
            .O(N__13719),
            .I(N__13684));
    InMux I__2629 (
            .O(N__13718),
            .I(N__13684));
    InMux I__2628 (
            .O(N__13717),
            .I(N__13684));
    InMux I__2627 (
            .O(N__13716),
            .I(N__13684));
    InMux I__2626 (
            .O(N__13715),
            .I(N__13681));
    Odrv4 I__2625 (
            .O(N__13712),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2624 (
            .O(N__13709),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2623 (
            .O(N__13706),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__2622 (
            .O(N__13703),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2621 (
            .O(N__13696),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2620 (
            .O(N__13693),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2619 (
            .O(N__13684),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2618 (
            .O(N__13681),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    InMux I__2617 (
            .O(N__13664),
            .I(N__13661));
    LocalMux I__2616 (
            .O(N__13661),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a2_x1 ));
    IoInMux I__2615 (
            .O(N__13658),
            .I(N__13655));
    LocalMux I__2614 (
            .O(N__13655),
            .I(N__13651));
    IoInMux I__2613 (
            .O(N__13654),
            .I(N__13648));
    IoSpan4Mux I__2612 (
            .O(N__13651),
            .I(N__13642));
    LocalMux I__2611 (
            .O(N__13648),
            .I(N__13642));
    IoInMux I__2610 (
            .O(N__13647),
            .I(N__13637));
    IoSpan4Mux I__2609 (
            .O(N__13642),
            .I(N__13632));
    IoInMux I__2608 (
            .O(N__13641),
            .I(N__13629));
    IoInMux I__2607 (
            .O(N__13640),
            .I(N__13626));
    LocalMux I__2606 (
            .O(N__13637),
            .I(N__13620));
    IoInMux I__2605 (
            .O(N__13636),
            .I(N__13617));
    IoInMux I__2604 (
            .O(N__13635),
            .I(N__13612));
    IoSpan4Mux I__2603 (
            .O(N__13632),
            .I(N__13607));
    LocalMux I__2602 (
            .O(N__13629),
            .I(N__13607));
    LocalMux I__2601 (
            .O(N__13626),
            .I(N__13604));
    IoInMux I__2600 (
            .O(N__13625),
            .I(N__13601));
    IoInMux I__2599 (
            .O(N__13624),
            .I(N__13598));
    IoInMux I__2598 (
            .O(N__13623),
            .I(N__13595));
    IoSpan4Mux I__2597 (
            .O(N__13620),
            .I(N__13587));
    LocalMux I__2596 (
            .O(N__13617),
            .I(N__13587));
    IoInMux I__2595 (
            .O(N__13616),
            .I(N__13584));
    IoInMux I__2594 (
            .O(N__13615),
            .I(N__13581));
    LocalMux I__2593 (
            .O(N__13612),
            .I(N__13577));
    IoSpan4Mux I__2592 (
            .O(N__13607),
            .I(N__13574));
    IoSpan4Mux I__2591 (
            .O(N__13604),
            .I(N__13567));
    LocalMux I__2590 (
            .O(N__13601),
            .I(N__13567));
    LocalMux I__2589 (
            .O(N__13598),
            .I(N__13567));
    LocalMux I__2588 (
            .O(N__13595),
            .I(N__13564));
    IoInMux I__2587 (
            .O(N__13594),
            .I(N__13561));
    IoInMux I__2586 (
            .O(N__13593),
            .I(N__13558));
    IoInMux I__2585 (
            .O(N__13592),
            .I(N__13555));
    IoSpan4Mux I__2584 (
            .O(N__13587),
            .I(N__13550));
    LocalMux I__2583 (
            .O(N__13584),
            .I(N__13550));
    LocalMux I__2582 (
            .O(N__13581),
            .I(N__13547));
    IoInMux I__2581 (
            .O(N__13580),
            .I(N__13544));
    Span4Mux_s3_v I__2580 (
            .O(N__13577),
            .I(N__13541));
    IoSpan4Mux I__2579 (
            .O(N__13574),
            .I(N__13536));
    IoSpan4Mux I__2578 (
            .O(N__13567),
            .I(N__13536));
    Span4Mux_s3_h I__2577 (
            .O(N__13564),
            .I(N__13533));
    LocalMux I__2576 (
            .O(N__13561),
            .I(N__13530));
    LocalMux I__2575 (
            .O(N__13558),
            .I(N__13527));
    LocalMux I__2574 (
            .O(N__13555),
            .I(N__13524));
    IoSpan4Mux I__2573 (
            .O(N__13550),
            .I(N__13517));
    IoSpan4Mux I__2572 (
            .O(N__13547),
            .I(N__13517));
    LocalMux I__2571 (
            .O(N__13544),
            .I(N__13517));
    Span4Mux_v I__2570 (
            .O(N__13541),
            .I(N__13514));
    Span4Mux_s3_h I__2569 (
            .O(N__13536),
            .I(N__13511));
    Span4Mux_v I__2568 (
            .O(N__13533),
            .I(N__13504));
    Span4Mux_s3_h I__2567 (
            .O(N__13530),
            .I(N__13504));
    Span4Mux_s3_h I__2566 (
            .O(N__13527),
            .I(N__13504));
    Span4Mux_s3_h I__2565 (
            .O(N__13524),
            .I(N__13501));
    IoSpan4Mux I__2564 (
            .O(N__13517),
            .I(N__13498));
    Span4Mux_v I__2563 (
            .O(N__13514),
            .I(N__13490));
    Span4Mux_h I__2562 (
            .O(N__13511),
            .I(N__13490));
    Span4Mux_h I__2561 (
            .O(N__13504),
            .I(N__13490));
    Span4Mux_h I__2560 (
            .O(N__13501),
            .I(N__13487));
    Span4Mux_s0_v I__2559 (
            .O(N__13498),
            .I(N__13484));
    IoInMux I__2558 (
            .O(N__13497),
            .I(N__13481));
    Span4Mux_h I__2557 (
            .O(N__13490),
            .I(N__13478));
    Span4Mux_h I__2556 (
            .O(N__13487),
            .I(N__13475));
    Sp12to4 I__2555 (
            .O(N__13484),
            .I(N__13470));
    LocalMux I__2554 (
            .O(N__13481),
            .I(N__13470));
    Span4Mux_h I__2553 (
            .O(N__13478),
            .I(N__13467));
    Span4Mux_h I__2552 (
            .O(N__13475),
            .I(N__13464));
    Span12Mux_s6_v I__2551 (
            .O(N__13470),
            .I(N__13461));
    Odrv4 I__2550 (
            .O(N__13467),
            .I(port_dmab_c_i));
    Odrv4 I__2549 (
            .O(N__13464),
            .I(port_dmab_c_i));
    Odrv12 I__2548 (
            .O(N__13461),
            .I(port_dmab_c_i));
    InMux I__2547 (
            .O(N__13454),
            .I(N__13449));
    InMux I__2546 (
            .O(N__13453),
            .I(N__13446));
    InMux I__2545 (
            .O(N__13452),
            .I(N__13442));
    LocalMux I__2544 (
            .O(N__13449),
            .I(N__13439));
    LocalMux I__2543 (
            .O(N__13446),
            .I(N__13435));
    InMux I__2542 (
            .O(N__13445),
            .I(N__13432));
    LocalMux I__2541 (
            .O(N__13442),
            .I(N__13429));
    Span4Mux_v I__2540 (
            .O(N__13439),
            .I(N__13419));
    InMux I__2539 (
            .O(N__13438),
            .I(N__13416));
    Span4Mux_h I__2538 (
            .O(N__13435),
            .I(N__13413));
    LocalMux I__2537 (
            .O(N__13432),
            .I(N__13410));
    Span4Mux_h I__2536 (
            .O(N__13429),
            .I(N__13407));
    InMux I__2535 (
            .O(N__13428),
            .I(N__13402));
    InMux I__2534 (
            .O(N__13427),
            .I(N__13402));
    InMux I__2533 (
            .O(N__13426),
            .I(N__13397));
    InMux I__2532 (
            .O(N__13425),
            .I(N__13397));
    InMux I__2531 (
            .O(N__13424),
            .I(N__13392));
    InMux I__2530 (
            .O(N__13423),
            .I(N__13392));
    InMux I__2529 (
            .O(N__13422),
            .I(N__13389));
    Odrv4 I__2528 (
            .O(N__13419),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2527 (
            .O(N__13416),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2526 (
            .O(N__13413),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2525 (
            .O(N__13410),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2524 (
            .O(N__13407),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2523 (
            .O(N__13402),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2522 (
            .O(N__13397),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2521 (
            .O(N__13392),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2520 (
            .O(N__13389),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    InMux I__2519 (
            .O(N__13370),
            .I(N__13367));
    LocalMux I__2518 (
            .O(N__13367),
            .I(N__13363));
    InMux I__2517 (
            .O(N__13366),
            .I(N__13360));
    Odrv4 I__2516 (
            .O(N__13363),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    LocalMux I__2515 (
            .O(N__13360),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    InMux I__2514 (
            .O(N__13355),
            .I(N__13349));
    InMux I__2513 (
            .O(N__13354),
            .I(N__13349));
    LocalMux I__2512 (
            .O(N__13349),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    InMux I__2511 (
            .O(N__13346),
            .I(un1_M_this_data_count_q_cry_0));
    InMux I__2510 (
            .O(N__13343),
            .I(un1_M_this_data_count_q_cry_1));
    InMux I__2509 (
            .O(N__13340),
            .I(bfn_15_22_0_));
    InMux I__2508 (
            .O(N__13337),
            .I(N__13326));
    InMux I__2507 (
            .O(N__13336),
            .I(N__13321));
    InMux I__2506 (
            .O(N__13335),
            .I(N__13321));
    InMux I__2505 (
            .O(N__13334),
            .I(N__13314));
    InMux I__2504 (
            .O(N__13333),
            .I(N__13314));
    InMux I__2503 (
            .O(N__13332),
            .I(N__13314));
    InMux I__2502 (
            .O(N__13331),
            .I(N__13311));
    InMux I__2501 (
            .O(N__13330),
            .I(N__13306));
    InMux I__2500 (
            .O(N__13329),
            .I(N__13306));
    LocalMux I__2499 (
            .O(N__13326),
            .I(N__13301));
    LocalMux I__2498 (
            .O(N__13321),
            .I(N__13301));
    LocalMux I__2497 (
            .O(N__13314),
            .I(N__13298));
    LocalMux I__2496 (
            .O(N__13311),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__2495 (
            .O(N__13306),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__2494 (
            .O(N__13301),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv12 I__2493 (
            .O(N__13298),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    CascadeMux I__2492 (
            .O(N__13289),
            .I(N__13286));
    InMux I__2491 (
            .O(N__13286),
            .I(N__13283));
    LocalMux I__2490 (
            .O(N__13283),
            .I(N__13278));
    InMux I__2489 (
            .O(N__13282),
            .I(N__13275));
    InMux I__2488 (
            .O(N__13281),
            .I(N__13272));
    Span4Mux_v I__2487 (
            .O(N__13278),
            .I(N__13269));
    LocalMux I__2486 (
            .O(N__13275),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    LocalMux I__2485 (
            .O(N__13272),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    Odrv4 I__2484 (
            .O(N__13269),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    InMux I__2483 (
            .O(N__13262),
            .I(N__13259));
    LocalMux I__2482 (
            .O(N__13259),
            .I(N__13255));
    InMux I__2481 (
            .O(N__13258),
            .I(N__13252));
    Span4Mux_h I__2480 (
            .O(N__13255),
            .I(N__13249));
    LocalMux I__2479 (
            .O(N__13252),
            .I(N__13246));
    Odrv4 I__2478 (
            .O(N__13249),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0 ));
    Odrv4 I__2477 (
            .O(N__13246),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_0 ));
    CascadeMux I__2476 (
            .O(N__13241),
            .I(N__13238));
    InMux I__2475 (
            .O(N__13238),
            .I(N__13235));
    LocalMux I__2474 (
            .O(N__13235),
            .I(N__13232));
    Odrv4 I__2473 (
            .O(N__13232),
            .I(\this_vga_signals.mult1_un54_sum_c2 ));
    InMux I__2472 (
            .O(N__13229),
            .I(N__13226));
    LocalMux I__2471 (
            .O(N__13226),
            .I(N__13223));
    Span4Mux_h I__2470 (
            .O(N__13223),
            .I(N__13217));
    InMux I__2469 (
            .O(N__13222),
            .I(N__13214));
    InMux I__2468 (
            .O(N__13221),
            .I(N__13209));
    InMux I__2467 (
            .O(N__13220),
            .I(N__13209));
    Odrv4 I__2466 (
            .O(N__13217),
            .I(\this_vga_signals.mult1_un47_sum_i_3 ));
    LocalMux I__2465 (
            .O(N__13214),
            .I(\this_vga_signals.mult1_un47_sum_i_3 ));
    LocalMux I__2464 (
            .O(N__13209),
            .I(\this_vga_signals.mult1_un47_sum_i_3 ));
    InMux I__2463 (
            .O(N__13202),
            .I(N__13185));
    InMux I__2462 (
            .O(N__13201),
            .I(N__13185));
    InMux I__2461 (
            .O(N__13200),
            .I(N__13185));
    InMux I__2460 (
            .O(N__13199),
            .I(N__13182));
    InMux I__2459 (
            .O(N__13198),
            .I(N__13178));
    InMux I__2458 (
            .O(N__13197),
            .I(N__13173));
    InMux I__2457 (
            .O(N__13196),
            .I(N__13173));
    InMux I__2456 (
            .O(N__13195),
            .I(N__13168));
    InMux I__2455 (
            .O(N__13194),
            .I(N__13168));
    InMux I__2454 (
            .O(N__13193),
            .I(N__13165));
    InMux I__2453 (
            .O(N__13192),
            .I(N__13162));
    LocalMux I__2452 (
            .O(N__13185),
            .I(N__13157));
    LocalMux I__2451 (
            .O(N__13182),
            .I(N__13157));
    InMux I__2450 (
            .O(N__13181),
            .I(N__13154));
    LocalMux I__2449 (
            .O(N__13178),
            .I(N__13151));
    LocalMux I__2448 (
            .O(N__13173),
            .I(N__13148));
    LocalMux I__2447 (
            .O(N__13168),
            .I(N__13145));
    LocalMux I__2446 (
            .O(N__13165),
            .I(N__13138));
    LocalMux I__2445 (
            .O(N__13162),
            .I(N__13138));
    Span4Mux_v I__2444 (
            .O(N__13157),
            .I(N__13138));
    LocalMux I__2443 (
            .O(N__13154),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv12 I__2442 (
            .O(N__13151),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__2441 (
            .O(N__13148),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__2440 (
            .O(N__13145),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__2439 (
            .O(N__13138),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    InMux I__2438 (
            .O(N__13127),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_1 ));
    CascadeMux I__2437 (
            .O(N__13124),
            .I(N__13117));
    CascadeMux I__2436 (
            .O(N__13123),
            .I(N__13110));
    CascadeMux I__2435 (
            .O(N__13122),
            .I(N__13107));
    InMux I__2434 (
            .O(N__13121),
            .I(N__13104));
    InMux I__2433 (
            .O(N__13120),
            .I(N__13101));
    InMux I__2432 (
            .O(N__13117),
            .I(N__13098));
    InMux I__2431 (
            .O(N__13116),
            .I(N__13093));
    InMux I__2430 (
            .O(N__13115),
            .I(N__13093));
    InMux I__2429 (
            .O(N__13114),
            .I(N__13090));
    InMux I__2428 (
            .O(N__13113),
            .I(N__13087));
    InMux I__2427 (
            .O(N__13110),
            .I(N__13081));
    InMux I__2426 (
            .O(N__13107),
            .I(N__13081));
    LocalMux I__2425 (
            .O(N__13104),
            .I(N__13077));
    LocalMux I__2424 (
            .O(N__13101),
            .I(N__13068));
    LocalMux I__2423 (
            .O(N__13098),
            .I(N__13068));
    LocalMux I__2422 (
            .O(N__13093),
            .I(N__13068));
    LocalMux I__2421 (
            .O(N__13090),
            .I(N__13068));
    LocalMux I__2420 (
            .O(N__13087),
            .I(N__13065));
    InMux I__2419 (
            .O(N__13086),
            .I(N__13062));
    LocalMux I__2418 (
            .O(N__13081),
            .I(N__13059));
    InMux I__2417 (
            .O(N__13080),
            .I(N__13056));
    Span4Mux_h I__2416 (
            .O(N__13077),
            .I(N__13051));
    Span4Mux_v I__2415 (
            .O(N__13068),
            .I(N__13051));
    Odrv4 I__2414 (
            .O(N__13065),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2413 (
            .O(N__13062),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2412 (
            .O(N__13059),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2411 (
            .O(N__13056),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2410 (
            .O(N__13051),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    InMux I__2409 (
            .O(N__13040),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_2 ));
    CascadeMux I__2408 (
            .O(N__13037),
            .I(N__13029));
    InMux I__2407 (
            .O(N__13036),
            .I(N__13022));
    CascadeMux I__2406 (
            .O(N__13035),
            .I(N__13014));
    CascadeMux I__2405 (
            .O(N__13034),
            .I(N__13011));
    InMux I__2404 (
            .O(N__13033),
            .I(N__13007));
    InMux I__2403 (
            .O(N__13032),
            .I(N__12996));
    InMux I__2402 (
            .O(N__13029),
            .I(N__12996));
    InMux I__2401 (
            .O(N__13028),
            .I(N__12996));
    InMux I__2400 (
            .O(N__13027),
            .I(N__12996));
    InMux I__2399 (
            .O(N__13026),
            .I(N__12996));
    InMux I__2398 (
            .O(N__13025),
            .I(N__12993));
    LocalMux I__2397 (
            .O(N__13022),
            .I(N__12990));
    InMux I__2396 (
            .O(N__13021),
            .I(N__12987));
    InMux I__2395 (
            .O(N__13020),
            .I(N__12984));
    InMux I__2394 (
            .O(N__13019),
            .I(N__12981));
    InMux I__2393 (
            .O(N__13018),
            .I(N__12976));
    InMux I__2392 (
            .O(N__13017),
            .I(N__12976));
    InMux I__2391 (
            .O(N__13014),
            .I(N__12971));
    InMux I__2390 (
            .O(N__13011),
            .I(N__12971));
    InMux I__2389 (
            .O(N__13010),
            .I(N__12968));
    LocalMux I__2388 (
            .O(N__13007),
            .I(N__12963));
    LocalMux I__2387 (
            .O(N__12996),
            .I(N__12963));
    LocalMux I__2386 (
            .O(N__12993),
            .I(N__12956));
    Span4Mux_h I__2385 (
            .O(N__12990),
            .I(N__12956));
    LocalMux I__2384 (
            .O(N__12987),
            .I(N__12956));
    LocalMux I__2383 (
            .O(N__12984),
            .I(N__12947));
    LocalMux I__2382 (
            .O(N__12981),
            .I(N__12947));
    LocalMux I__2381 (
            .O(N__12976),
            .I(N__12947));
    LocalMux I__2380 (
            .O(N__12971),
            .I(N__12947));
    LocalMux I__2379 (
            .O(N__12968),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv12 I__2378 (
            .O(N__12963),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2377 (
            .O(N__12956),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2376 (
            .O(N__12947),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    InMux I__2375 (
            .O(N__12938),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3 ));
    InMux I__2374 (
            .O(N__12935),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4 ));
    InMux I__2373 (
            .O(N__12932),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5 ));
    InMux I__2372 (
            .O(N__12929),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6 ));
    InMux I__2371 (
            .O(N__12926),
            .I(N__12907));
    InMux I__2370 (
            .O(N__12925),
            .I(N__12907));
    InMux I__2369 (
            .O(N__12924),
            .I(N__12907));
    InMux I__2368 (
            .O(N__12923),
            .I(N__12907));
    InMux I__2367 (
            .O(N__12922),
            .I(N__12902));
    InMux I__2366 (
            .O(N__12921),
            .I(N__12902));
    InMux I__2365 (
            .O(N__12920),
            .I(N__12897));
    InMux I__2364 (
            .O(N__12919),
            .I(N__12897));
    InMux I__2363 (
            .O(N__12918),
            .I(N__12892));
    InMux I__2362 (
            .O(N__12917),
            .I(N__12889));
    InMux I__2361 (
            .O(N__12916),
            .I(N__12886));
    LocalMux I__2360 (
            .O(N__12907),
            .I(N__12876));
    LocalMux I__2359 (
            .O(N__12902),
            .I(N__12876));
    LocalMux I__2358 (
            .O(N__12897),
            .I(N__12876));
    InMux I__2357 (
            .O(N__12896),
            .I(N__12873));
    InMux I__2356 (
            .O(N__12895),
            .I(N__12870));
    LocalMux I__2355 (
            .O(N__12892),
            .I(N__12865));
    LocalMux I__2354 (
            .O(N__12889),
            .I(N__12865));
    LocalMux I__2353 (
            .O(N__12886),
            .I(N__12862));
    InMux I__2352 (
            .O(N__12885),
            .I(N__12857));
    InMux I__2351 (
            .O(N__12884),
            .I(N__12857));
    CascadeMux I__2350 (
            .O(N__12883),
            .I(N__12854));
    Span4Mux_h I__2349 (
            .O(N__12876),
            .I(N__12850));
    LocalMux I__2348 (
            .O(N__12873),
            .I(N__12847));
    LocalMux I__2347 (
            .O(N__12870),
            .I(N__12844));
    Span4Mux_h I__2346 (
            .O(N__12865),
            .I(N__12837));
    Span4Mux_v I__2345 (
            .O(N__12862),
            .I(N__12837));
    LocalMux I__2344 (
            .O(N__12857),
            .I(N__12837));
    InMux I__2343 (
            .O(N__12854),
            .I(N__12832));
    InMux I__2342 (
            .O(N__12853),
            .I(N__12832));
    Span4Mux_h I__2341 (
            .O(N__12850),
            .I(N__12829));
    Span12Mux_v I__2340 (
            .O(N__12847),
            .I(N__12826));
    Span4Mux_v I__2339 (
            .O(N__12844),
            .I(N__12821));
    Span4Mux_h I__2338 (
            .O(N__12837),
            .I(N__12821));
    LocalMux I__2337 (
            .O(N__12832),
            .I(\this_vga_signals.GZ0Z_296 ));
    Odrv4 I__2336 (
            .O(N__12829),
            .I(\this_vga_signals.GZ0Z_296 ));
    Odrv12 I__2335 (
            .O(N__12826),
            .I(\this_vga_signals.GZ0Z_296 ));
    Odrv4 I__2334 (
            .O(N__12821),
            .I(\this_vga_signals.GZ0Z_296 ));
    InMux I__2333 (
            .O(N__12812),
            .I(bfn_15_21_0_));
    InMux I__2332 (
            .O(N__12809),
            .I(N__12802));
    InMux I__2331 (
            .O(N__12808),
            .I(N__12802));
    CascadeMux I__2330 (
            .O(N__12807),
            .I(N__12799));
    LocalMux I__2329 (
            .O(N__12802),
            .I(N__12796));
    InMux I__2328 (
            .O(N__12799),
            .I(N__12793));
    Span4Mux_h I__2327 (
            .O(N__12796),
            .I(N__12788));
    LocalMux I__2326 (
            .O(N__12793),
            .I(N__12788));
    Odrv4 I__2325 (
            .O(N__12788),
            .I(\this_vga_signals.mult1_un40_sum_c3 ));
    CascadeMux I__2324 (
            .O(N__12785),
            .I(\this_vga_signals.mult1_un40_sum_c3_cascade_ ));
    CascadeMux I__2323 (
            .O(N__12782),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a2_x0_cascade_ ));
    CascadeMux I__2322 (
            .O(N__12779),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a2_ns_cascade_ ));
    CascadeMux I__2321 (
            .O(N__12776),
            .I(N__12773));
    InMux I__2320 (
            .O(N__12773),
            .I(N__12770));
    LocalMux I__2319 (
            .O(N__12770),
            .I(\this_vga_signals.mult1_un47_sum_axb2_0_3_1_1 ));
    CascadeMux I__2318 (
            .O(N__12767),
            .I(N__12762));
    InMux I__2317 (
            .O(N__12766),
            .I(N__12759));
    InMux I__2316 (
            .O(N__12765),
            .I(N__12756));
    InMux I__2315 (
            .O(N__12762),
            .I(N__12753));
    LocalMux I__2314 (
            .O(N__12759),
            .I(N__12746));
    LocalMux I__2313 (
            .O(N__12756),
            .I(N__12746));
    LocalMux I__2312 (
            .O(N__12753),
            .I(N__12746));
    Odrv12 I__2311 (
            .O(N__12746),
            .I(\this_vga_signals.M_hcounter_d6_0 ));
    InMux I__2310 (
            .O(N__12743),
            .I(N__12739));
    InMux I__2309 (
            .O(N__12742),
            .I(N__12735));
    LocalMux I__2308 (
            .O(N__12739),
            .I(N__12732));
    InMux I__2307 (
            .O(N__12738),
            .I(N__12729));
    LocalMux I__2306 (
            .O(N__12735),
            .I(N__12726));
    Odrv12 I__2305 (
            .O(N__12732),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__2304 (
            .O(N__12729),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv4 I__2303 (
            .O(N__12726),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    CascadeMux I__2302 (
            .O(N__12719),
            .I(N__12714));
    CascadeMux I__2301 (
            .O(N__12718),
            .I(N__12709));
    CascadeMux I__2300 (
            .O(N__12717),
            .I(N__12706));
    InMux I__2299 (
            .O(N__12714),
            .I(N__12703));
    InMux I__2298 (
            .O(N__12713),
            .I(N__12700));
    CascadeMux I__2297 (
            .O(N__12712),
            .I(N__12697));
    InMux I__2296 (
            .O(N__12709),
            .I(N__12694));
    InMux I__2295 (
            .O(N__12706),
            .I(N__12691));
    LocalMux I__2294 (
            .O(N__12703),
            .I(N__12685));
    LocalMux I__2293 (
            .O(N__12700),
            .I(N__12685));
    InMux I__2292 (
            .O(N__12697),
            .I(N__12682));
    LocalMux I__2291 (
            .O(N__12694),
            .I(N__12679));
    LocalMux I__2290 (
            .O(N__12691),
            .I(N__12676));
    InMux I__2289 (
            .O(N__12690),
            .I(N__12673));
    Span4Mux_v I__2288 (
            .O(N__12685),
            .I(N__12668));
    LocalMux I__2287 (
            .O(N__12682),
            .I(N__12668));
    Odrv4 I__2286 (
            .O(N__12679),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__2285 (
            .O(N__12676),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__2284 (
            .O(N__12673),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__2283 (
            .O(N__12668),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    InMux I__2282 (
            .O(N__12659),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_0 ));
    InMux I__2281 (
            .O(N__12656),
            .I(N__12653));
    LocalMux I__2280 (
            .O(N__12653),
            .I(\this_vga_signals.mult1_un75_sum_c2 ));
    CascadeMux I__2279 (
            .O(N__12650),
            .I(\this_vga_signals.mult1_un82_sum_c3_cascade_ ));
    CascadeMux I__2278 (
            .O(N__12647),
            .I(N__12644));
    CascadeBuf I__2277 (
            .O(N__12644),
            .I(N__12641));
    CascadeMux I__2276 (
            .O(N__12641),
            .I(N__12638));
    CascadeBuf I__2275 (
            .O(N__12638),
            .I(N__12635));
    CascadeMux I__2274 (
            .O(N__12635),
            .I(N__12632));
    CascadeBuf I__2273 (
            .O(N__12632),
            .I(N__12629));
    CascadeMux I__2272 (
            .O(N__12629),
            .I(N__12626));
    CascadeBuf I__2271 (
            .O(N__12626),
            .I(N__12623));
    CascadeMux I__2270 (
            .O(N__12623),
            .I(N__12620));
    CascadeBuf I__2269 (
            .O(N__12620),
            .I(N__12617));
    CascadeMux I__2268 (
            .O(N__12617),
            .I(N__12614));
    CascadeBuf I__2267 (
            .O(N__12614),
            .I(N__12611));
    CascadeMux I__2266 (
            .O(N__12611),
            .I(N__12608));
    CascadeBuf I__2265 (
            .O(N__12608),
            .I(N__12605));
    CascadeMux I__2264 (
            .O(N__12605),
            .I(N__12602));
    CascadeBuf I__2263 (
            .O(N__12602),
            .I(N__12599));
    CascadeMux I__2262 (
            .O(N__12599),
            .I(N__12596));
    CascadeBuf I__2261 (
            .O(N__12596),
            .I(N__12593));
    CascadeMux I__2260 (
            .O(N__12593),
            .I(N__12590));
    CascadeBuf I__2259 (
            .O(N__12590),
            .I(N__12587));
    CascadeMux I__2258 (
            .O(N__12587),
            .I(N__12584));
    CascadeBuf I__2257 (
            .O(N__12584),
            .I(N__12581));
    CascadeMux I__2256 (
            .O(N__12581),
            .I(N__12578));
    CascadeBuf I__2255 (
            .O(N__12578),
            .I(N__12575));
    CascadeMux I__2254 (
            .O(N__12575),
            .I(N__12572));
    CascadeBuf I__2253 (
            .O(N__12572),
            .I(N__12569));
    CascadeMux I__2252 (
            .O(N__12569),
            .I(N__12566));
    CascadeBuf I__2251 (
            .O(N__12566),
            .I(N__12563));
    CascadeMux I__2250 (
            .O(N__12563),
            .I(N__12560));
    CascadeBuf I__2249 (
            .O(N__12560),
            .I(N__12557));
    CascadeMux I__2248 (
            .O(N__12557),
            .I(N__12554));
    InMux I__2247 (
            .O(N__12554),
            .I(N__12551));
    LocalMux I__2246 (
            .O(N__12551),
            .I(N__12548));
    Span4Mux_v I__2245 (
            .O(N__12548),
            .I(N__12545));
    Sp12to4 I__2244 (
            .O(N__12545),
            .I(N__12542));
    Span12Mux_h I__2243 (
            .O(N__12542),
            .I(N__12539));
    Odrv12 I__2242 (
            .O(N__12539),
            .I(M_this_vga_signals_address_7));
    InMux I__2241 (
            .O(N__12536),
            .I(N__12533));
    LocalMux I__2240 (
            .O(N__12533),
            .I(\this_vga_signals.mult1_un68_sum_axbxc1 ));
    CascadeMux I__2239 (
            .O(N__12530),
            .I(\this_vga_signals.mult1_un75_sum_c3_0_cascade_ ));
    InMux I__2238 (
            .O(N__12527),
            .I(N__12524));
    LocalMux I__2237 (
            .O(N__12524),
            .I(\this_vga_signals.mult1_un82_sum_i_1_3 ));
    InMux I__2236 (
            .O(N__12521),
            .I(N__12517));
    InMux I__2235 (
            .O(N__12520),
            .I(N__12514));
    LocalMux I__2234 (
            .O(N__12517),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    LocalMux I__2233 (
            .O(N__12514),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    CascadeMux I__2232 (
            .O(N__12509),
            .I(N__12506));
    InMux I__2231 (
            .O(N__12506),
            .I(N__12503));
    LocalMux I__2230 (
            .O(N__12503),
            .I(N__12499));
    InMux I__2229 (
            .O(N__12502),
            .I(N__12496));
    Odrv4 I__2228 (
            .O(N__12499),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0_0 ));
    LocalMux I__2227 (
            .O(N__12496),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0_0 ));
    InMux I__2226 (
            .O(N__12491),
            .I(N__12484));
    InMux I__2225 (
            .O(N__12490),
            .I(N__12481));
    InMux I__2224 (
            .O(N__12489),
            .I(N__12474));
    InMux I__2223 (
            .O(N__12488),
            .I(N__12474));
    InMux I__2222 (
            .O(N__12487),
            .I(N__12474));
    LocalMux I__2221 (
            .O(N__12484),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3 ));
    LocalMux I__2220 (
            .O(N__12481),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3 ));
    LocalMux I__2219 (
            .O(N__12474),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3 ));
    CascadeMux I__2218 (
            .O(N__12467),
            .I(N__12464));
    CascadeBuf I__2217 (
            .O(N__12464),
            .I(N__12461));
    CascadeMux I__2216 (
            .O(N__12461),
            .I(N__12458));
    CascadeBuf I__2215 (
            .O(N__12458),
            .I(N__12455));
    CascadeMux I__2214 (
            .O(N__12455),
            .I(N__12452));
    CascadeBuf I__2213 (
            .O(N__12452),
            .I(N__12449));
    CascadeMux I__2212 (
            .O(N__12449),
            .I(N__12446));
    CascadeBuf I__2211 (
            .O(N__12446),
            .I(N__12443));
    CascadeMux I__2210 (
            .O(N__12443),
            .I(N__12440));
    CascadeBuf I__2209 (
            .O(N__12440),
            .I(N__12437));
    CascadeMux I__2208 (
            .O(N__12437),
            .I(N__12434));
    CascadeBuf I__2207 (
            .O(N__12434),
            .I(N__12431));
    CascadeMux I__2206 (
            .O(N__12431),
            .I(N__12428));
    CascadeBuf I__2205 (
            .O(N__12428),
            .I(N__12425));
    CascadeMux I__2204 (
            .O(N__12425),
            .I(N__12422));
    CascadeBuf I__2203 (
            .O(N__12422),
            .I(N__12419));
    CascadeMux I__2202 (
            .O(N__12419),
            .I(N__12416));
    CascadeBuf I__2201 (
            .O(N__12416),
            .I(N__12413));
    CascadeMux I__2200 (
            .O(N__12413),
            .I(N__12410));
    CascadeBuf I__2199 (
            .O(N__12410),
            .I(N__12407));
    CascadeMux I__2198 (
            .O(N__12407),
            .I(N__12404));
    CascadeBuf I__2197 (
            .O(N__12404),
            .I(N__12401));
    CascadeMux I__2196 (
            .O(N__12401),
            .I(N__12398));
    CascadeBuf I__2195 (
            .O(N__12398),
            .I(N__12395));
    CascadeMux I__2194 (
            .O(N__12395),
            .I(N__12392));
    CascadeBuf I__2193 (
            .O(N__12392),
            .I(N__12389));
    CascadeMux I__2192 (
            .O(N__12389),
            .I(N__12386));
    CascadeBuf I__2191 (
            .O(N__12386),
            .I(N__12383));
    CascadeMux I__2190 (
            .O(N__12383),
            .I(N__12380));
    CascadeBuf I__2189 (
            .O(N__12380),
            .I(N__12377));
    CascadeMux I__2188 (
            .O(N__12377),
            .I(N__12374));
    InMux I__2187 (
            .O(N__12374),
            .I(N__12371));
    LocalMux I__2186 (
            .O(N__12371),
            .I(N__12368));
    Span4Mux_s2_v I__2185 (
            .O(N__12368),
            .I(N__12365));
    Span4Mux_v I__2184 (
            .O(N__12365),
            .I(N__12362));
    Sp12to4 I__2183 (
            .O(N__12362),
            .I(N__12359));
    Span12Mux_h I__2182 (
            .O(N__12359),
            .I(N__12356));
    Odrv12 I__2181 (
            .O(N__12356),
            .I(M_this_vga_signals_address_10));
    InMux I__2180 (
            .O(N__12353),
            .I(N__12350));
    LocalMux I__2179 (
            .O(N__12350),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_bm ));
    InMux I__2178 (
            .O(N__12347),
            .I(N__12343));
    InMux I__2177 (
            .O(N__12346),
            .I(N__12340));
    LocalMux I__2176 (
            .O(N__12343),
            .I(\this_vga_signals.mult1_un61_sum_axb2 ));
    LocalMux I__2175 (
            .O(N__12340),
            .I(\this_vga_signals.mult1_un61_sum_axb2 ));
    CascadeMux I__2174 (
            .O(N__12335),
            .I(N__12332));
    InMux I__2173 (
            .O(N__12332),
            .I(N__12325));
    InMux I__2172 (
            .O(N__12331),
            .I(N__12325));
    InMux I__2171 (
            .O(N__12330),
            .I(N__12322));
    LocalMux I__2170 (
            .O(N__12325),
            .I(\this_vga_signals.mult1_un61_sum_c2 ));
    LocalMux I__2169 (
            .O(N__12322),
            .I(\this_vga_signals.mult1_un61_sum_c2 ));
    InMux I__2168 (
            .O(N__12317),
            .I(N__12314));
    LocalMux I__2167 (
            .O(N__12314),
            .I(\this_vga_signals.if_N_10 ));
    CascadeMux I__2166 (
            .O(N__12311),
            .I(N__12308));
    CascadeBuf I__2165 (
            .O(N__12308),
            .I(N__12305));
    CascadeMux I__2164 (
            .O(N__12305),
            .I(N__12302));
    CascadeBuf I__2163 (
            .O(N__12302),
            .I(N__12299));
    CascadeMux I__2162 (
            .O(N__12299),
            .I(N__12296));
    CascadeBuf I__2161 (
            .O(N__12296),
            .I(N__12293));
    CascadeMux I__2160 (
            .O(N__12293),
            .I(N__12290));
    CascadeBuf I__2159 (
            .O(N__12290),
            .I(N__12287));
    CascadeMux I__2158 (
            .O(N__12287),
            .I(N__12284));
    CascadeBuf I__2157 (
            .O(N__12284),
            .I(N__12281));
    CascadeMux I__2156 (
            .O(N__12281),
            .I(N__12278));
    CascadeBuf I__2155 (
            .O(N__12278),
            .I(N__12275));
    CascadeMux I__2154 (
            .O(N__12275),
            .I(N__12272));
    CascadeBuf I__2153 (
            .O(N__12272),
            .I(N__12269));
    CascadeMux I__2152 (
            .O(N__12269),
            .I(N__12266));
    CascadeBuf I__2151 (
            .O(N__12266),
            .I(N__12263));
    CascadeMux I__2150 (
            .O(N__12263),
            .I(N__12260));
    CascadeBuf I__2149 (
            .O(N__12260),
            .I(N__12257));
    CascadeMux I__2148 (
            .O(N__12257),
            .I(N__12254));
    CascadeBuf I__2147 (
            .O(N__12254),
            .I(N__12251));
    CascadeMux I__2146 (
            .O(N__12251),
            .I(N__12248));
    CascadeBuf I__2145 (
            .O(N__12248),
            .I(N__12245));
    CascadeMux I__2144 (
            .O(N__12245),
            .I(N__12242));
    CascadeBuf I__2143 (
            .O(N__12242),
            .I(N__12239));
    CascadeMux I__2142 (
            .O(N__12239),
            .I(N__12236));
    CascadeBuf I__2141 (
            .O(N__12236),
            .I(N__12233));
    CascadeMux I__2140 (
            .O(N__12233),
            .I(N__12230));
    CascadeBuf I__2139 (
            .O(N__12230),
            .I(N__12227));
    CascadeMux I__2138 (
            .O(N__12227),
            .I(N__12224));
    CascadeBuf I__2137 (
            .O(N__12224),
            .I(N__12221));
    CascadeMux I__2136 (
            .O(N__12221),
            .I(N__12218));
    InMux I__2135 (
            .O(N__12218),
            .I(N__12215));
    LocalMux I__2134 (
            .O(N__12215),
            .I(N__12212));
    Span4Mux_s3_v I__2133 (
            .O(N__12212),
            .I(N__12209));
    Sp12to4 I__2132 (
            .O(N__12209),
            .I(N__12206));
    Span12Mux_h I__2131 (
            .O(N__12206),
            .I(N__12203));
    Odrv12 I__2130 (
            .O(N__12203),
            .I(M_this_vga_signals_address_9));
    InMux I__2129 (
            .O(N__12200),
            .I(N__12194));
    InMux I__2128 (
            .O(N__12199),
            .I(N__12194));
    LocalMux I__2127 (
            .O(N__12194),
            .I(\this_vga_signals.mult1_un68_sum_axbxc2_0 ));
    InMux I__2126 (
            .O(N__12191),
            .I(N__12183));
    InMux I__2125 (
            .O(N__12190),
            .I(N__12176));
    InMux I__2124 (
            .O(N__12189),
            .I(N__12176));
    InMux I__2123 (
            .O(N__12188),
            .I(N__12176));
    InMux I__2122 (
            .O(N__12187),
            .I(N__12171));
    InMux I__2121 (
            .O(N__12186),
            .I(N__12171));
    LocalMux I__2120 (
            .O(N__12183),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0 ));
    LocalMux I__2119 (
            .O(N__12176),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0 ));
    LocalMux I__2118 (
            .O(N__12171),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0 ));
    InMux I__2117 (
            .O(N__12164),
            .I(N__12161));
    LocalMux I__2116 (
            .O(N__12161),
            .I(\this_vga_signals.mult1_un68_sum_axbxc2 ));
    InMux I__2115 (
            .O(N__12158),
            .I(N__12155));
    LocalMux I__2114 (
            .O(N__12155),
            .I(\this_vga_signals.mult1_un75_sum_c3_0 ));
    CascadeMux I__2113 (
            .O(N__12152),
            .I(\this_vga_signals.mult1_un68_sum_axbxc2_cascade_ ));
    InMux I__2112 (
            .O(N__12149),
            .I(N__12144));
    InMux I__2111 (
            .O(N__12148),
            .I(N__12141));
    InMux I__2110 (
            .O(N__12147),
            .I(N__12138));
    LocalMux I__2109 (
            .O(N__12144),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_0 ));
    LocalMux I__2108 (
            .O(N__12141),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_0 ));
    LocalMux I__2107 (
            .O(N__12138),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_0 ));
    CascadeMux I__2106 (
            .O(N__12131),
            .I(N__12128));
    CascadeBuf I__2105 (
            .O(N__12128),
            .I(N__12125));
    CascadeMux I__2104 (
            .O(N__12125),
            .I(N__12122));
    CascadeBuf I__2103 (
            .O(N__12122),
            .I(N__12119));
    CascadeMux I__2102 (
            .O(N__12119),
            .I(N__12116));
    CascadeBuf I__2101 (
            .O(N__12116),
            .I(N__12113));
    CascadeMux I__2100 (
            .O(N__12113),
            .I(N__12110));
    CascadeBuf I__2099 (
            .O(N__12110),
            .I(N__12107));
    CascadeMux I__2098 (
            .O(N__12107),
            .I(N__12104));
    CascadeBuf I__2097 (
            .O(N__12104),
            .I(N__12101));
    CascadeMux I__2096 (
            .O(N__12101),
            .I(N__12098));
    CascadeBuf I__2095 (
            .O(N__12098),
            .I(N__12095));
    CascadeMux I__2094 (
            .O(N__12095),
            .I(N__12092));
    CascadeBuf I__2093 (
            .O(N__12092),
            .I(N__12089));
    CascadeMux I__2092 (
            .O(N__12089),
            .I(N__12086));
    CascadeBuf I__2091 (
            .O(N__12086),
            .I(N__12083));
    CascadeMux I__2090 (
            .O(N__12083),
            .I(N__12080));
    CascadeBuf I__2089 (
            .O(N__12080),
            .I(N__12077));
    CascadeMux I__2088 (
            .O(N__12077),
            .I(N__12074));
    CascadeBuf I__2087 (
            .O(N__12074),
            .I(N__12071));
    CascadeMux I__2086 (
            .O(N__12071),
            .I(N__12068));
    CascadeBuf I__2085 (
            .O(N__12068),
            .I(N__12065));
    CascadeMux I__2084 (
            .O(N__12065),
            .I(N__12062));
    CascadeBuf I__2083 (
            .O(N__12062),
            .I(N__12059));
    CascadeMux I__2082 (
            .O(N__12059),
            .I(N__12056));
    CascadeBuf I__2081 (
            .O(N__12056),
            .I(N__12053));
    CascadeMux I__2080 (
            .O(N__12053),
            .I(N__12050));
    CascadeBuf I__2079 (
            .O(N__12050),
            .I(N__12047));
    CascadeMux I__2078 (
            .O(N__12047),
            .I(N__12044));
    CascadeBuf I__2077 (
            .O(N__12044),
            .I(N__12041));
    CascadeMux I__2076 (
            .O(N__12041),
            .I(N__12038));
    InMux I__2075 (
            .O(N__12038),
            .I(N__12035));
    LocalMux I__2074 (
            .O(N__12035),
            .I(N__12032));
    Span4Mux_h I__2073 (
            .O(N__12032),
            .I(N__12029));
    Span4Mux_h I__2072 (
            .O(N__12029),
            .I(N__12026));
    Sp12to4 I__2071 (
            .O(N__12026),
            .I(N__12023));
    Span12Mux_v I__2070 (
            .O(N__12023),
            .I(N__12020));
    Odrv12 I__2069 (
            .O(N__12020),
            .I(M_this_vga_signals_address_8));
    CascadeMux I__2068 (
            .O(N__12017),
            .I(\this_vga_signals.M_vcounter_d7lt9_cascade_ ));
    InMux I__2067 (
            .O(N__12014),
            .I(N__12011));
    LocalMux I__2066 (
            .O(N__12011),
            .I(\this_vga_signals.M_vcounter_d7lto8_1 ));
    CascadeMux I__2065 (
            .O(N__12008),
            .I(\this_vga_signals.un6_vvisibilitylt9_0_cascade_ ));
    InMux I__2064 (
            .O(N__12005),
            .I(N__12001));
    InMux I__2063 (
            .O(N__12004),
            .I(N__11998));
    LocalMux I__2062 (
            .O(N__12001),
            .I(\this_vga_signals.vaddress_c5_i ));
    LocalMux I__2061 (
            .O(N__11998),
            .I(\this_vga_signals.vaddress_c5_i ));
    InMux I__2060 (
            .O(N__11993),
            .I(N__11990));
    LocalMux I__2059 (
            .O(N__11990),
            .I(N__11985));
    InMux I__2058 (
            .O(N__11989),
            .I(N__11982));
    InMux I__2057 (
            .O(N__11988),
            .I(N__11979));
    Span4Mux_h I__2056 (
            .O(N__11985),
            .I(N__11976));
    LocalMux I__2055 (
            .O(N__11982),
            .I(N__11973));
    LocalMux I__2054 (
            .O(N__11979),
            .I(N__11969));
    Span4Mux_v I__2053 (
            .O(N__11976),
            .I(N__11964));
    Span4Mux_v I__2052 (
            .O(N__11973),
            .I(N__11964));
    InMux I__2051 (
            .O(N__11972),
            .I(N__11961));
    Span12Mux_h I__2050 (
            .O(N__11969),
            .I(N__11958));
    Span4Mux_h I__2049 (
            .O(N__11964),
            .I(N__11953));
    LocalMux I__2048 (
            .O(N__11961),
            .I(N__11953));
    Odrv12 I__2047 (
            .O(N__11958),
            .I(\this_vga_signals.vvisibility ));
    Odrv4 I__2046 (
            .O(N__11953),
            .I(\this_vga_signals.vvisibility ));
    CascadeMux I__2045 (
            .O(N__11948),
            .I(\this_vga_signals.vsync_1_0_cascade_ ));
    InMux I__2044 (
            .O(N__11945),
            .I(N__11942));
    LocalMux I__2043 (
            .O(N__11942),
            .I(\this_vga_signals.vsync_1_4 ));
    InMux I__2042 (
            .O(N__11939),
            .I(N__11936));
    LocalMux I__2041 (
            .O(N__11936),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_ns_1 ));
    InMux I__2040 (
            .O(N__11933),
            .I(N__11924));
    InMux I__2039 (
            .O(N__11932),
            .I(N__11924));
    InMux I__2038 (
            .O(N__11931),
            .I(N__11924));
    LocalMux I__2037 (
            .O(N__11924),
            .I(N__11921));
    Odrv4 I__2036 (
            .O(N__11921),
            .I(\this_vga_signals.SUM_2 ));
    InMux I__2035 (
            .O(N__11918),
            .I(N__11915));
    LocalMux I__2034 (
            .O(N__11915),
            .I(\this_vga_signals.mult1_un47_sum_c2 ));
    InMux I__2033 (
            .O(N__11912),
            .I(N__11908));
    InMux I__2032 (
            .O(N__11911),
            .I(N__11905));
    LocalMux I__2031 (
            .O(N__11908),
            .I(\this_vga_signals.mult1_un47_sum_axb2_0_3 ));
    LocalMux I__2030 (
            .O(N__11905),
            .I(\this_vga_signals.mult1_un47_sum_axb2_0_3 ));
    CascadeMux I__2029 (
            .O(N__11900),
            .I(\this_vga_signals.mult1_un47_sum_c2_cascade_ ));
    InMux I__2028 (
            .O(N__11897),
            .I(N__11891));
    InMux I__2027 (
            .O(N__11896),
            .I(N__11891));
    LocalMux I__2026 (
            .O(N__11891),
            .I(N__11888));
    Odrv4 I__2025 (
            .O(N__11888),
            .I(\this_vga_signals.vaddress_6 ));
    InMux I__2024 (
            .O(N__11885),
            .I(N__11882));
    LocalMux I__2023 (
            .O(N__11882),
            .I(\this_vga_signals.mult1_un47_sum_axb2_3_tz ));
    CascadeMux I__2022 (
            .O(N__11879),
            .I(N__11875));
    CascadeMux I__2021 (
            .O(N__11878),
            .I(N__11872));
    InMux I__2020 (
            .O(N__11875),
            .I(N__11863));
    InMux I__2019 (
            .O(N__11872),
            .I(N__11863));
    InMux I__2018 (
            .O(N__11871),
            .I(N__11863));
    CascadeMux I__2017 (
            .O(N__11870),
            .I(N__11860));
    LocalMux I__2016 (
            .O(N__11863),
            .I(N__11857));
    InMux I__2015 (
            .O(N__11860),
            .I(N__11854));
    Odrv4 I__2014 (
            .O(N__11857),
            .I(\this_vga_signals.vaddress_7 ));
    LocalMux I__2013 (
            .O(N__11854),
            .I(\this_vga_signals.vaddress_7 ));
    CascadeMux I__2012 (
            .O(N__11849),
            .I(\this_vga_signals.M_vcounter_d7lt8_0_cascade_ ));
    CascadeMux I__2011 (
            .O(N__11846),
            .I(\this_vga_signals.mult1_un54_sum_c2_cascade_ ));
    CascadeMux I__2010 (
            .O(N__11843),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_cascade_ ));
    CascadeMux I__2009 (
            .O(N__11840),
            .I(\this_vga_signals.mult1_un61_sum_c2_cascade_ ));
    InMux I__2008 (
            .O(N__11837),
            .I(N__11832));
    InMux I__2007 (
            .O(N__11836),
            .I(N__11827));
    InMux I__2006 (
            .O(N__11835),
            .I(N__11827));
    LocalMux I__2005 (
            .O(N__11832),
            .I(\this_vga_signals.mult1_un54_sum_axb1_i ));
    LocalMux I__2004 (
            .O(N__11827),
            .I(\this_vga_signals.mult1_un54_sum_axb1_i ));
    InMux I__2003 (
            .O(N__11822),
            .I(N__11818));
    InMux I__2002 (
            .O(N__11821),
            .I(N__11815));
    LocalMux I__2001 (
            .O(N__11818),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1_2 ));
    LocalMux I__2000 (
            .O(N__11815),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1_2 ));
    CascadeMux I__1999 (
            .O(N__11810),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1_2_cascade_ ));
    CascadeMux I__1998 (
            .O(N__11807),
            .I(N__11804));
    InMux I__1997 (
            .O(N__11804),
            .I(N__11799));
    InMux I__1996 (
            .O(N__11803),
            .I(N__11794));
    InMux I__1995 (
            .O(N__11802),
            .I(N__11794));
    LocalMux I__1994 (
            .O(N__11799),
            .I(\this_vga_signals.mult1_un40_sum_c2 ));
    LocalMux I__1993 (
            .O(N__11794),
            .I(\this_vga_signals.mult1_un40_sum_c2 ));
    InMux I__1992 (
            .O(N__11789),
            .I(N__11785));
    InMux I__1991 (
            .O(N__11788),
            .I(N__11782));
    LocalMux I__1990 (
            .O(N__11785),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3 ));
    LocalMux I__1989 (
            .O(N__11782),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3 ));
    CascadeMux I__1988 (
            .O(N__11777),
            .I(\this_vga_signals.mult1_un54_sum_axb1_0_cascade_ ));
    InMux I__1987 (
            .O(N__11774),
            .I(N__11769));
    InMux I__1986 (
            .O(N__11773),
            .I(N__11764));
    InMux I__1985 (
            .O(N__11772),
            .I(N__11764));
    LocalMux I__1984 (
            .O(N__11769),
            .I(\this_vga_signals.mult1_un47_sum_ac0_4 ));
    LocalMux I__1983 (
            .O(N__11764),
            .I(\this_vga_signals.mult1_un47_sum_ac0_4 ));
    CascadeMux I__1982 (
            .O(N__11759),
            .I(N__11756));
    InMux I__1981 (
            .O(N__11756),
            .I(N__11753));
    LocalMux I__1980 (
            .O(N__11753),
            .I(\this_vga_signals.un2_vsynclt8 ));
    IoInMux I__1979 (
            .O(N__11750),
            .I(N__11747));
    LocalMux I__1978 (
            .O(N__11747),
            .I(N__11744));
    Span4Mux_s0_v I__1977 (
            .O(N__11744),
            .I(N__11741));
    Sp12to4 I__1976 (
            .O(N__11741),
            .I(N__11738));
    Span12Mux_h I__1975 (
            .O(N__11738),
            .I(N__11735));
    Odrv12 I__1974 (
            .O(N__11735),
            .I(this_vga_signals_vsync_1_i));
    CascadeMux I__1973 (
            .O(N__11732),
            .I(N__11729));
    CascadeBuf I__1972 (
            .O(N__11729),
            .I(N__11726));
    CascadeMux I__1971 (
            .O(N__11726),
            .I(N__11723));
    CascadeBuf I__1970 (
            .O(N__11723),
            .I(N__11720));
    CascadeMux I__1969 (
            .O(N__11720),
            .I(N__11717));
    CascadeBuf I__1968 (
            .O(N__11717),
            .I(N__11714));
    CascadeMux I__1967 (
            .O(N__11714),
            .I(N__11711));
    CascadeBuf I__1966 (
            .O(N__11711),
            .I(N__11708));
    CascadeMux I__1965 (
            .O(N__11708),
            .I(N__11705));
    CascadeBuf I__1964 (
            .O(N__11705),
            .I(N__11702));
    CascadeMux I__1963 (
            .O(N__11702),
            .I(N__11699));
    CascadeBuf I__1962 (
            .O(N__11699),
            .I(N__11696));
    CascadeMux I__1961 (
            .O(N__11696),
            .I(N__11693));
    CascadeBuf I__1960 (
            .O(N__11693),
            .I(N__11690));
    CascadeMux I__1959 (
            .O(N__11690),
            .I(N__11687));
    CascadeBuf I__1958 (
            .O(N__11687),
            .I(N__11684));
    CascadeMux I__1957 (
            .O(N__11684),
            .I(N__11681));
    CascadeBuf I__1956 (
            .O(N__11681),
            .I(N__11678));
    CascadeMux I__1955 (
            .O(N__11678),
            .I(N__11675));
    CascadeBuf I__1954 (
            .O(N__11675),
            .I(N__11672));
    CascadeMux I__1953 (
            .O(N__11672),
            .I(N__11669));
    CascadeBuf I__1952 (
            .O(N__11669),
            .I(N__11666));
    CascadeMux I__1951 (
            .O(N__11666),
            .I(N__11663));
    CascadeBuf I__1950 (
            .O(N__11663),
            .I(N__11660));
    CascadeMux I__1949 (
            .O(N__11660),
            .I(N__11657));
    CascadeBuf I__1948 (
            .O(N__11657),
            .I(N__11654));
    CascadeMux I__1947 (
            .O(N__11654),
            .I(N__11651));
    CascadeBuf I__1946 (
            .O(N__11651),
            .I(N__11648));
    CascadeMux I__1945 (
            .O(N__11648),
            .I(N__11645));
    CascadeBuf I__1944 (
            .O(N__11645),
            .I(N__11642));
    CascadeMux I__1943 (
            .O(N__11642),
            .I(N__11639));
    InMux I__1942 (
            .O(N__11639),
            .I(N__11636));
    LocalMux I__1941 (
            .O(N__11636),
            .I(N__11633));
    Span4Mux_v I__1940 (
            .O(N__11633),
            .I(N__11630));
    Sp12to4 I__1939 (
            .O(N__11630),
            .I(N__11627));
    Span12Mux_h I__1938 (
            .O(N__11627),
            .I(N__11624));
    Odrv12 I__1937 (
            .O(N__11624),
            .I(M_this_vga_signals_address_6));
    InMux I__1936 (
            .O(N__11621),
            .I(N__11618));
    LocalMux I__1935 (
            .O(N__11618),
            .I(\this_vga_signals.if_N_9 ));
    CascadeMux I__1934 (
            .O(N__11615),
            .I(\this_vga_signals.if_N_10_cascade_ ));
    CascadeMux I__1933 (
            .O(N__11612),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_0_cascade_ ));
    IoInMux I__1932 (
            .O(N__11609),
            .I(N__11606));
    LocalMux I__1931 (
            .O(N__11606),
            .I(N__11603));
    IoSpan4Mux I__1930 (
            .O(N__11603),
            .I(N__11598));
    InMux I__1929 (
            .O(N__11602),
            .I(N__11595));
    InMux I__1928 (
            .O(N__11601),
            .I(N__11592));
    Span4Mux_s2_v I__1927 (
            .O(N__11598),
            .I(N__11589));
    LocalMux I__1926 (
            .O(N__11595),
            .I(N__11586));
    LocalMux I__1925 (
            .O(N__11592),
            .I(N__11583));
    Sp12to4 I__1924 (
            .O(N__11589),
            .I(N__11580));
    Span4Mux_h I__1923 (
            .O(N__11586),
            .I(N__11577));
    Span4Mux_h I__1922 (
            .O(N__11583),
            .I(N__11574));
    Span12Mux_v I__1921 (
            .O(N__11580),
            .I(N__11570));
    Span4Mux_h I__1920 (
            .O(N__11577),
            .I(N__11565));
    Span4Mux_h I__1919 (
            .O(N__11574),
            .I(N__11565));
    InMux I__1918 (
            .O(N__11573),
            .I(N__11562));
    Odrv12 I__1917 (
            .O(N__11570),
            .I(debug_c_1));
    Odrv4 I__1916 (
            .O(N__11565),
            .I(debug_c_1));
    LocalMux I__1915 (
            .O(N__11562),
            .I(debug_c_1));
    CascadeMux I__1914 (
            .O(N__11555),
            .I(N__11551));
    CascadeMux I__1913 (
            .O(N__11554),
            .I(N__11545));
    InMux I__1912 (
            .O(N__11551),
            .I(N__11542));
    CascadeMux I__1911 (
            .O(N__11550),
            .I(N__11538));
    InMux I__1910 (
            .O(N__11549),
            .I(N__11535));
    InMux I__1909 (
            .O(N__11548),
            .I(N__11532));
    InMux I__1908 (
            .O(N__11545),
            .I(N__11529));
    LocalMux I__1907 (
            .O(N__11542),
            .I(N__11525));
    InMux I__1906 (
            .O(N__11541),
            .I(N__11522));
    InMux I__1905 (
            .O(N__11538),
            .I(N__11519));
    LocalMux I__1904 (
            .O(N__11535),
            .I(N__11514));
    LocalMux I__1903 (
            .O(N__11532),
            .I(N__11514));
    LocalMux I__1902 (
            .O(N__11529),
            .I(N__11510));
    InMux I__1901 (
            .O(N__11528),
            .I(N__11507));
    Span4Mux_v I__1900 (
            .O(N__11525),
            .I(N__11498));
    LocalMux I__1899 (
            .O(N__11522),
            .I(N__11498));
    LocalMux I__1898 (
            .O(N__11519),
            .I(N__11498));
    Span4Mux_h I__1897 (
            .O(N__11514),
            .I(N__11498));
    InMux I__1896 (
            .O(N__11513),
            .I(N__11495));
    Span4Mux_h I__1895 (
            .O(N__11510),
            .I(N__11492));
    LocalMux I__1894 (
            .O(N__11507),
            .I(N__11487));
    Span4Mux_h I__1893 (
            .O(N__11498),
            .I(N__11487));
    LocalMux I__1892 (
            .O(N__11495),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__1891 (
            .O(N__11492),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__1890 (
            .O(N__11487),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    CascadeMux I__1889 (
            .O(N__11480),
            .I(N__11477));
    InMux I__1888 (
            .O(N__11477),
            .I(N__11472));
    InMux I__1887 (
            .O(N__11476),
            .I(N__11464));
    InMux I__1886 (
            .O(N__11475),
            .I(N__11461));
    LocalMux I__1885 (
            .O(N__11472),
            .I(N__11458));
    InMux I__1884 (
            .O(N__11471),
            .I(N__11455));
    InMux I__1883 (
            .O(N__11470),
            .I(N__11452));
    InMux I__1882 (
            .O(N__11469),
            .I(N__11447));
    InMux I__1881 (
            .O(N__11468),
            .I(N__11447));
    CascadeMux I__1880 (
            .O(N__11467),
            .I(N__11442));
    LocalMux I__1879 (
            .O(N__11464),
            .I(N__11436));
    LocalMux I__1878 (
            .O(N__11461),
            .I(N__11436));
    Span4Mux_h I__1877 (
            .O(N__11458),
            .I(N__11431));
    LocalMux I__1876 (
            .O(N__11455),
            .I(N__11431));
    LocalMux I__1875 (
            .O(N__11452),
            .I(N__11428));
    LocalMux I__1874 (
            .O(N__11447),
            .I(N__11425));
    InMux I__1873 (
            .O(N__11446),
            .I(N__11422));
    InMux I__1872 (
            .O(N__11445),
            .I(N__11419));
    InMux I__1871 (
            .O(N__11442),
            .I(N__11415));
    InMux I__1870 (
            .O(N__11441),
            .I(N__11412));
    Span4Mux_v I__1869 (
            .O(N__11436),
            .I(N__11409));
    Span4Mux_h I__1868 (
            .O(N__11431),
            .I(N__11406));
    Span4Mux_h I__1867 (
            .O(N__11428),
            .I(N__11397));
    Span4Mux_h I__1866 (
            .O(N__11425),
            .I(N__11397));
    LocalMux I__1865 (
            .O(N__11422),
            .I(N__11397));
    LocalMux I__1864 (
            .O(N__11419),
            .I(N__11397));
    InMux I__1863 (
            .O(N__11418),
            .I(N__11394));
    LocalMux I__1862 (
            .O(N__11415),
            .I(N__11391));
    LocalMux I__1861 (
            .O(N__11412),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__1860 (
            .O(N__11409),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__1859 (
            .O(N__11406),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__1858 (
            .O(N__11397),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__1857 (
            .O(N__11394),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv12 I__1856 (
            .O(N__11391),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    InMux I__1855 (
            .O(N__11378),
            .I(N__11375));
    LocalMux I__1854 (
            .O(N__11375),
            .I(\this_vga_signals.g0_0_a2_1 ));
    InMux I__1853 (
            .O(N__11372),
            .I(N__11369));
    LocalMux I__1852 (
            .O(N__11369),
            .I(N__11366));
    Span4Mux_v I__1851 (
            .O(N__11366),
            .I(N__11363));
    Sp12to4 I__1850 (
            .O(N__11363),
            .I(N__11360));
    Odrv12 I__1849 (
            .O(N__11360),
            .I(\this_delay_clk.M_pipe_qZ0Z_1 ));
    InMux I__1848 (
            .O(N__11357),
            .I(N__11354));
    LocalMux I__1847 (
            .O(N__11354),
            .I(\this_delay_clk.M_pipe_qZ0Z_2 ));
    CascadeMux I__1846 (
            .O(N__11351),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0_0_cascade_ ));
    CascadeMux I__1845 (
            .O(N__11348),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_cascade_ ));
    InMux I__1844 (
            .O(N__11345),
            .I(N__11342));
    LocalMux I__1843 (
            .O(N__11342),
            .I(N__11330));
    SRMux I__1842 (
            .O(N__11341),
            .I(N__11309));
    SRMux I__1841 (
            .O(N__11340),
            .I(N__11309));
    SRMux I__1840 (
            .O(N__11339),
            .I(N__11309));
    SRMux I__1839 (
            .O(N__11338),
            .I(N__11309));
    SRMux I__1838 (
            .O(N__11337),
            .I(N__11309));
    SRMux I__1837 (
            .O(N__11336),
            .I(N__11309));
    SRMux I__1836 (
            .O(N__11335),
            .I(N__11309));
    SRMux I__1835 (
            .O(N__11334),
            .I(N__11309));
    SRMux I__1834 (
            .O(N__11333),
            .I(N__11309));
    Glb2LocalMux I__1833 (
            .O(N__11330),
            .I(N__11309));
    GlobalMux I__1832 (
            .O(N__11309),
            .I(N__11306));
    gio2CtrlBuf I__1831 (
            .O(N__11306),
            .I(\this_vga_signals.N_583_g ));
    InMux I__1830 (
            .O(N__11303),
            .I(N__11298));
    InMux I__1829 (
            .O(N__11302),
            .I(N__11295));
    InMux I__1828 (
            .O(N__11301),
            .I(N__11292));
    LocalMux I__1827 (
            .O(N__11298),
            .I(N__11289));
    LocalMux I__1826 (
            .O(N__11295),
            .I(N__11284));
    LocalMux I__1825 (
            .O(N__11292),
            .I(N__11284));
    Sp12to4 I__1824 (
            .O(N__11289),
            .I(N__11281));
    Odrv4 I__1823 (
            .O(N__11284),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRDZ0 ));
    Odrv12 I__1822 (
            .O(N__11281),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRDZ0 ));
    InMux I__1821 (
            .O(N__11276),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    InMux I__1820 (
            .O(N__11273),
            .I(N__11268));
    InMux I__1819 (
            .O(N__11272),
            .I(N__11263));
    InMux I__1818 (
            .O(N__11271),
            .I(N__11263));
    LocalMux I__1817 (
            .O(N__11268),
            .I(N__11260));
    LocalMux I__1816 (
            .O(N__11263),
            .I(N__11257));
    Span4Mux_h I__1815 (
            .O(N__11260),
            .I(N__11254));
    Span4Mux_h I__1814 (
            .O(N__11257),
            .I(N__11251));
    Odrv4 I__1813 (
            .O(N__11254),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0 ));
    Odrv4 I__1812 (
            .O(N__11251),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0 ));
    InMux I__1811 (
            .O(N__11246),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    InMux I__1810 (
            .O(N__11243),
            .I(N__11236));
    InMux I__1809 (
            .O(N__11242),
            .I(N__11236));
    InMux I__1808 (
            .O(N__11241),
            .I(N__11233));
    LocalMux I__1807 (
            .O(N__11236),
            .I(N__11228));
    LocalMux I__1806 (
            .O(N__11233),
            .I(N__11228));
    Span4Mux_h I__1805 (
            .O(N__11228),
            .I(N__11225));
    Odrv4 I__1804 (
            .O(N__11225),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0 ));
    InMux I__1803 (
            .O(N__11222),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__1802 (
            .O(N__11219),
            .I(N__11214));
    InMux I__1801 (
            .O(N__11218),
            .I(N__11211));
    InMux I__1800 (
            .O(N__11217),
            .I(N__11208));
    LocalMux I__1799 (
            .O(N__11214),
            .I(N__11205));
    LocalMux I__1798 (
            .O(N__11211),
            .I(N__11202));
    LocalMux I__1797 (
            .O(N__11208),
            .I(N__11199));
    Span4Mux_h I__1796 (
            .O(N__11205),
            .I(N__11196));
    Span4Mux_v I__1795 (
            .O(N__11202),
            .I(N__11191));
    Span4Mux_h I__1794 (
            .O(N__11199),
            .I(N__11191));
    Odrv4 I__1793 (
            .O(N__11196),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0 ));
    Odrv4 I__1792 (
            .O(N__11191),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0 ));
    InMux I__1791 (
            .O(N__11186),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__1790 (
            .O(N__11183),
            .I(bfn_12_21_0_));
    InMux I__1789 (
            .O(N__11180),
            .I(N__11175));
    InMux I__1788 (
            .O(N__11179),
            .I(N__11172));
    InMux I__1787 (
            .O(N__11178),
            .I(N__11169));
    LocalMux I__1786 (
            .O(N__11175),
            .I(N__11164));
    LocalMux I__1785 (
            .O(N__11172),
            .I(N__11164));
    LocalMux I__1784 (
            .O(N__11169),
            .I(N__11161));
    Span4Mux_h I__1783 (
            .O(N__11164),
            .I(N__11158));
    Span4Mux_v I__1782 (
            .O(N__11161),
            .I(N__11155));
    Odrv4 I__1781 (
            .O(N__11158),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0 ));
    Odrv4 I__1780 (
            .O(N__11155),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0 ));
    CascadeMux I__1779 (
            .O(N__11150),
            .I(N__11145));
    InMux I__1778 (
            .O(N__11149),
            .I(N__11139));
    InMux I__1777 (
            .O(N__11148),
            .I(N__11136));
    InMux I__1776 (
            .O(N__11145),
            .I(N__11133));
    CascadeMux I__1775 (
            .O(N__11144),
            .I(N__11128));
    CascadeMux I__1774 (
            .O(N__11143),
            .I(N__11125));
    CascadeMux I__1773 (
            .O(N__11142),
            .I(N__11119));
    LocalMux I__1772 (
            .O(N__11139),
            .I(N__11111));
    LocalMux I__1771 (
            .O(N__11136),
            .I(N__11111));
    LocalMux I__1770 (
            .O(N__11133),
            .I(N__11107));
    InMux I__1769 (
            .O(N__11132),
            .I(N__11100));
    InMux I__1768 (
            .O(N__11131),
            .I(N__11100));
    InMux I__1767 (
            .O(N__11128),
            .I(N__11100));
    InMux I__1766 (
            .O(N__11125),
            .I(N__11097));
    InMux I__1765 (
            .O(N__11124),
            .I(N__11094));
    CascadeMux I__1764 (
            .O(N__11123),
            .I(N__11089));
    InMux I__1763 (
            .O(N__11122),
            .I(N__11081));
    InMux I__1762 (
            .O(N__11119),
            .I(N__11072));
    InMux I__1761 (
            .O(N__11118),
            .I(N__11072));
    InMux I__1760 (
            .O(N__11117),
            .I(N__11072));
    InMux I__1759 (
            .O(N__11116),
            .I(N__11072));
    Span4Mux_v I__1758 (
            .O(N__11111),
            .I(N__11069));
    InMux I__1757 (
            .O(N__11110),
            .I(N__11066));
    Span4Mux_h I__1756 (
            .O(N__11107),
            .I(N__11061));
    LocalMux I__1755 (
            .O(N__11100),
            .I(N__11061));
    LocalMux I__1754 (
            .O(N__11097),
            .I(N__11058));
    LocalMux I__1753 (
            .O(N__11094),
            .I(N__11055));
    InMux I__1752 (
            .O(N__11093),
            .I(N__11050));
    InMux I__1751 (
            .O(N__11092),
            .I(N__11050));
    InMux I__1750 (
            .O(N__11089),
            .I(N__11047));
    InMux I__1749 (
            .O(N__11088),
            .I(N__11042));
    InMux I__1748 (
            .O(N__11087),
            .I(N__11042));
    InMux I__1747 (
            .O(N__11086),
            .I(N__11037));
    InMux I__1746 (
            .O(N__11085),
            .I(N__11037));
    InMux I__1745 (
            .O(N__11084),
            .I(N__11034));
    LocalMux I__1744 (
            .O(N__11081),
            .I(N__11027));
    LocalMux I__1743 (
            .O(N__11072),
            .I(N__11027));
    Span4Mux_h I__1742 (
            .O(N__11069),
            .I(N__11027));
    LocalMux I__1741 (
            .O(N__11066),
            .I(N__11022));
    Span4Mux_h I__1740 (
            .O(N__11061),
            .I(N__11022));
    Span4Mux_v I__1739 (
            .O(N__11058),
            .I(N__11013));
    Span4Mux_v I__1738 (
            .O(N__11055),
            .I(N__11013));
    LocalMux I__1737 (
            .O(N__11050),
            .I(N__11013));
    LocalMux I__1736 (
            .O(N__11047),
            .I(N__11013));
    LocalMux I__1735 (
            .O(N__11042),
            .I(N__11010));
    LocalMux I__1734 (
            .O(N__11037),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__1733 (
            .O(N__11034),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1732 (
            .O(N__11027),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1731 (
            .O(N__11022),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1730 (
            .O(N__11013),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv12 I__1729 (
            .O(N__11010),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    CascadeMux I__1728 (
            .O(N__10997),
            .I(N__10993));
    InMux I__1727 (
            .O(N__10996),
            .I(N__10987));
    InMux I__1726 (
            .O(N__10993),
            .I(N__10984));
    CascadeMux I__1725 (
            .O(N__10992),
            .I(N__10976));
    CascadeMux I__1724 (
            .O(N__10991),
            .I(N__10969));
    CascadeMux I__1723 (
            .O(N__10990),
            .I(N__10966));
    LocalMux I__1722 (
            .O(N__10987),
            .I(N__10958));
    LocalMux I__1721 (
            .O(N__10984),
            .I(N__10958));
    InMux I__1720 (
            .O(N__10983),
            .I(N__10955));
    InMux I__1719 (
            .O(N__10982),
            .I(N__10952));
    InMux I__1718 (
            .O(N__10981),
            .I(N__10949));
    InMux I__1717 (
            .O(N__10980),
            .I(N__10946));
    CascadeMux I__1716 (
            .O(N__10979),
            .I(N__10942));
    InMux I__1715 (
            .O(N__10976),
            .I(N__10939));
    InMux I__1714 (
            .O(N__10975),
            .I(N__10936));
    InMux I__1713 (
            .O(N__10974),
            .I(N__10933));
    CascadeMux I__1712 (
            .O(N__10973),
            .I(N__10928));
    CascadeMux I__1711 (
            .O(N__10972),
            .I(N__10925));
    InMux I__1710 (
            .O(N__10969),
            .I(N__10916));
    InMux I__1709 (
            .O(N__10966),
            .I(N__10916));
    InMux I__1708 (
            .O(N__10965),
            .I(N__10916));
    InMux I__1707 (
            .O(N__10964),
            .I(N__10911));
    InMux I__1706 (
            .O(N__10963),
            .I(N__10911));
    Span4Mux_h I__1705 (
            .O(N__10958),
            .I(N__10899));
    LocalMux I__1704 (
            .O(N__10955),
            .I(N__10899));
    LocalMux I__1703 (
            .O(N__10952),
            .I(N__10899));
    LocalMux I__1702 (
            .O(N__10949),
            .I(N__10894));
    LocalMux I__1701 (
            .O(N__10946),
            .I(N__10894));
    InMux I__1700 (
            .O(N__10945),
            .I(N__10889));
    InMux I__1699 (
            .O(N__10942),
            .I(N__10889));
    LocalMux I__1698 (
            .O(N__10939),
            .I(N__10886));
    LocalMux I__1697 (
            .O(N__10936),
            .I(N__10883));
    LocalMux I__1696 (
            .O(N__10933),
            .I(N__10880));
    InMux I__1695 (
            .O(N__10932),
            .I(N__10877));
    InMux I__1694 (
            .O(N__10931),
            .I(N__10874));
    InMux I__1693 (
            .O(N__10928),
            .I(N__10867));
    InMux I__1692 (
            .O(N__10925),
            .I(N__10867));
    InMux I__1691 (
            .O(N__10924),
            .I(N__10867));
    InMux I__1690 (
            .O(N__10923),
            .I(N__10864));
    LocalMux I__1689 (
            .O(N__10916),
            .I(N__10861));
    LocalMux I__1688 (
            .O(N__10911),
            .I(N__10858));
    InMux I__1687 (
            .O(N__10910),
            .I(N__10855));
    InMux I__1686 (
            .O(N__10909),
            .I(N__10852));
    InMux I__1685 (
            .O(N__10908),
            .I(N__10847));
    InMux I__1684 (
            .O(N__10907),
            .I(N__10847));
    InMux I__1683 (
            .O(N__10906),
            .I(N__10844));
    Span4Mux_h I__1682 (
            .O(N__10899),
            .I(N__10841));
    Span4Mux_v I__1681 (
            .O(N__10894),
            .I(N__10834));
    LocalMux I__1680 (
            .O(N__10889),
            .I(N__10834));
    Span4Mux_h I__1679 (
            .O(N__10886),
            .I(N__10834));
    Span4Mux_h I__1678 (
            .O(N__10883),
            .I(N__10831));
    Span4Mux_v I__1677 (
            .O(N__10880),
            .I(N__10826));
    LocalMux I__1676 (
            .O(N__10877),
            .I(N__10826));
    LocalMux I__1675 (
            .O(N__10874),
            .I(N__10821));
    LocalMux I__1674 (
            .O(N__10867),
            .I(N__10821));
    LocalMux I__1673 (
            .O(N__10864),
            .I(N__10814));
    Span4Mux_h I__1672 (
            .O(N__10861),
            .I(N__10814));
    Span4Mux_h I__1671 (
            .O(N__10858),
            .I(N__10814));
    LocalMux I__1670 (
            .O(N__10855),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1669 (
            .O(N__10852),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1668 (
            .O(N__10847),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1667 (
            .O(N__10844),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1666 (
            .O(N__10841),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1665 (
            .O(N__10834),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1664 (
            .O(N__10831),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1663 (
            .O(N__10826),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv12 I__1662 (
            .O(N__10821),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1661 (
            .O(N__10814),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    CascadeMux I__1660 (
            .O(N__10793),
            .I(N__10790));
    InMux I__1659 (
            .O(N__10790),
            .I(N__10787));
    LocalMux I__1658 (
            .O(N__10787),
            .I(\this_vga_signals.g0_4_0 ));
    CascadeMux I__1657 (
            .O(N__10784),
            .I(N__10781));
    CascadeBuf I__1656 (
            .O(N__10781),
            .I(N__10778));
    CascadeMux I__1655 (
            .O(N__10778),
            .I(N__10775));
    CascadeBuf I__1654 (
            .O(N__10775),
            .I(N__10772));
    CascadeMux I__1653 (
            .O(N__10772),
            .I(N__10769));
    CascadeBuf I__1652 (
            .O(N__10769),
            .I(N__10766));
    CascadeMux I__1651 (
            .O(N__10766),
            .I(N__10763));
    CascadeBuf I__1650 (
            .O(N__10763),
            .I(N__10760));
    CascadeMux I__1649 (
            .O(N__10760),
            .I(N__10757));
    CascadeBuf I__1648 (
            .O(N__10757),
            .I(N__10754));
    CascadeMux I__1647 (
            .O(N__10754),
            .I(N__10751));
    CascadeBuf I__1646 (
            .O(N__10751),
            .I(N__10748));
    CascadeMux I__1645 (
            .O(N__10748),
            .I(N__10745));
    CascadeBuf I__1644 (
            .O(N__10745),
            .I(N__10742));
    CascadeMux I__1643 (
            .O(N__10742),
            .I(N__10739));
    CascadeBuf I__1642 (
            .O(N__10739),
            .I(N__10736));
    CascadeMux I__1641 (
            .O(N__10736),
            .I(N__10733));
    CascadeBuf I__1640 (
            .O(N__10733),
            .I(N__10730));
    CascadeMux I__1639 (
            .O(N__10730),
            .I(N__10727));
    CascadeBuf I__1638 (
            .O(N__10727),
            .I(N__10724));
    CascadeMux I__1637 (
            .O(N__10724),
            .I(N__10721));
    CascadeBuf I__1636 (
            .O(N__10721),
            .I(N__10718));
    CascadeMux I__1635 (
            .O(N__10718),
            .I(N__10715));
    CascadeBuf I__1634 (
            .O(N__10715),
            .I(N__10712));
    CascadeMux I__1633 (
            .O(N__10712),
            .I(N__10709));
    CascadeBuf I__1632 (
            .O(N__10709),
            .I(N__10706));
    CascadeMux I__1631 (
            .O(N__10706),
            .I(N__10703));
    CascadeBuf I__1630 (
            .O(N__10703),
            .I(N__10700));
    CascadeMux I__1629 (
            .O(N__10700),
            .I(N__10697));
    CascadeBuf I__1628 (
            .O(N__10697),
            .I(N__10694));
    CascadeMux I__1627 (
            .O(N__10694),
            .I(N__10691));
    InMux I__1626 (
            .O(N__10691),
            .I(N__10688));
    LocalMux I__1625 (
            .O(N__10688),
            .I(N__10685));
    Span4Mux_v I__1624 (
            .O(N__10685),
            .I(N__10682));
    Sp12to4 I__1623 (
            .O(N__10682),
            .I(N__10679));
    Span12Mux_h I__1622 (
            .O(N__10679),
            .I(N__10676));
    Odrv12 I__1621 (
            .O(N__10676),
            .I(M_this_vga_signals_address_0));
    InMux I__1620 (
            .O(N__10673),
            .I(N__10667));
    InMux I__1619 (
            .O(N__10672),
            .I(N__10662));
    InMux I__1618 (
            .O(N__10671),
            .I(N__10662));
    InMux I__1617 (
            .O(N__10670),
            .I(N__10659));
    LocalMux I__1616 (
            .O(N__10667),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0 ));
    LocalMux I__1615 (
            .O(N__10662),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0 ));
    LocalMux I__1614 (
            .O(N__10659),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0 ));
    InMux I__1613 (
            .O(N__10652),
            .I(N__10644));
    InMux I__1612 (
            .O(N__10651),
            .I(N__10641));
    InMux I__1611 (
            .O(N__10650),
            .I(N__10634));
    InMux I__1610 (
            .O(N__10649),
            .I(N__10634));
    InMux I__1609 (
            .O(N__10648),
            .I(N__10634));
    InMux I__1608 (
            .O(N__10647),
            .I(N__10631));
    LocalMux I__1607 (
            .O(N__10644),
            .I(\this_vga_signals.mult1_un82_sum_axb2_i ));
    LocalMux I__1606 (
            .O(N__10641),
            .I(\this_vga_signals.mult1_un82_sum_axb2_i ));
    LocalMux I__1605 (
            .O(N__10634),
            .I(\this_vga_signals.mult1_un82_sum_axb2_i ));
    LocalMux I__1604 (
            .O(N__10631),
            .I(\this_vga_signals.mult1_un82_sum_axb2_i ));
    CascadeMux I__1603 (
            .O(N__10622),
            .I(N__10619));
    InMux I__1602 (
            .O(N__10619),
            .I(N__10616));
    LocalMux I__1601 (
            .O(N__10616),
            .I(N__10613));
    Span4Mux_h I__1600 (
            .O(N__10613),
            .I(N__10606));
    InMux I__1599 (
            .O(N__10612),
            .I(N__10603));
    InMux I__1598 (
            .O(N__10611),
            .I(N__10600));
    InMux I__1597 (
            .O(N__10610),
            .I(N__10595));
    InMux I__1596 (
            .O(N__10609),
            .I(N__10595));
    Odrv4 I__1595 (
            .O(N__10606),
            .I(\this_vga_signals.mult1_un82_sum_ac0_1 ));
    LocalMux I__1594 (
            .O(N__10603),
            .I(\this_vga_signals.mult1_un82_sum_ac0_1 ));
    LocalMux I__1593 (
            .O(N__10600),
            .I(\this_vga_signals.mult1_un82_sum_ac0_1 ));
    LocalMux I__1592 (
            .O(N__10595),
            .I(\this_vga_signals.mult1_un82_sum_ac0_1 ));
    CascadeMux I__1591 (
            .O(N__10586),
            .I(N__10581));
    InMux I__1590 (
            .O(N__10585),
            .I(N__10577));
    InMux I__1589 (
            .O(N__10584),
            .I(N__10572));
    InMux I__1588 (
            .O(N__10581),
            .I(N__10572));
    InMux I__1587 (
            .O(N__10580),
            .I(N__10569));
    LocalMux I__1586 (
            .O(N__10577),
            .I(\this_vga_signals.mult1_un82_sum_ac0_3_0_0 ));
    LocalMux I__1585 (
            .O(N__10572),
            .I(\this_vga_signals.mult1_un82_sum_ac0_3_0_0 ));
    LocalMux I__1584 (
            .O(N__10569),
            .I(\this_vga_signals.mult1_un82_sum_ac0_3_0_0 ));
    CascadeMux I__1583 (
            .O(N__10562),
            .I(N__10559));
    CascadeBuf I__1582 (
            .O(N__10559),
            .I(N__10556));
    CascadeMux I__1581 (
            .O(N__10556),
            .I(N__10553));
    CascadeBuf I__1580 (
            .O(N__10553),
            .I(N__10550));
    CascadeMux I__1579 (
            .O(N__10550),
            .I(N__10547));
    CascadeBuf I__1578 (
            .O(N__10547),
            .I(N__10544));
    CascadeMux I__1577 (
            .O(N__10544),
            .I(N__10541));
    CascadeBuf I__1576 (
            .O(N__10541),
            .I(N__10538));
    CascadeMux I__1575 (
            .O(N__10538),
            .I(N__10535));
    CascadeBuf I__1574 (
            .O(N__10535),
            .I(N__10532));
    CascadeMux I__1573 (
            .O(N__10532),
            .I(N__10529));
    CascadeBuf I__1572 (
            .O(N__10529),
            .I(N__10526));
    CascadeMux I__1571 (
            .O(N__10526),
            .I(N__10523));
    CascadeBuf I__1570 (
            .O(N__10523),
            .I(N__10520));
    CascadeMux I__1569 (
            .O(N__10520),
            .I(N__10517));
    CascadeBuf I__1568 (
            .O(N__10517),
            .I(N__10514));
    CascadeMux I__1567 (
            .O(N__10514),
            .I(N__10511));
    CascadeBuf I__1566 (
            .O(N__10511),
            .I(N__10508));
    CascadeMux I__1565 (
            .O(N__10508),
            .I(N__10505));
    CascadeBuf I__1564 (
            .O(N__10505),
            .I(N__10502));
    CascadeMux I__1563 (
            .O(N__10502),
            .I(N__10499));
    CascadeBuf I__1562 (
            .O(N__10499),
            .I(N__10496));
    CascadeMux I__1561 (
            .O(N__10496),
            .I(N__10493));
    CascadeBuf I__1560 (
            .O(N__10493),
            .I(N__10490));
    CascadeMux I__1559 (
            .O(N__10490),
            .I(N__10487));
    CascadeBuf I__1558 (
            .O(N__10487),
            .I(N__10484));
    CascadeMux I__1557 (
            .O(N__10484),
            .I(N__10481));
    CascadeBuf I__1556 (
            .O(N__10481),
            .I(N__10478));
    CascadeMux I__1555 (
            .O(N__10478),
            .I(N__10475));
    CascadeBuf I__1554 (
            .O(N__10475),
            .I(N__10472));
    CascadeMux I__1553 (
            .O(N__10472),
            .I(N__10469));
    InMux I__1552 (
            .O(N__10469),
            .I(N__10466));
    LocalMux I__1551 (
            .O(N__10466),
            .I(N__10463));
    Span4Mux_v I__1550 (
            .O(N__10463),
            .I(N__10460));
    Span4Mux_v I__1549 (
            .O(N__10460),
            .I(N__10457));
    Sp12to4 I__1548 (
            .O(N__10457),
            .I(N__10454));
    Span12Mux_h I__1547 (
            .O(N__10454),
            .I(N__10451));
    Odrv12 I__1546 (
            .O(N__10451),
            .I(M_this_vga_signals_address_1));
    CascadeMux I__1545 (
            .O(N__10448),
            .I(N__10441));
    InMux I__1544 (
            .O(N__10447),
            .I(N__10436));
    InMux I__1543 (
            .O(N__10446),
            .I(N__10433));
    InMux I__1542 (
            .O(N__10445),
            .I(N__10428));
    InMux I__1541 (
            .O(N__10444),
            .I(N__10428));
    InMux I__1540 (
            .O(N__10441),
            .I(N__10421));
    InMux I__1539 (
            .O(N__10440),
            .I(N__10421));
    InMux I__1538 (
            .O(N__10439),
            .I(N__10421));
    LocalMux I__1537 (
            .O(N__10436),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_i ));
    LocalMux I__1536 (
            .O(N__10433),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_i ));
    LocalMux I__1535 (
            .O(N__10428),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_i ));
    LocalMux I__1534 (
            .O(N__10421),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_i ));
    InMux I__1533 (
            .O(N__10412),
            .I(N__10407));
    CascadeMux I__1532 (
            .O(N__10411),
            .I(N__10404));
    CascadeMux I__1531 (
            .O(N__10410),
            .I(N__10401));
    LocalMux I__1530 (
            .O(N__10407),
            .I(N__10393));
    InMux I__1529 (
            .O(N__10404),
            .I(N__10386));
    InMux I__1528 (
            .O(N__10401),
            .I(N__10386));
    InMux I__1527 (
            .O(N__10400),
            .I(N__10386));
    InMux I__1526 (
            .O(N__10399),
            .I(N__10377));
    InMux I__1525 (
            .O(N__10398),
            .I(N__10377));
    InMux I__1524 (
            .O(N__10397),
            .I(N__10377));
    InMux I__1523 (
            .O(N__10396),
            .I(N__10377));
    Odrv4 I__1522 (
            .O(N__10393),
            .I(\this_vga_signals.mult1_un75_sum_c3 ));
    LocalMux I__1521 (
            .O(N__10386),
            .I(\this_vga_signals.mult1_un75_sum_c3 ));
    LocalMux I__1520 (
            .O(N__10377),
            .I(\this_vga_signals.mult1_un75_sum_c3 ));
    CascadeMux I__1519 (
            .O(N__10370),
            .I(N__10367));
    CascadeBuf I__1518 (
            .O(N__10367),
            .I(N__10364));
    CascadeMux I__1517 (
            .O(N__10364),
            .I(N__10361));
    CascadeBuf I__1516 (
            .O(N__10361),
            .I(N__10358));
    CascadeMux I__1515 (
            .O(N__10358),
            .I(N__10355));
    CascadeBuf I__1514 (
            .O(N__10355),
            .I(N__10352));
    CascadeMux I__1513 (
            .O(N__10352),
            .I(N__10349));
    CascadeBuf I__1512 (
            .O(N__10349),
            .I(N__10346));
    CascadeMux I__1511 (
            .O(N__10346),
            .I(N__10343));
    CascadeBuf I__1510 (
            .O(N__10343),
            .I(N__10340));
    CascadeMux I__1509 (
            .O(N__10340),
            .I(N__10337));
    CascadeBuf I__1508 (
            .O(N__10337),
            .I(N__10334));
    CascadeMux I__1507 (
            .O(N__10334),
            .I(N__10331));
    CascadeBuf I__1506 (
            .O(N__10331),
            .I(N__10328));
    CascadeMux I__1505 (
            .O(N__10328),
            .I(N__10325));
    CascadeBuf I__1504 (
            .O(N__10325),
            .I(N__10322));
    CascadeMux I__1503 (
            .O(N__10322),
            .I(N__10319));
    CascadeBuf I__1502 (
            .O(N__10319),
            .I(N__10316));
    CascadeMux I__1501 (
            .O(N__10316),
            .I(N__10313));
    CascadeBuf I__1500 (
            .O(N__10313),
            .I(N__10310));
    CascadeMux I__1499 (
            .O(N__10310),
            .I(N__10307));
    CascadeBuf I__1498 (
            .O(N__10307),
            .I(N__10304));
    CascadeMux I__1497 (
            .O(N__10304),
            .I(N__10301));
    CascadeBuf I__1496 (
            .O(N__10301),
            .I(N__10298));
    CascadeMux I__1495 (
            .O(N__10298),
            .I(N__10295));
    CascadeBuf I__1494 (
            .O(N__10295),
            .I(N__10292));
    CascadeMux I__1493 (
            .O(N__10292),
            .I(N__10289));
    CascadeBuf I__1492 (
            .O(N__10289),
            .I(N__10286));
    CascadeMux I__1491 (
            .O(N__10286),
            .I(N__10283));
    CascadeBuf I__1490 (
            .O(N__10283),
            .I(N__10280));
    CascadeMux I__1489 (
            .O(N__10280),
            .I(N__10277));
    InMux I__1488 (
            .O(N__10277),
            .I(N__10274));
    LocalMux I__1487 (
            .O(N__10274),
            .I(N__10271));
    Span4Mux_h I__1486 (
            .O(N__10271),
            .I(N__10268));
    Sp12to4 I__1485 (
            .O(N__10268),
            .I(N__10265));
    Span12Mux_s9_v I__1484 (
            .O(N__10265),
            .I(N__10262));
    Odrv12 I__1483 (
            .O(N__10262),
            .I(M_this_vga_signals_address_2));
    InMux I__1482 (
            .O(N__10259),
            .I(N__10256));
    LocalMux I__1481 (
            .O(N__10256),
            .I(N__10252));
    CascadeMux I__1480 (
            .O(N__10255),
            .I(N__10247));
    Span4Mux_v I__1479 (
            .O(N__10252),
            .I(N__10243));
    InMux I__1478 (
            .O(N__10251),
            .I(N__10240));
    InMux I__1477 (
            .O(N__10250),
            .I(N__10237));
    InMux I__1476 (
            .O(N__10247),
            .I(N__10232));
    InMux I__1475 (
            .O(N__10246),
            .I(N__10232));
    Odrv4 I__1474 (
            .O(N__10243),
            .I(\this_vga_signals.mult1_un61_sum_ac0_1 ));
    LocalMux I__1473 (
            .O(N__10240),
            .I(\this_vga_signals.mult1_un61_sum_ac0_1 ));
    LocalMux I__1472 (
            .O(N__10237),
            .I(\this_vga_signals.mult1_un61_sum_ac0_1 ));
    LocalMux I__1471 (
            .O(N__10232),
            .I(\this_vga_signals.mult1_un61_sum_ac0_1 ));
    InMux I__1470 (
            .O(N__10223),
            .I(N__10216));
    InMux I__1469 (
            .O(N__10222),
            .I(N__10212));
    InMux I__1468 (
            .O(N__10221),
            .I(N__10209));
    InMux I__1467 (
            .O(N__10220),
            .I(N__10203));
    InMux I__1466 (
            .O(N__10219),
            .I(N__10203));
    LocalMux I__1465 (
            .O(N__10216),
            .I(N__10196));
    InMux I__1464 (
            .O(N__10215),
            .I(N__10193));
    LocalMux I__1463 (
            .O(N__10212),
            .I(N__10190));
    LocalMux I__1462 (
            .O(N__10209),
            .I(N__10187));
    InMux I__1461 (
            .O(N__10208),
            .I(N__10184));
    LocalMux I__1460 (
            .O(N__10203),
            .I(N__10181));
    InMux I__1459 (
            .O(N__10202),
            .I(N__10178));
    InMux I__1458 (
            .O(N__10201),
            .I(N__10175));
    CascadeMux I__1457 (
            .O(N__10200),
            .I(N__10172));
    InMux I__1456 (
            .O(N__10199),
            .I(N__10165));
    Span4Mux_v I__1455 (
            .O(N__10196),
            .I(N__10154));
    LocalMux I__1454 (
            .O(N__10193),
            .I(N__10154));
    Span4Mux_v I__1453 (
            .O(N__10190),
            .I(N__10141));
    Span4Mux_v I__1452 (
            .O(N__10187),
            .I(N__10141));
    LocalMux I__1451 (
            .O(N__10184),
            .I(N__10141));
    Span4Mux_h I__1450 (
            .O(N__10181),
            .I(N__10141));
    LocalMux I__1449 (
            .O(N__10178),
            .I(N__10141));
    LocalMux I__1448 (
            .O(N__10175),
            .I(N__10141));
    InMux I__1447 (
            .O(N__10172),
            .I(N__10136));
    InMux I__1446 (
            .O(N__10171),
            .I(N__10136));
    InMux I__1445 (
            .O(N__10170),
            .I(N__10129));
    InMux I__1444 (
            .O(N__10169),
            .I(N__10129));
    InMux I__1443 (
            .O(N__10168),
            .I(N__10129));
    LocalMux I__1442 (
            .O(N__10165),
            .I(N__10126));
    InMux I__1441 (
            .O(N__10164),
            .I(N__10123));
    InMux I__1440 (
            .O(N__10163),
            .I(N__10120));
    InMux I__1439 (
            .O(N__10162),
            .I(N__10111));
    InMux I__1438 (
            .O(N__10161),
            .I(N__10111));
    InMux I__1437 (
            .O(N__10160),
            .I(N__10111));
    InMux I__1436 (
            .O(N__10159),
            .I(N__10111));
    Odrv4 I__1435 (
            .O(N__10154),
            .I(\this_vga_signals.mult1_un54_sum_i_0_3 ));
    Odrv4 I__1434 (
            .O(N__10141),
            .I(\this_vga_signals.mult1_un54_sum_i_0_3 ));
    LocalMux I__1433 (
            .O(N__10136),
            .I(\this_vga_signals.mult1_un54_sum_i_0_3 ));
    LocalMux I__1432 (
            .O(N__10129),
            .I(\this_vga_signals.mult1_un54_sum_i_0_3 ));
    Odrv4 I__1431 (
            .O(N__10126),
            .I(\this_vga_signals.mult1_un54_sum_i_0_3 ));
    LocalMux I__1430 (
            .O(N__10123),
            .I(\this_vga_signals.mult1_un54_sum_i_0_3 ));
    LocalMux I__1429 (
            .O(N__10120),
            .I(\this_vga_signals.mult1_un54_sum_i_0_3 ));
    LocalMux I__1428 (
            .O(N__10111),
            .I(\this_vga_signals.mult1_un54_sum_i_0_3 ));
    CascadeMux I__1427 (
            .O(N__10094),
            .I(N__10090));
    InMux I__1426 (
            .O(N__10093),
            .I(N__10087));
    InMux I__1425 (
            .O(N__10090),
            .I(N__10083));
    LocalMux I__1424 (
            .O(N__10087),
            .I(N__10080));
    InMux I__1423 (
            .O(N__10086),
            .I(N__10077));
    LocalMux I__1422 (
            .O(N__10083),
            .I(N__10074));
    Span4Mux_v I__1421 (
            .O(N__10080),
            .I(N__10071));
    LocalMux I__1420 (
            .O(N__10077),
            .I(N__10068));
    Odrv12 I__1419 (
            .O(N__10074),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c ));
    Odrv4 I__1418 (
            .O(N__10071),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c ));
    Odrv4 I__1417 (
            .O(N__10068),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c ));
    InMux I__1416 (
            .O(N__10061),
            .I(N__10057));
    InMux I__1415 (
            .O(N__10060),
            .I(N__10046));
    LocalMux I__1414 (
            .O(N__10057),
            .I(N__10043));
    InMux I__1413 (
            .O(N__10056),
            .I(N__10034));
    InMux I__1412 (
            .O(N__10055),
            .I(N__10034));
    InMux I__1411 (
            .O(N__10054),
            .I(N__10034));
    InMux I__1410 (
            .O(N__10053),
            .I(N__10034));
    InMux I__1409 (
            .O(N__10052),
            .I(N__10029));
    CascadeMux I__1408 (
            .O(N__10051),
            .I(N__10023));
    InMux I__1407 (
            .O(N__10050),
            .I(N__10020));
    InMux I__1406 (
            .O(N__10049),
            .I(N__10017));
    LocalMux I__1405 (
            .O(N__10046),
            .I(N__10014));
    Span4Mux_v I__1404 (
            .O(N__10043),
            .I(N__10009));
    LocalMux I__1403 (
            .O(N__10034),
            .I(N__10009));
    InMux I__1402 (
            .O(N__10033),
            .I(N__10004));
    InMux I__1401 (
            .O(N__10032),
            .I(N__10004));
    LocalMux I__1400 (
            .O(N__10029),
            .I(N__10001));
    InMux I__1399 (
            .O(N__10028),
            .I(N__9996));
    InMux I__1398 (
            .O(N__10027),
            .I(N__9996));
    InMux I__1397 (
            .O(N__10026),
            .I(N__9991));
    InMux I__1396 (
            .O(N__10023),
            .I(N__9991));
    LocalMux I__1395 (
            .O(N__10020),
            .I(\this_vga_signals.mult1_un54_sum_m_ns_1 ));
    LocalMux I__1394 (
            .O(N__10017),
            .I(\this_vga_signals.mult1_un54_sum_m_ns_1 ));
    Odrv4 I__1393 (
            .O(N__10014),
            .I(\this_vga_signals.mult1_un54_sum_m_ns_1 ));
    Odrv4 I__1392 (
            .O(N__10009),
            .I(\this_vga_signals.mult1_un54_sum_m_ns_1 ));
    LocalMux I__1391 (
            .O(N__10004),
            .I(\this_vga_signals.mult1_un54_sum_m_ns_1 ));
    Odrv4 I__1390 (
            .O(N__10001),
            .I(\this_vga_signals.mult1_un54_sum_m_ns_1 ));
    LocalMux I__1389 (
            .O(N__9996),
            .I(\this_vga_signals.mult1_un54_sum_m_ns_1 ));
    LocalMux I__1388 (
            .O(N__9991),
            .I(\this_vga_signals.mult1_un54_sum_m_ns_1 ));
    CascadeMux I__1387 (
            .O(N__9974),
            .I(N__9971));
    CascadeBuf I__1386 (
            .O(N__9971),
            .I(N__9968));
    CascadeMux I__1385 (
            .O(N__9968),
            .I(N__9965));
    CascadeBuf I__1384 (
            .O(N__9965),
            .I(N__9962));
    CascadeMux I__1383 (
            .O(N__9962),
            .I(N__9959));
    CascadeBuf I__1382 (
            .O(N__9959),
            .I(N__9956));
    CascadeMux I__1381 (
            .O(N__9956),
            .I(N__9953));
    CascadeBuf I__1380 (
            .O(N__9953),
            .I(N__9950));
    CascadeMux I__1379 (
            .O(N__9950),
            .I(N__9947));
    CascadeBuf I__1378 (
            .O(N__9947),
            .I(N__9944));
    CascadeMux I__1377 (
            .O(N__9944),
            .I(N__9941));
    CascadeBuf I__1376 (
            .O(N__9941),
            .I(N__9938));
    CascadeMux I__1375 (
            .O(N__9938),
            .I(N__9935));
    CascadeBuf I__1374 (
            .O(N__9935),
            .I(N__9932));
    CascadeMux I__1373 (
            .O(N__9932),
            .I(N__9929));
    CascadeBuf I__1372 (
            .O(N__9929),
            .I(N__9926));
    CascadeMux I__1371 (
            .O(N__9926),
            .I(N__9923));
    CascadeBuf I__1370 (
            .O(N__9923),
            .I(N__9920));
    CascadeMux I__1369 (
            .O(N__9920),
            .I(N__9917));
    CascadeBuf I__1368 (
            .O(N__9917),
            .I(N__9914));
    CascadeMux I__1367 (
            .O(N__9914),
            .I(N__9911));
    CascadeBuf I__1366 (
            .O(N__9911),
            .I(N__9908));
    CascadeMux I__1365 (
            .O(N__9908),
            .I(N__9905));
    CascadeBuf I__1364 (
            .O(N__9905),
            .I(N__9902));
    CascadeMux I__1363 (
            .O(N__9902),
            .I(N__9899));
    CascadeBuf I__1362 (
            .O(N__9899),
            .I(N__9896));
    CascadeMux I__1361 (
            .O(N__9896),
            .I(N__9893));
    CascadeBuf I__1360 (
            .O(N__9893),
            .I(N__9890));
    CascadeMux I__1359 (
            .O(N__9890),
            .I(N__9887));
    CascadeBuf I__1358 (
            .O(N__9887),
            .I(N__9884));
    CascadeMux I__1357 (
            .O(N__9884),
            .I(N__9881));
    InMux I__1356 (
            .O(N__9881),
            .I(N__9878));
    LocalMux I__1355 (
            .O(N__9878),
            .I(N__9875));
    Span4Mux_v I__1354 (
            .O(N__9875),
            .I(N__9872));
    Span4Mux_h I__1353 (
            .O(N__9872),
            .I(N__9869));
    Sp12to4 I__1352 (
            .O(N__9869),
            .I(N__9866));
    Span12Mux_h I__1351 (
            .O(N__9866),
            .I(N__9863));
    Odrv12 I__1350 (
            .O(N__9863),
            .I(M_this_vga_signals_address_4));
    InMux I__1349 (
            .O(N__9860),
            .I(N__9855));
    CascadeMux I__1348 (
            .O(N__9859),
            .I(N__9851));
    CascadeMux I__1347 (
            .O(N__9858),
            .I(N__9847));
    LocalMux I__1346 (
            .O(N__9855),
            .I(N__9844));
    InMux I__1345 (
            .O(N__9854),
            .I(N__9841));
    InMux I__1344 (
            .O(N__9851),
            .I(N__9834));
    InMux I__1343 (
            .O(N__9850),
            .I(N__9834));
    InMux I__1342 (
            .O(N__9847),
            .I(N__9831));
    Span4Mux_v I__1341 (
            .O(N__9844),
            .I(N__9826));
    LocalMux I__1340 (
            .O(N__9841),
            .I(N__9826));
    InMux I__1339 (
            .O(N__9840),
            .I(N__9821));
    InMux I__1338 (
            .O(N__9839),
            .I(N__9821));
    LocalMux I__1337 (
            .O(N__9834),
            .I(N__9816));
    LocalMux I__1336 (
            .O(N__9831),
            .I(N__9816));
    Span4Mux_h I__1335 (
            .O(N__9826),
            .I(N__9813));
    LocalMux I__1334 (
            .O(N__9821),
            .I(\this_vga_signals.new_pixel_1 ));
    Odrv4 I__1333 (
            .O(N__9816),
            .I(\this_vga_signals.new_pixel_1 ));
    Odrv4 I__1332 (
            .O(N__9813),
            .I(\this_vga_signals.new_pixel_1 ));
    InMux I__1331 (
            .O(N__9806),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    InMux I__1330 (
            .O(N__9803),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    InMux I__1329 (
            .O(N__9800),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    CascadeMux I__1328 (
            .O(N__9797),
            .I(N__9787));
    CascadeMux I__1327 (
            .O(N__9796),
            .I(N__9782));
    InMux I__1326 (
            .O(N__9795),
            .I(N__9774));
    InMux I__1325 (
            .O(N__9794),
            .I(N__9774));
    InMux I__1324 (
            .O(N__9793),
            .I(N__9769));
    InMux I__1323 (
            .O(N__9792),
            .I(N__9769));
    InMux I__1322 (
            .O(N__9791),
            .I(N__9764));
    InMux I__1321 (
            .O(N__9790),
            .I(N__9764));
    InMux I__1320 (
            .O(N__9787),
            .I(N__9757));
    InMux I__1319 (
            .O(N__9786),
            .I(N__9757));
    InMux I__1318 (
            .O(N__9785),
            .I(N__9757));
    InMux I__1317 (
            .O(N__9782),
            .I(N__9752));
    InMux I__1316 (
            .O(N__9781),
            .I(N__9752));
    InMux I__1315 (
            .O(N__9780),
            .I(N__9749));
    InMux I__1314 (
            .O(N__9779),
            .I(N__9746));
    LocalMux I__1313 (
            .O(N__9774),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    LocalMux I__1312 (
            .O(N__9769),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    LocalMux I__1311 (
            .O(N__9764),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    LocalMux I__1310 (
            .O(N__9757),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    LocalMux I__1309 (
            .O(N__9752),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    LocalMux I__1308 (
            .O(N__9749),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    LocalMux I__1307 (
            .O(N__9746),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    InMux I__1306 (
            .O(N__9731),
            .I(N__9725));
    InMux I__1305 (
            .O(N__9730),
            .I(N__9725));
    LocalMux I__1304 (
            .O(N__9725),
            .I(\this_vga_signals.N_19 ));
    InMux I__1303 (
            .O(N__9722),
            .I(N__9718));
    InMux I__1302 (
            .O(N__9721),
            .I(N__9715));
    LocalMux I__1301 (
            .O(N__9718),
            .I(\this_vga_signals.mult1_un75_sum_ac0_3_0_1 ));
    LocalMux I__1300 (
            .O(N__9715),
            .I(\this_vga_signals.mult1_un75_sum_ac0_3_0_1 ));
    CascadeMux I__1299 (
            .O(N__9710),
            .I(\this_vga_signals.mult1_un75_sum_axb2_i_0_cascade_ ));
    InMux I__1298 (
            .O(N__9707),
            .I(N__9701));
    InMux I__1297 (
            .O(N__9706),
            .I(N__9701));
    LocalMux I__1296 (
            .O(N__9701),
            .I(\this_vga_signals.mult1_un75_sum_ac0_1_0 ));
    CascadeMux I__1295 (
            .O(N__9698),
            .I(\this_vga_signals.g0_i_x2_0_0_a2_3_cascade_ ));
    InMux I__1294 (
            .O(N__9695),
            .I(N__9689));
    InMux I__1293 (
            .O(N__9694),
            .I(N__9689));
    LocalMux I__1292 (
            .O(N__9689),
            .I(\this_vga_signals.mult1_un75_sum_c3_0_0 ));
    CascadeMux I__1291 (
            .O(N__9686),
            .I(\this_vga_signals.if_i4_mux_0_cascade_ ));
    InMux I__1290 (
            .O(N__9683),
            .I(N__9680));
    LocalMux I__1289 (
            .O(N__9680),
            .I(\this_vga_signals.g1_0_a2 ));
    CascadeMux I__1288 (
            .O(N__9677),
            .I(N__9674));
    InMux I__1287 (
            .O(N__9674),
            .I(N__9671));
    LocalMux I__1286 (
            .O(N__9671),
            .I(\this_vga_signals.g0_i_x2_0_0_a2_0 ));
    CascadeMux I__1285 (
            .O(N__9668),
            .I(N__9665));
    InMux I__1284 (
            .O(N__9665),
            .I(N__9662));
    LocalMux I__1283 (
            .O(N__9662),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0 ));
    InMux I__1282 (
            .O(N__9659),
            .I(N__9656));
    LocalMux I__1281 (
            .O(N__9656),
            .I(N__9652));
    InMux I__1280 (
            .O(N__9655),
            .I(N__9649));
    Odrv4 I__1279 (
            .O(N__9652),
            .I(\this_vga_signals.g1_1 ));
    LocalMux I__1278 (
            .O(N__9649),
            .I(\this_vga_signals.g1_1 ));
    InMux I__1277 (
            .O(N__9644),
            .I(N__9641));
    LocalMux I__1276 (
            .O(N__9641),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_0 ));
    CascadeMux I__1275 (
            .O(N__9638),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_0_cascade_ ));
    InMux I__1274 (
            .O(N__9635),
            .I(N__9628));
    InMux I__1273 (
            .O(N__9634),
            .I(N__9628));
    InMux I__1272 (
            .O(N__9633),
            .I(N__9625));
    LocalMux I__1271 (
            .O(N__9628),
            .I(\this_vga_signals.mult1_un68_sum_0_3 ));
    LocalMux I__1270 (
            .O(N__9625),
            .I(\this_vga_signals.mult1_un68_sum_0_3 ));
    InMux I__1269 (
            .O(N__9620),
            .I(N__9617));
    LocalMux I__1268 (
            .O(N__9617),
            .I(\this_vga_signals.g0_0_a2_4 ));
    InMux I__1267 (
            .O(N__9614),
            .I(N__9608));
    InMux I__1266 (
            .O(N__9613),
            .I(N__9608));
    LocalMux I__1265 (
            .O(N__9608),
            .I(N__9604));
    InMux I__1264 (
            .O(N__9607),
            .I(N__9601));
    Span4Mux_h I__1263 (
            .O(N__9604),
            .I(N__9598));
    LocalMux I__1262 (
            .O(N__9601),
            .I(\this_vga_signals.mult1_un89_sum_axbxc3_0 ));
    Odrv4 I__1261 (
            .O(N__9598),
            .I(\this_vga_signals.mult1_un89_sum_axbxc3_0 ));
    CascadeMux I__1260 (
            .O(N__9593),
            .I(N__9590));
    InMux I__1259 (
            .O(N__9590),
            .I(N__9583));
    InMux I__1258 (
            .O(N__9589),
            .I(N__9583));
    InMux I__1257 (
            .O(N__9588),
            .I(N__9578));
    LocalMux I__1256 (
            .O(N__9583),
            .I(N__9575));
    InMux I__1255 (
            .O(N__9582),
            .I(N__9570));
    InMux I__1254 (
            .O(N__9581),
            .I(N__9570));
    LocalMux I__1253 (
            .O(N__9578),
            .I(\this_vga_signals.mult1_un89_sum_c3 ));
    Odrv12 I__1252 (
            .O(N__9575),
            .I(\this_vga_signals.mult1_un89_sum_c3 ));
    LocalMux I__1251 (
            .O(N__9570),
            .I(\this_vga_signals.mult1_un89_sum_c3 ));
    InMux I__1250 (
            .O(N__9563),
            .I(N__9560));
    LocalMux I__1249 (
            .O(N__9560),
            .I(N__9555));
    InMux I__1248 (
            .O(N__9559),
            .I(N__9550));
    InMux I__1247 (
            .O(N__9558),
            .I(N__9550));
    Span4Mux_v I__1246 (
            .O(N__9555),
            .I(N__9544));
    LocalMux I__1245 (
            .O(N__9550),
            .I(N__9544));
    InMux I__1244 (
            .O(N__9549),
            .I(N__9541));
    Odrv4 I__1243 (
            .O(N__9544),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3 ));
    LocalMux I__1242 (
            .O(N__9541),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3 ));
    InMux I__1241 (
            .O(N__9536),
            .I(N__9533));
    LocalMux I__1240 (
            .O(N__9533),
            .I(N__9530));
    Span4Mux_v I__1239 (
            .O(N__9530),
            .I(N__9527));
    Odrv4 I__1238 (
            .O(N__9527),
            .I(\this_vga_signals.mult1_un75_sum_ac0_1_1 ));
    InMux I__1237 (
            .O(N__9524),
            .I(N__9521));
    LocalMux I__1236 (
            .O(N__9521),
            .I(\this_vga_signals.g0_13_N_4L5 ));
    CascadeMux I__1235 (
            .O(N__9518),
            .I(\this_vga_signals.mult1_un75_sum_ac0_1_1_cascade_ ));
    InMux I__1234 (
            .O(N__9515),
            .I(N__9512));
    LocalMux I__1233 (
            .O(N__9512),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_3 ));
    InMux I__1232 (
            .O(N__9509),
            .I(N__9503));
    InMux I__1231 (
            .O(N__9508),
            .I(N__9500));
    InMux I__1230 (
            .O(N__9507),
            .I(N__9495));
    InMux I__1229 (
            .O(N__9506),
            .I(N__9495));
    LocalMux I__1228 (
            .O(N__9503),
            .I(\this_vga_signals.mult1_un68_sum_1_3 ));
    LocalMux I__1227 (
            .O(N__9500),
            .I(\this_vga_signals.mult1_un68_sum_1_3 ));
    LocalMux I__1226 (
            .O(N__9495),
            .I(\this_vga_signals.mult1_un68_sum_1_3 ));
    InMux I__1225 (
            .O(N__9488),
            .I(N__9485));
    LocalMux I__1224 (
            .O(N__9485),
            .I(\this_vga_signals.mult1_un75_sum_axb2_i_1_0_0 ));
    InMux I__1223 (
            .O(N__9482),
            .I(N__9479));
    LocalMux I__1222 (
            .O(N__9479),
            .I(\this_vga_signals.g4 ));
    CascadeMux I__1221 (
            .O(N__9476),
            .I(\this_vga_signals.g0_0_2_cascade_ ));
    InMux I__1220 (
            .O(N__9473),
            .I(N__9470));
    LocalMux I__1219 (
            .O(N__9470),
            .I(\this_vga_signals.g1_1_1_0_0 ));
    CascadeMux I__1218 (
            .O(N__9467),
            .I(N__9463));
    InMux I__1217 (
            .O(N__9466),
            .I(N__9458));
    InMux I__1216 (
            .O(N__9463),
            .I(N__9458));
    LocalMux I__1215 (
            .O(N__9458),
            .I(N__9455));
    Odrv4 I__1214 (
            .O(N__9455),
            .I(\this_vga_signals.N_4_0_0 ));
    InMux I__1213 (
            .O(N__9452),
            .I(N__9449));
    LocalMux I__1212 (
            .O(N__9449),
            .I(N__9446));
    Odrv4 I__1211 (
            .O(N__9446),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0 ));
    CascadeMux I__1210 (
            .O(N__9443),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_cascade_ ));
    CascadeMux I__1209 (
            .O(N__9440),
            .I(\this_vga_signals.mult1_un68_sum_0_3_cascade_ ));
    InMux I__1208 (
            .O(N__9437),
            .I(N__9434));
    LocalMux I__1207 (
            .O(N__9434),
            .I(N__9431));
    Odrv4 I__1206 (
            .O(N__9431),
            .I(\this_vga_signals.g1_0_a2_0 ));
    InMux I__1205 (
            .O(N__9428),
            .I(N__9425));
    LocalMux I__1204 (
            .O(N__9425),
            .I(N__9421));
    CascadeMux I__1203 (
            .O(N__9424),
            .I(N__9418));
    Span4Mux_h I__1202 (
            .O(N__9421),
            .I(N__9415));
    InMux I__1201 (
            .O(N__9418),
            .I(N__9412));
    Odrv4 I__1200 (
            .O(N__9415),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_6 ));
    LocalMux I__1199 (
            .O(N__9412),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_6 ));
    InMux I__1198 (
            .O(N__9407),
            .I(N__9404));
    LocalMux I__1197 (
            .O(N__9404),
            .I(N__9401));
    Odrv4 I__1196 (
            .O(N__9401),
            .I(\this_vga_signals.M_hcounter_q_fast_esr_RNI52HLZ0Z_9 ));
    InMux I__1195 (
            .O(N__9398),
            .I(N__9394));
    CascadeMux I__1194 (
            .O(N__9397),
            .I(N__9389));
    LocalMux I__1193 (
            .O(N__9394),
            .I(N__9386));
    InMux I__1192 (
            .O(N__9393),
            .I(N__9383));
    InMux I__1191 (
            .O(N__9392),
            .I(N__9378));
    InMux I__1190 (
            .O(N__9389),
            .I(N__9378));
    Odrv4 I__1189 (
            .O(N__9386),
            .I(\this_vga_signals.m8_0_1_0 ));
    LocalMux I__1188 (
            .O(N__9383),
            .I(\this_vga_signals.m8_0_1_0 ));
    LocalMux I__1187 (
            .O(N__9378),
            .I(\this_vga_signals.m8_0_1_0 ));
    InMux I__1186 (
            .O(N__9371),
            .I(N__9364));
    InMux I__1185 (
            .O(N__9370),
            .I(N__9359));
    InMux I__1184 (
            .O(N__9369),
            .I(N__9359));
    InMux I__1183 (
            .O(N__9368),
            .I(N__9352));
    InMux I__1182 (
            .O(N__9367),
            .I(N__9352));
    LocalMux I__1181 (
            .O(N__9364),
            .I(N__9347));
    LocalMux I__1180 (
            .O(N__9359),
            .I(N__9347));
    InMux I__1179 (
            .O(N__9358),
            .I(N__9342));
    InMux I__1178 (
            .O(N__9357),
            .I(N__9342));
    LocalMux I__1177 (
            .O(N__9352),
            .I(\this_vga_signals.M_hcounter_q_8_repZ0Z1 ));
    Odrv4 I__1176 (
            .O(N__9347),
            .I(\this_vga_signals.M_hcounter_q_8_repZ0Z1 ));
    LocalMux I__1175 (
            .O(N__9342),
            .I(\this_vga_signals.M_hcounter_q_8_repZ0Z1 ));
    InMux I__1174 (
            .O(N__9335),
            .I(N__9331));
    InMux I__1173 (
            .O(N__9334),
            .I(N__9328));
    LocalMux I__1172 (
            .O(N__9331),
            .I(\this_vga_signals.m8_0_3 ));
    LocalMux I__1171 (
            .O(N__9328),
            .I(\this_vga_signals.m8_0_3 ));
    InMux I__1170 (
            .O(N__9323),
            .I(N__9320));
    LocalMux I__1169 (
            .O(N__9320),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_3 ));
    CascadeMux I__1168 (
            .O(N__9317),
            .I(N__9314));
    InMux I__1167 (
            .O(N__9314),
            .I(N__9311));
    LocalMux I__1166 (
            .O(N__9311),
            .I(\this_vga_signals.g1_1_0_0 ));
    InMux I__1165 (
            .O(N__9308),
            .I(N__9305));
    LocalMux I__1164 (
            .O(N__9305),
            .I(N__9302));
    Span4Mux_h I__1163 (
            .O(N__9302),
            .I(N__9299));
    Odrv4 I__1162 (
            .O(N__9299),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_2_0 ));
    CascadeMux I__1161 (
            .O(N__9296),
            .I(\this_vga_signals.g1_0_0_cascade_ ));
    InMux I__1160 (
            .O(N__9293),
            .I(N__9290));
    LocalMux I__1159 (
            .O(N__9290),
            .I(\this_vga_signals.g1_6_0 ));
    InMux I__1158 (
            .O(N__9287),
            .I(N__9284));
    LocalMux I__1157 (
            .O(N__9284),
            .I(\this_vga_signals.g4_1 ));
    InMux I__1156 (
            .O(N__9281),
            .I(N__9278));
    LocalMux I__1155 (
            .O(N__9278),
            .I(N__9274));
    InMux I__1154 (
            .O(N__9277),
            .I(N__9268));
    Span4Mux_v I__1153 (
            .O(N__9274),
            .I(N__9265));
    InMux I__1152 (
            .O(N__9273),
            .I(N__9262));
    InMux I__1151 (
            .O(N__9272),
            .I(N__9257));
    InMux I__1150 (
            .O(N__9271),
            .I(N__9257));
    LocalMux I__1149 (
            .O(N__9268),
            .I(N__9254));
    Odrv4 I__1148 (
            .O(N__9265),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    LocalMux I__1147 (
            .O(N__9262),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    LocalMux I__1146 (
            .O(N__9257),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    Odrv4 I__1145 (
            .O(N__9254),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    InMux I__1144 (
            .O(N__9245),
            .I(N__9241));
    InMux I__1143 (
            .O(N__9244),
            .I(N__9238));
    LocalMux I__1142 (
            .O(N__9241),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_9 ));
    LocalMux I__1141 (
            .O(N__9238),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_9 ));
    CascadeMux I__1140 (
            .O(N__9233),
            .I(N__9228));
    CascadeMux I__1139 (
            .O(N__9232),
            .I(N__9225));
    CascadeMux I__1138 (
            .O(N__9231),
            .I(N__9219));
    InMux I__1137 (
            .O(N__9228),
            .I(N__9216));
    InMux I__1136 (
            .O(N__9225),
            .I(N__9213));
    InMux I__1135 (
            .O(N__9224),
            .I(N__9210));
    InMux I__1134 (
            .O(N__9223),
            .I(N__9207));
    InMux I__1133 (
            .O(N__9222),
            .I(N__9204));
    InMux I__1132 (
            .O(N__9219),
            .I(N__9201));
    LocalMux I__1131 (
            .O(N__9216),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_7 ));
    LocalMux I__1130 (
            .O(N__9213),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_7 ));
    LocalMux I__1129 (
            .O(N__9210),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_7 ));
    LocalMux I__1128 (
            .O(N__9207),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_7 ));
    LocalMux I__1127 (
            .O(N__9204),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_7 ));
    LocalMux I__1126 (
            .O(N__9201),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_7 ));
    CascadeMux I__1125 (
            .O(N__9188),
            .I(N__9182));
    InMux I__1124 (
            .O(N__9187),
            .I(N__9176));
    InMux I__1123 (
            .O(N__9186),
            .I(N__9171));
    InMux I__1122 (
            .O(N__9185),
            .I(N__9171));
    InMux I__1121 (
            .O(N__9182),
            .I(N__9168));
    InMux I__1120 (
            .O(N__9181),
            .I(N__9165));
    InMux I__1119 (
            .O(N__9180),
            .I(N__9162));
    InMux I__1118 (
            .O(N__9179),
            .I(N__9159));
    LocalMux I__1117 (
            .O(N__9176),
            .I(\this_vga_signals.M_hcounter_q_6_repZ0Z1 ));
    LocalMux I__1116 (
            .O(N__9171),
            .I(\this_vga_signals.M_hcounter_q_6_repZ0Z1 ));
    LocalMux I__1115 (
            .O(N__9168),
            .I(\this_vga_signals.M_hcounter_q_6_repZ0Z1 ));
    LocalMux I__1114 (
            .O(N__9165),
            .I(\this_vga_signals.M_hcounter_q_6_repZ0Z1 ));
    LocalMux I__1113 (
            .O(N__9162),
            .I(\this_vga_signals.M_hcounter_q_6_repZ0Z1 ));
    LocalMux I__1112 (
            .O(N__9159),
            .I(\this_vga_signals.M_hcounter_q_6_repZ0Z1 ));
    CascadeMux I__1111 (
            .O(N__9146),
            .I(N__9139));
    InMux I__1110 (
            .O(N__9145),
            .I(N__9136));
    InMux I__1109 (
            .O(N__9144),
            .I(N__9130));
    InMux I__1108 (
            .O(N__9143),
            .I(N__9125));
    InMux I__1107 (
            .O(N__9142),
            .I(N__9125));
    InMux I__1106 (
            .O(N__9139),
            .I(N__9122));
    LocalMux I__1105 (
            .O(N__9136),
            .I(N__9119));
    InMux I__1104 (
            .O(N__9135),
            .I(N__9114));
    InMux I__1103 (
            .O(N__9134),
            .I(N__9114));
    InMux I__1102 (
            .O(N__9133),
            .I(N__9111));
    LocalMux I__1101 (
            .O(N__9130),
            .I(\this_vga_signals.M_hcounter_q_9_repZ0Z1 ));
    LocalMux I__1100 (
            .O(N__9125),
            .I(\this_vga_signals.M_hcounter_q_9_repZ0Z1 ));
    LocalMux I__1099 (
            .O(N__9122),
            .I(\this_vga_signals.M_hcounter_q_9_repZ0Z1 ));
    Odrv4 I__1098 (
            .O(N__9119),
            .I(\this_vga_signals.M_hcounter_q_9_repZ0Z1 ));
    LocalMux I__1097 (
            .O(N__9114),
            .I(\this_vga_signals.M_hcounter_q_9_repZ0Z1 ));
    LocalMux I__1096 (
            .O(N__9111),
            .I(\this_vga_signals.M_hcounter_q_9_repZ0Z1 ));
    CascadeMux I__1095 (
            .O(N__9098),
            .I(\this_vga_signals.M_hcounter_q_fast_esr_RNIHH441Z0Z_5_cascade_ ));
    InMux I__1094 (
            .O(N__9095),
            .I(N__9092));
    LocalMux I__1093 (
            .O(N__9092),
            .I(\this_vga_signals.M_hcounter_q_fast_esr_RNIN6RRZ0Z_7 ));
    InMux I__1092 (
            .O(N__9089),
            .I(N__9086));
    LocalMux I__1091 (
            .O(N__9086),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_5 ));
    InMux I__1090 (
            .O(N__9083),
            .I(N__9080));
    LocalMux I__1089 (
            .O(N__9080),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_8 ));
    CEMux I__1088 (
            .O(N__9077),
            .I(N__9073));
    CEMux I__1087 (
            .O(N__9076),
            .I(N__9070));
    LocalMux I__1086 (
            .O(N__9073),
            .I(N__9063));
    LocalMux I__1085 (
            .O(N__9070),
            .I(N__9063));
    CEMux I__1084 (
            .O(N__9069),
            .I(N__9059));
    CEMux I__1083 (
            .O(N__9068),
            .I(N__9055));
    Span4Mux_v I__1082 (
            .O(N__9063),
            .I(N__9051));
    CEMux I__1081 (
            .O(N__9062),
            .I(N__9048));
    LocalMux I__1080 (
            .O(N__9059),
            .I(N__9045));
    CEMux I__1079 (
            .O(N__9058),
            .I(N__9042));
    LocalMux I__1078 (
            .O(N__9055),
            .I(N__9039));
    CEMux I__1077 (
            .O(N__9054),
            .I(N__9036));
    Span4Mux_h I__1076 (
            .O(N__9051),
            .I(N__9033));
    LocalMux I__1075 (
            .O(N__9048),
            .I(N__9030));
    Span4Mux_v I__1074 (
            .O(N__9045),
            .I(N__9023));
    LocalMux I__1073 (
            .O(N__9042),
            .I(N__9023));
    Span4Mux_v I__1072 (
            .O(N__9039),
            .I(N__9023));
    LocalMux I__1071 (
            .O(N__9036),
            .I(N__9020));
    Odrv4 I__1070 (
            .O(N__9033),
            .I(\this_vga_signals.N_550_1 ));
    Odrv4 I__1069 (
            .O(N__9030),
            .I(\this_vga_signals.N_550_1 ));
    Odrv4 I__1068 (
            .O(N__9023),
            .I(\this_vga_signals.N_550_1 ));
    Odrv4 I__1067 (
            .O(N__9020),
            .I(\this_vga_signals.N_550_1 ));
    InMux I__1066 (
            .O(N__9011),
            .I(N__9007));
    InMux I__1065 (
            .O(N__9010),
            .I(N__9002));
    LocalMux I__1064 (
            .O(N__9007),
            .I(N__8999));
    InMux I__1063 (
            .O(N__9006),
            .I(N__8996));
    InMux I__1062 (
            .O(N__9005),
            .I(N__8993));
    LocalMux I__1061 (
            .O(N__9002),
            .I(\this_vga_signals.m8_0_2 ));
    Odrv4 I__1060 (
            .O(N__8999),
            .I(\this_vga_signals.m8_0_2 ));
    LocalMux I__1059 (
            .O(N__8996),
            .I(\this_vga_signals.m8_0_2 ));
    LocalMux I__1058 (
            .O(N__8993),
            .I(\this_vga_signals.m8_0_2 ));
    InMux I__1057 (
            .O(N__8984),
            .I(N__8981));
    LocalMux I__1056 (
            .O(N__8981),
            .I(N__8978));
    Odrv4 I__1055 (
            .O(N__8978),
            .I(\this_vga_signals.g1_0_1 ));
    CascadeMux I__1054 (
            .O(N__8975),
            .I(\this_vga_signals.g4_1_1_cascade_ ));
    InMux I__1053 (
            .O(N__8972),
            .I(N__8967));
    InMux I__1052 (
            .O(N__8971),
            .I(N__8964));
    InMux I__1051 (
            .O(N__8970),
            .I(N__8961));
    LocalMux I__1050 (
            .O(N__8967),
            .I(\this_vga_signals.un1_haddress_0 ));
    LocalMux I__1049 (
            .O(N__8964),
            .I(\this_vga_signals.un1_haddress_0 ));
    LocalMux I__1048 (
            .O(N__8961),
            .I(\this_vga_signals.un1_haddress_0 ));
    CascadeMux I__1047 (
            .O(N__8954),
            .I(\this_vga_signals.mult1_un89_sum_axbxc3_0_cascade_ ));
    CascadeMux I__1046 (
            .O(N__8951),
            .I(N__8948));
    InMux I__1045 (
            .O(N__8948),
            .I(N__8945));
    LocalMux I__1044 (
            .O(N__8945),
            .I(\this_vga_signals.un1_haddress_0_cry_1_c_RNOZ0 ));
    CascadeMux I__1043 (
            .O(N__8942),
            .I(N__8939));
    InMux I__1042 (
            .O(N__8939),
            .I(N__8935));
    InMux I__1041 (
            .O(N__8938),
            .I(N__8932));
    LocalMux I__1040 (
            .O(N__8935),
            .I(N__8929));
    LocalMux I__1039 (
            .O(N__8932),
            .I(\this_vga_signals.m8_0_1_tz ));
    Odrv12 I__1038 (
            .O(N__8929),
            .I(\this_vga_signals.m8_0_1_tz ));
    InMux I__1037 (
            .O(N__8924),
            .I(N__8921));
    LocalMux I__1036 (
            .O(N__8921),
            .I(\this_vga_signals.ANC2_4_1 ));
    CascadeMux I__1035 (
            .O(N__8918),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2_cascade_ ));
    CascadeMux I__1034 (
            .O(N__8915),
            .I(N__8910));
    InMux I__1033 (
            .O(N__8914),
            .I(N__8907));
    CascadeMux I__1032 (
            .O(N__8913),
            .I(N__8904));
    InMux I__1031 (
            .O(N__8910),
            .I(N__8901));
    LocalMux I__1030 (
            .O(N__8907),
            .I(N__8898));
    InMux I__1029 (
            .O(N__8904),
            .I(N__8895));
    LocalMux I__1028 (
            .O(N__8901),
            .I(\this_vga_signals.M_hcounter_q_7_repZ0Z1 ));
    Odrv4 I__1027 (
            .O(N__8898),
            .I(\this_vga_signals.M_hcounter_q_7_repZ0Z1 ));
    LocalMux I__1026 (
            .O(N__8895),
            .I(\this_vga_signals.M_hcounter_q_7_repZ0Z1 ));
    InMux I__1025 (
            .O(N__8888),
            .I(N__8877));
    InMux I__1024 (
            .O(N__8887),
            .I(N__8877));
    InMux I__1023 (
            .O(N__8886),
            .I(N__8872));
    InMux I__1022 (
            .O(N__8885),
            .I(N__8872));
    InMux I__1021 (
            .O(N__8884),
            .I(N__8867));
    InMux I__1020 (
            .O(N__8883),
            .I(N__8867));
    InMux I__1019 (
            .O(N__8882),
            .I(N__8864));
    LocalMux I__1018 (
            .O(N__8877),
            .I(N__8861));
    LocalMux I__1017 (
            .O(N__8872),
            .I(\this_vga_signals.M_hcounter_q_5_repZ0Z1 ));
    LocalMux I__1016 (
            .O(N__8867),
            .I(\this_vga_signals.M_hcounter_q_5_repZ0Z1 ));
    LocalMux I__1015 (
            .O(N__8864),
            .I(\this_vga_signals.M_hcounter_q_5_repZ0Z1 ));
    Odrv4 I__1014 (
            .O(N__8861),
            .I(\this_vga_signals.M_hcounter_q_5_repZ0Z1 ));
    InMux I__1013 (
            .O(N__8852),
            .I(N__8846));
    InMux I__1012 (
            .O(N__8851),
            .I(N__8846));
    LocalMux I__1011 (
            .O(N__8846),
            .I(\this_vga_signals.mult1_un75_sum_axb1 ));
    CascadeMux I__1010 (
            .O(N__8843),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_i_cascade_ ));
    CascadeMux I__1009 (
            .O(N__8840),
            .I(\this_vga_signals.mult1_un82_sum_ac0_3_0_0_cascade_ ));
    CascadeMux I__1008 (
            .O(N__8837),
            .I(\this_vga_signals.new_pixel_1_axb_1_N_4L5_xZ0Z1_cascade_ ));
    InMux I__1007 (
            .O(N__8834),
            .I(N__8831));
    LocalMux I__1006 (
            .O(N__8831),
            .I(\this_vga_signals.M_hcounter_q_RNIPIQRNRZ0Z_2 ));
    InMux I__1005 (
            .O(N__8828),
            .I(N__8825));
    LocalMux I__1004 (
            .O(N__8825),
            .I(\this_vga_signals.M_hcounter_q_RNI5HOBQCZ0Z_1 ));
    CascadeMux I__1003 (
            .O(N__8822),
            .I(\this_vga_signals.M_hcounter_q_RNI8TTVN32Z0Z_2_cascade_ ));
    InMux I__1002 (
            .O(N__8819),
            .I(N__8816));
    LocalMux I__1001 (
            .O(N__8816),
            .I(N__8813));
    Span4Mux_h I__1000 (
            .O(N__8813),
            .I(N__8810));
    Odrv4 I__999 (
            .O(N__8810),
            .I(\this_vga_signals.new_pixel_1_axb_1 ));
    CascadeMux I__998 (
            .O(N__8807),
            .I(\this_vga_signals.N_510_cascade_ ));
    InMux I__997 (
            .O(N__8804),
            .I(N__8801));
    LocalMux I__996 (
            .O(N__8801),
            .I(N__8797));
    InMux I__995 (
            .O(N__8800),
            .I(N__8794));
    Odrv4 I__994 (
            .O(N__8797),
            .I(\this_vga_signals.un1_haddress_0_axb_6 ));
    LocalMux I__993 (
            .O(N__8794),
            .I(\this_vga_signals.un1_haddress_0_axb_6 ));
    CascadeMux I__992 (
            .O(N__8789),
            .I(\this_vga_signals.mult1_un75_sum_axb2_i_cascade_ ));
    InMux I__991 (
            .O(N__8786),
            .I(N__8781));
    InMux I__990 (
            .O(N__8785),
            .I(N__8778));
    InMux I__989 (
            .O(N__8784),
            .I(N__8771));
    LocalMux I__988 (
            .O(N__8781),
            .I(N__8766));
    LocalMux I__987 (
            .O(N__8778),
            .I(N__8766));
    InMux I__986 (
            .O(N__8777),
            .I(N__8763));
    InMux I__985 (
            .O(N__8776),
            .I(N__8758));
    InMux I__984 (
            .O(N__8775),
            .I(N__8758));
    InMux I__983 (
            .O(N__8774),
            .I(N__8755));
    LocalMux I__982 (
            .O(N__8771),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0 ));
    Odrv4 I__981 (
            .O(N__8766),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0 ));
    LocalMux I__980 (
            .O(N__8763),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0 ));
    LocalMux I__979 (
            .O(N__8758),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0 ));
    LocalMux I__978 (
            .O(N__8755),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0 ));
    InMux I__977 (
            .O(N__8744),
            .I(N__8741));
    LocalMux I__976 (
            .O(N__8741),
            .I(\this_vga_signals.mult1_un75_sum_ac0_3_0_1_x1 ));
    CascadeMux I__975 (
            .O(N__8738),
            .I(\this_vga_signals.mult1_un75_sum_ac0_3_0_1_x0_cascade_ ));
    InMux I__974 (
            .O(N__8735),
            .I(N__8729));
    InMux I__973 (
            .O(N__8734),
            .I(N__8729));
    LocalMux I__972 (
            .O(N__8729),
            .I(\this_vga_signals.mult1_un75_sum_ac0_1 ));
    CascadeMux I__971 (
            .O(N__8726),
            .I(\this_vga_signals.mult1_un75_sum_ac0_3_0_1_cascade_ ));
    InMux I__970 (
            .O(N__8723),
            .I(N__8720));
    LocalMux I__969 (
            .O(N__8720),
            .I(\this_vga_signals.mult1_un75_sum_axb2_i ));
    InMux I__968 (
            .O(N__8717),
            .I(N__8714));
    LocalMux I__967 (
            .O(N__8714),
            .I(\this_vga_signals.mult1_un75_sum_axbxc2 ));
    InMux I__966 (
            .O(N__8711),
            .I(N__8705));
    InMux I__965 (
            .O(N__8710),
            .I(N__8700));
    InMux I__964 (
            .O(N__8709),
            .I(N__8700));
    InMux I__963 (
            .O(N__8708),
            .I(N__8697));
    LocalMux I__962 (
            .O(N__8705),
            .I(\this_vga_signals.N_510_i ));
    LocalMux I__961 (
            .O(N__8700),
            .I(\this_vga_signals.N_510_i ));
    LocalMux I__960 (
            .O(N__8697),
            .I(\this_vga_signals.N_510_i ));
    CascadeMux I__959 (
            .O(N__8690),
            .I(N__8687));
    InMux I__958 (
            .O(N__8687),
            .I(N__8681));
    InMux I__957 (
            .O(N__8686),
            .I(N__8681));
    LocalMux I__956 (
            .O(N__8681),
            .I(N__8673));
    InMux I__955 (
            .O(N__8680),
            .I(N__8670));
    InMux I__954 (
            .O(N__8679),
            .I(N__8665));
    InMux I__953 (
            .O(N__8678),
            .I(N__8665));
    InMux I__952 (
            .O(N__8677),
            .I(N__8659));
    InMux I__951 (
            .O(N__8676),
            .I(N__8656));
    Span4Mux_v I__950 (
            .O(N__8673),
            .I(N__8649));
    LocalMux I__949 (
            .O(N__8670),
            .I(N__8649));
    LocalMux I__948 (
            .O(N__8665),
            .I(N__8649));
    InMux I__947 (
            .O(N__8664),
            .I(N__8642));
    InMux I__946 (
            .O(N__8663),
            .I(N__8642));
    InMux I__945 (
            .O(N__8662),
            .I(N__8642));
    LocalMux I__944 (
            .O(N__8659),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__943 (
            .O(N__8656),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    Odrv4 I__942 (
            .O(N__8649),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__941 (
            .O(N__8642),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    CascadeMux I__940 (
            .O(N__8633),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_cascade_ ));
    InMux I__939 (
            .O(N__8630),
            .I(N__8627));
    LocalMux I__938 (
            .O(N__8627),
            .I(\this_vga_signals.mult1_un75_sum_axb2_0_0 ));
    CascadeMux I__937 (
            .O(N__8624),
            .I(\this_vga_signals.mult1_un75_sum_axb2_0_0_cascade_ ));
    InMux I__936 (
            .O(N__8621),
            .I(N__8615));
    InMux I__935 (
            .O(N__8620),
            .I(N__8610));
    InMux I__934 (
            .O(N__8619),
            .I(N__8610));
    InMux I__933 (
            .O(N__8618),
            .I(N__8607));
    LocalMux I__932 (
            .O(N__8615),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5 ));
    LocalMux I__931 (
            .O(N__8610),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5 ));
    LocalMux I__930 (
            .O(N__8607),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5 ));
    CascadeMux I__929 (
            .O(N__8600),
            .I(N__8595));
    InMux I__928 (
            .O(N__8599),
            .I(N__8588));
    InMux I__927 (
            .O(N__8598),
            .I(N__8588));
    InMux I__926 (
            .O(N__8595),
            .I(N__8581));
    InMux I__925 (
            .O(N__8594),
            .I(N__8581));
    InMux I__924 (
            .O(N__8593),
            .I(N__8581));
    LocalMux I__923 (
            .O(N__8588),
            .I(\this_vga_signals.if_m2_0 ));
    LocalMux I__922 (
            .O(N__8581),
            .I(\this_vga_signals.if_m2_0 ));
    CascadeMux I__921 (
            .O(N__8576),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5_cascade_ ));
    InMux I__920 (
            .O(N__8573),
            .I(N__8570));
    LocalMux I__919 (
            .O(N__8570),
            .I(\this_vga_signals.g0_10_3_0_a2_0_0 ));
    InMux I__918 (
            .O(N__8567),
            .I(N__8564));
    LocalMux I__917 (
            .O(N__8564),
            .I(N__8561));
    Span4Mux_v I__916 (
            .O(N__8561),
            .I(N__8558));
    Odrv4 I__915 (
            .O(N__8558),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_1 ));
    InMux I__914 (
            .O(N__8555),
            .I(N__8551));
    InMux I__913 (
            .O(N__8554),
            .I(N__8548));
    LocalMux I__912 (
            .O(N__8551),
            .I(N__8545));
    LocalMux I__911 (
            .O(N__8548),
            .I(\this_vga_signals.g1_0 ));
    Odrv12 I__910 (
            .O(N__8545),
            .I(\this_vga_signals.g1_0 ));
    CascadeMux I__909 (
            .O(N__8540),
            .I(\this_vga_signals.g0_10_3_0_a2_0_0_cascade_ ));
    InMux I__908 (
            .O(N__8537),
            .I(N__8534));
    LocalMux I__907 (
            .O(N__8534),
            .I(\this_vga_signals.mult1_un75_sum_axb2_x0 ));
    CascadeMux I__906 (
            .O(N__8531),
            .I(N__8528));
    InMux I__905 (
            .O(N__8528),
            .I(N__8525));
    LocalMux I__904 (
            .O(N__8525),
            .I(\this_vga_signals.mult1_un75_sum_axb2_x1 ));
    CascadeMux I__903 (
            .O(N__8522),
            .I(\this_vga_signals.M_hcounter_q_7_rep1_esr_RNIJOMZ0Z71_cascade_ ));
    CascadeMux I__902 (
            .O(N__8519),
            .I(\this_vga_signals.m8_0_2_cascade_ ));
    CascadeMux I__901 (
            .O(N__8516),
            .I(\this_vga_signals.mult1_un61_sum_ac0_1_cascade_ ));
    CascadeMux I__900 (
            .O(N__8513),
            .I(\this_vga_signals.mult1_un54_sum_i_0_3_cascade_ ));
    CascadeMux I__899 (
            .O(N__8510),
            .I(\this_vga_signals.g1_6_0_cascade_ ));
    InMux I__898 (
            .O(N__8507),
            .I(N__8504));
    LocalMux I__897 (
            .O(N__8504),
            .I(N__8500));
    InMux I__896 (
            .O(N__8503),
            .I(N__8497));
    Odrv4 I__895 (
            .O(N__8500),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3 ));
    LocalMux I__894 (
            .O(N__8497),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3 ));
    InMux I__893 (
            .O(N__8492),
            .I(N__8489));
    LocalMux I__892 (
            .O(N__8489),
            .I(\this_vga_signals.g0_13_N_3L3_ns ));
    CascadeMux I__891 (
            .O(N__8486),
            .I(\this_vga_signals.g0_13_N_2L1_cascade_ ));
    CascadeMux I__890 (
            .O(N__8483),
            .I(\this_vga_signals.N_75_cascade_ ));
    InMux I__889 (
            .O(N__8480),
            .I(N__8477));
    LocalMux I__888 (
            .O(N__8477),
            .I(\this_vga_signals.mult1_un54_sum_m_1_1 ));
    CascadeMux I__887 (
            .O(N__8474),
            .I(\this_vga_signals.mult1_un54_sum_m_1_1_cascade_ ));
    InMux I__886 (
            .O(N__8471),
            .I(N__8468));
    LocalMux I__885 (
            .O(N__8468),
            .I(\this_vga_signals.N_75 ));
    CascadeMux I__884 (
            .O(N__8465),
            .I(\this_vga_signals.mult1_un54_sum_m_x0_1_cascade_ ));
    InMux I__883 (
            .O(N__8462),
            .I(N__8459));
    LocalMux I__882 (
            .O(N__8459),
            .I(\this_vga_signals.mult1_un54_sum_m_x1_1 ));
    InMux I__881 (
            .O(N__8456),
            .I(\this_vga_signals.un1_haddress_0_cry_5 ));
    InMux I__880 (
            .O(N__8453),
            .I(N__8449));
    CascadeMux I__879 (
            .O(N__8452),
            .I(N__8446));
    LocalMux I__878 (
            .O(N__8449),
            .I(N__8443));
    InMux I__877 (
            .O(N__8446),
            .I(N__8440));
    Odrv12 I__876 (
            .O(N__8443),
            .I(\this_vga_signals.un1_haddress_0_axb_7 ));
    LocalMux I__875 (
            .O(N__8440),
            .I(\this_vga_signals.un1_haddress_0_axb_7 ));
    InMux I__874 (
            .O(N__8435),
            .I(N__8432));
    LocalMux I__873 (
            .O(N__8432),
            .I(N__8429));
    Span4Mux_h I__872 (
            .O(N__8429),
            .I(N__8426));
    Odrv4 I__871 (
            .O(N__8426),
            .I(\this_vga_signals.un1_haddress_0_cry_6_c_RNI5KQUZ0 ));
    InMux I__870 (
            .O(N__8423),
            .I(\this_vga_signals.un1_haddress_0_cry_6 ));
    InMux I__869 (
            .O(N__8420),
            .I(N__8416));
    CascadeMux I__868 (
            .O(N__8419),
            .I(N__8413));
    LocalMux I__867 (
            .O(N__8416),
            .I(N__8410));
    InMux I__866 (
            .O(N__8413),
            .I(N__8407));
    Odrv4 I__865 (
            .O(N__8410),
            .I(\this_vga_signals.un1_haddress_0_cry_7_i ));
    LocalMux I__864 (
            .O(N__8407),
            .I(\this_vga_signals.un1_haddress_0_cry_7_i ));
    InMux I__863 (
            .O(N__8402),
            .I(\this_vga_signals.un1_haddress_0_cry_7 ));
    CascadeMux I__862 (
            .O(N__8399),
            .I(N__8396));
    InMux I__861 (
            .O(N__8396),
            .I(N__8393));
    LocalMux I__860 (
            .O(N__8393),
            .I(N__8390));
    Span4Mux_h I__859 (
            .O(N__8390),
            .I(N__8387));
    Odrv4 I__858 (
            .O(N__8387),
            .I(\this_vga_signals.un1_haddress_0_cry_7_c_RNIRVBSZ0Z7 ));
    CascadeMux I__857 (
            .O(N__8384),
            .I(\this_vga_signals.m8_0_1_tz_cascade_ ));
    CascadeMux I__856 (
            .O(N__8381),
            .I(\this_vga_signals.g1_cascade_ ));
    CascadeMux I__855 (
            .O(N__8378),
            .I(\this_vga_signals.g1_1_0_cascade_ ));
    CascadeMux I__854 (
            .O(N__8375),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIGF3C6Z0Z_9_cascade_ ));
    InMux I__853 (
            .O(N__8372),
            .I(N__8369));
    LocalMux I__852 (
            .O(N__8369),
            .I(N__8366));
    Span4Mux_h I__851 (
            .O(N__8366),
            .I(N__8363));
    Odrv4 I__850 (
            .O(N__8363),
            .I(\this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TAZ0Z7 ));
    InMux I__849 (
            .O(N__8360),
            .I(N__8357));
    LocalMux I__848 (
            .O(N__8357),
            .I(\this_vga_signals.mult1_un75_sum_i_0_3 ));
    CascadeMux I__847 (
            .O(N__8354),
            .I(N__8351));
    InMux I__846 (
            .O(N__8351),
            .I(N__8348));
    LocalMux I__845 (
            .O(N__8348),
            .I(\this_vga_signals.un1_haddress_0_axb_2_l_ofxZ0 ));
    InMux I__844 (
            .O(N__8345),
            .I(N__8342));
    LocalMux I__843 (
            .O(N__8342),
            .I(N__8339));
    Span4Mux_h I__842 (
            .O(N__8339),
            .I(N__8336));
    Odrv4 I__841 (
            .O(N__8336),
            .I(\this_vga_signals.un1_haddress_0_cry_1_c_RNIDP44VZ0Z02 ));
    InMux I__840 (
            .O(N__8333),
            .I(\this_vga_signals.un1_haddress_0_cry_1 ));
    InMux I__839 (
            .O(N__8330),
            .I(N__8327));
    LocalMux I__838 (
            .O(N__8327),
            .I(\this_vga_signals.un1_haddress_0_axb_3_l_fxZ0 ));
    CascadeMux I__837 (
            .O(N__8324),
            .I(N__8321));
    InMux I__836 (
            .O(N__8321),
            .I(N__8317));
    CascadeMux I__835 (
            .O(N__8320),
            .I(N__8314));
    LocalMux I__834 (
            .O(N__8317),
            .I(N__8311));
    InMux I__833 (
            .O(N__8314),
            .I(N__8308));
    Odrv4 I__832 (
            .O(N__8311),
            .I(\this_vga_signals.mult1_un68_sum_i_3 ));
    LocalMux I__831 (
            .O(N__8308),
            .I(\this_vga_signals.mult1_un68_sum_i_3 ));
    InMux I__830 (
            .O(N__8303),
            .I(N__8300));
    LocalMux I__829 (
            .O(N__8300),
            .I(N__8297));
    Span4Mux_v I__828 (
            .O(N__8297),
            .I(N__8294));
    Odrv4 I__827 (
            .O(N__8294),
            .I(\this_vga_signals.un1_haddress_0_cry_2_c_RNIVPNA9DZ0 ));
    InMux I__826 (
            .O(N__8291),
            .I(\this_vga_signals.un1_haddress_0_cry_2 ));
    CascadeMux I__825 (
            .O(N__8288),
            .I(N__8285));
    InMux I__824 (
            .O(N__8285),
            .I(N__8282));
    LocalMux I__823 (
            .O(N__8282),
            .I(N__8279));
    Odrv12 I__822 (
            .O(N__8279),
            .I(\this_vga_signals.un1_haddress_0_axb_4_l_fxZ0 ));
    InMux I__821 (
            .O(N__8276),
            .I(N__8273));
    LocalMux I__820 (
            .O(N__8273),
            .I(N__8270));
    Span4Mux_v I__819 (
            .O(N__8270),
            .I(N__8267));
    Odrv4 I__818 (
            .O(N__8267),
            .I(\this_vga_signals.un1_haddress_0_cry_3_c_RNIBO4TZ0Z72 ));
    InMux I__817 (
            .O(N__8264),
            .I(\this_vga_signals.un1_haddress_0_cry_3 ));
    InMux I__816 (
            .O(N__8261),
            .I(N__8258));
    LocalMux I__815 (
            .O(N__8258),
            .I(N__8255));
    Span4Mux_h I__814 (
            .O(N__8255),
            .I(N__8252));
    Odrv4 I__813 (
            .O(N__8252),
            .I(\this_vga_signals.un1_haddress_0_cry_4_c_RNI5SHJLZ0 ));
    InMux I__812 (
            .O(N__8249),
            .I(\this_vga_signals.un1_haddress_0_cry_4 ));
    CascadeMux I__811 (
            .O(N__8246),
            .I(N__8243));
    InMux I__810 (
            .O(N__8243),
            .I(N__8240));
    LocalMux I__809 (
            .O(N__8240),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIGF3C6Z0Z_9 ));
    InMux I__808 (
            .O(N__8237),
            .I(N__8231));
    InMux I__807 (
            .O(N__8236),
            .I(N__8231));
    LocalMux I__806 (
            .O(N__8231),
            .I(\this_vga_signals.un1_haddress_0_cry_5_THRU_CO ));
    CascadeMux I__805 (
            .O(N__8228),
            .I(\this_vga_signals.mult1_un75_sum_axb2_i_1_cascade_ ));
    InMux I__804 (
            .O(N__8225),
            .I(N__8222));
    LocalMux I__803 (
            .O(N__8222),
            .I(N__8219));
    Odrv12 I__802 (
            .O(N__8219),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_1 ));
    CascadeMux I__801 (
            .O(N__8216),
            .I(\this_vga_signals.N_4_i_1_cascade_ ));
    CascadeMux I__800 (
            .O(N__8213),
            .I(\this_vga_signals.mult1_un82_sum_ac0_1_cascade_ ));
    InMux I__799 (
            .O(N__8210),
            .I(N__8207));
    LocalMux I__798 (
            .O(N__8207),
            .I(\this_vga_signals.N_4_i ));
    CascadeMux I__797 (
            .O(N__8204),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_cascade_ ));
    CascadeMux I__796 (
            .O(N__8201),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_cascade_ ));
    CascadeMux I__795 (
            .O(N__8198),
            .I(N__8195));
    CascadeBuf I__794 (
            .O(N__8195),
            .I(N__8192));
    CascadeMux I__793 (
            .O(N__8192),
            .I(N__8189));
    CascadeBuf I__792 (
            .O(N__8189),
            .I(N__8186));
    CascadeMux I__791 (
            .O(N__8186),
            .I(N__8183));
    CascadeBuf I__790 (
            .O(N__8183),
            .I(N__8180));
    CascadeMux I__789 (
            .O(N__8180),
            .I(N__8177));
    CascadeBuf I__788 (
            .O(N__8177),
            .I(N__8174));
    CascadeMux I__787 (
            .O(N__8174),
            .I(N__8171));
    CascadeBuf I__786 (
            .O(N__8171),
            .I(N__8168));
    CascadeMux I__785 (
            .O(N__8168),
            .I(N__8165));
    CascadeBuf I__784 (
            .O(N__8165),
            .I(N__8162));
    CascadeMux I__783 (
            .O(N__8162),
            .I(N__8159));
    CascadeBuf I__782 (
            .O(N__8159),
            .I(N__8156));
    CascadeMux I__781 (
            .O(N__8156),
            .I(N__8153));
    CascadeBuf I__780 (
            .O(N__8153),
            .I(N__8150));
    CascadeMux I__779 (
            .O(N__8150),
            .I(N__8147));
    CascadeBuf I__778 (
            .O(N__8147),
            .I(N__8144));
    CascadeMux I__777 (
            .O(N__8144),
            .I(N__8141));
    CascadeBuf I__776 (
            .O(N__8141),
            .I(N__8138));
    CascadeMux I__775 (
            .O(N__8138),
            .I(N__8135));
    CascadeBuf I__774 (
            .O(N__8135),
            .I(N__8132));
    CascadeMux I__773 (
            .O(N__8132),
            .I(N__8129));
    CascadeBuf I__772 (
            .O(N__8129),
            .I(N__8126));
    CascadeMux I__771 (
            .O(N__8126),
            .I(N__8123));
    CascadeBuf I__770 (
            .O(N__8123),
            .I(N__8120));
    CascadeMux I__769 (
            .O(N__8120),
            .I(N__8117));
    CascadeBuf I__768 (
            .O(N__8117),
            .I(N__8114));
    CascadeMux I__767 (
            .O(N__8114),
            .I(N__8111));
    CascadeBuf I__766 (
            .O(N__8111),
            .I(N__8108));
    CascadeMux I__765 (
            .O(N__8108),
            .I(N__8105));
    InMux I__764 (
            .O(N__8105),
            .I(N__8102));
    LocalMux I__763 (
            .O(N__8102),
            .I(N__8099));
    Span12Mux_s10_h I__762 (
            .O(N__8099),
            .I(N__8096));
    Span12Mux_v I__761 (
            .O(N__8096),
            .I(N__8093));
    Span12Mux_h I__760 (
            .O(N__8093),
            .I(N__8090));
    Odrv12 I__759 (
            .O(N__8090),
            .I(M_this_vga_signals_address_3));
    CascadeMux I__758 (
            .O(N__8087),
            .I(\this_vga_signals.M_hcounter_d6lt9_cascade_ ));
    InMux I__757 (
            .O(N__8084),
            .I(N__8081));
    LocalMux I__756 (
            .O(N__8081),
            .I(N__8078));
    Span4Mux_v I__755 (
            .O(N__8078),
            .I(N__8073));
    InMux I__754 (
            .O(N__8077),
            .I(N__8068));
    InMux I__753 (
            .O(N__8076),
            .I(N__8068));
    Span4Mux_h I__752 (
            .O(N__8073),
            .I(N__8065));
    LocalMux I__751 (
            .O(N__8068),
            .I(this_pixel_clock_M_counter_q_i_1));
    Odrv4 I__750 (
            .O(N__8065),
            .I(this_pixel_clock_M_counter_q_i_1));
    InMux I__749 (
            .O(N__8060),
            .I(N__8055));
    InMux I__748 (
            .O(N__8059),
            .I(N__8049));
    InMux I__747 (
            .O(N__8058),
            .I(N__8049));
    LocalMux I__746 (
            .O(N__8055),
            .I(N__8046));
    InMux I__745 (
            .O(N__8054),
            .I(N__8043));
    LocalMux I__744 (
            .O(N__8049),
            .I(N__8040));
    Span4Mux_h I__743 (
            .O(N__8046),
            .I(N__8037));
    LocalMux I__742 (
            .O(N__8043),
            .I(this_pixel_clock_M_counter_q_0));
    Odrv4 I__741 (
            .O(N__8040),
            .I(this_pixel_clock_M_counter_q_0));
    Odrv4 I__740 (
            .O(N__8037),
            .I(this_pixel_clock_M_counter_q_0));
    CascadeMux I__739 (
            .O(N__8030),
            .I(\this_vga_signals.M_hcounter_d6_0_cascade_ ));
    IoInMux I__738 (
            .O(N__8027),
            .I(N__8024));
    LocalMux I__737 (
            .O(N__8024),
            .I(N__8021));
    IoSpan4Mux I__736 (
            .O(N__8021),
            .I(N__8018));
    Span4Mux_s2_h I__735 (
            .O(N__8018),
            .I(N__8015));
    Sp12to4 I__734 (
            .O(N__8015),
            .I(N__8012));
    Span12Mux_s5_h I__733 (
            .O(N__8012),
            .I(N__8009));
    Span12Mux_h I__732 (
            .O(N__8009),
            .I(N__8006));
    Odrv12 I__731 (
            .O(N__8006),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIUKG82Z0Z_9 ));
    CascadeMux I__730 (
            .O(N__8003),
            .I(\this_vga_signals.mult1_un75_sum_ac0_1_sx_cascade_ ));
    CascadeMux I__729 (
            .O(N__8000),
            .I(\this_vga_signals.if_m2_0_cascade_ ));
    CascadeMux I__728 (
            .O(N__7997),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_5_cascade_ ));
    CascadeMux I__727 (
            .O(N__7994),
            .I(\this_vga_signals.g0_13_N_3L3_x0_cascade_ ));
    InMux I__726 (
            .O(N__7991),
            .I(N__7987));
    InMux I__725 (
            .O(N__7990),
            .I(N__7984));
    LocalMux I__724 (
            .O(N__7987),
            .I(N__7981));
    LocalMux I__723 (
            .O(N__7984),
            .I(N__7978));
    Odrv4 I__722 (
            .O(N__7981),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_2_0_0 ));
    Odrv4 I__721 (
            .O(N__7978),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_2_0_0 ));
    InMux I__720 (
            .O(N__7973),
            .I(N__7970));
    LocalMux I__719 (
            .O(N__7970),
            .I(\this_vga_signals.g0_13_N_3L3_x1 ));
    CascadeMux I__718 (
            .O(N__7967),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_cascade_ ));
    InMux I__717 (
            .O(N__7964),
            .I(N__7961));
    LocalMux I__716 (
            .O(N__7961),
            .I(\this_vga_signals.M_hcounter_q_RNIUA42NDZ0Z_1 ));
    InMux I__715 (
            .O(N__7958),
            .I(N__7955));
    LocalMux I__714 (
            .O(N__7955),
            .I(\this_vga_signals.new_pixel_1_cry_0_c_RNOZ0 ));
    InMux I__713 (
            .O(N__7952),
            .I(N__7949));
    LocalMux I__712 (
            .O(N__7949),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIG53KZ0Z_9 ));
    CascadeMux I__711 (
            .O(N__7946),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_1_cascade_ ));
    CascadeMux I__710 (
            .O(N__7943),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_1_cascade_ ));
    CascadeMux I__709 (
            .O(N__7940),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_4_cascade_ ));
    IoInMux I__708 (
            .O(N__7937),
            .I(N__7934));
    LocalMux I__707 (
            .O(N__7934),
            .I(N__7931));
    IoSpan4Mux I__706 (
            .O(N__7931),
            .I(N__7928));
    Span4Mux_s1_v I__705 (
            .O(N__7928),
            .I(N__7925));
    Span4Mux_v I__704 (
            .O(N__7925),
            .I(N__7922));
    Odrv4 I__703 (
            .O(N__7922),
            .I(debug_c_i_1));
    CascadeMux I__702 (
            .O(N__7919),
            .I(N__7916));
    InMux I__701 (
            .O(N__7916),
            .I(N__7913));
    LocalMux I__700 (
            .O(N__7913),
            .I(\this_vga_signals.M_hcounter_q_esr_RNIG53K_1Z0Z_9 ));
    InMux I__699 (
            .O(N__7910),
            .I(N__7907));
    LocalMux I__698 (
            .O(N__7907),
            .I(\this_vga_signals.un3_hsynclt8_0 ));
    InMux I__697 (
            .O(N__7904),
            .I(N__7901));
    LocalMux I__696 (
            .O(N__7901),
            .I(N__7898));
    Odrv4 I__695 (
            .O(N__7898),
            .I(\this_vga_signals.new_pixel_1_i_0 ));
    InMux I__694 (
            .O(N__7895),
            .I(N__7892));
    LocalMux I__693 (
            .O(N__7892),
            .I(\this_vga_signals.new_pixel_1_5 ));
    InMux I__692 (
            .O(N__7889),
            .I(\this_vga_signals.new_pixel_1_cry_4 ));
    InMux I__691 (
            .O(N__7886),
            .I(N__7883));
    LocalMux I__690 (
            .O(N__7883),
            .I(\this_vga_signals.new_pixel_1_6 ));
    InMux I__689 (
            .O(N__7880),
            .I(\this_vga_signals.new_pixel_1_cry_5 ));
    CascadeMux I__688 (
            .O(N__7877),
            .I(N__7874));
    InMux I__687 (
            .O(N__7874),
            .I(N__7871));
    LocalMux I__686 (
            .O(N__7871),
            .I(\this_vga_signals.M_hcounter_q_i_7 ));
    InMux I__685 (
            .O(N__7868),
            .I(N__7865));
    LocalMux I__684 (
            .O(N__7865),
            .I(\this_vga_signals.new_pixel_1_7 ));
    InMux I__683 (
            .O(N__7862),
            .I(\this_vga_signals.new_pixel_1_cry_6 ));
    InMux I__682 (
            .O(N__7859),
            .I(N__7856));
    LocalMux I__681 (
            .O(N__7856),
            .I(\this_vga_signals.new_pixel_1_8 ));
    InMux I__680 (
            .O(N__7853),
            .I(bfn_6_22_0_));
    InMux I__679 (
            .O(N__7850),
            .I(N__7847));
    LocalMux I__678 (
            .O(N__7847),
            .I(\this_vga_signals.new_pixel_1_9 ));
    InMux I__677 (
            .O(N__7844),
            .I(\this_vga_signals.new_pixel_1_cry_8 ));
    InMux I__676 (
            .O(N__7841),
            .I(N__7838));
    LocalMux I__675 (
            .O(N__7838),
            .I(\this_vga_signals.new_pixel_1_10 ));
    InMux I__674 (
            .O(N__7835),
            .I(\this_vga_signals.new_pixel_1_cry_9 ));
    InMux I__673 (
            .O(N__7832),
            .I(\this_vga_signals.new_pixel_1_cry_10 ));
    InMux I__672 (
            .O(N__7829),
            .I(N__7826));
    LocalMux I__671 (
            .O(N__7826),
            .I(\this_vga_signals.new_pixel_1_11 ));
    InMux I__670 (
            .O(N__7823),
            .I(N__7820));
    LocalMux I__669 (
            .O(N__7820),
            .I(N__7817));
    Odrv12 I__668 (
            .O(N__7817),
            .I(\this_vga_signals.un4_hsynclt8_0 ));
    IoInMux I__667 (
            .O(N__7814),
            .I(N__7811));
    LocalMux I__666 (
            .O(N__7811),
            .I(N__7808));
    Span4Mux_s3_v I__665 (
            .O(N__7808),
            .I(N__7805));
    Span4Mux_h I__664 (
            .O(N__7805),
            .I(N__7802));
    Span4Mux_v I__663 (
            .O(N__7802),
            .I(N__7799));
    Odrv4 I__662 (
            .O(N__7799),
            .I(this_vga_signals_hsync_1_i));
    CascadeMux I__661 (
            .O(N__7796),
            .I(N_50_cascade_));
    IoInMux I__660 (
            .O(N__7793),
            .I(N__7790));
    LocalMux I__659 (
            .O(N__7790),
            .I(N__7787));
    Span4Mux_s0_v I__658 (
            .O(N__7787),
            .I(N__7784));
    Sp12to4 I__657 (
            .O(N__7784),
            .I(N__7781));
    Span12Mux_h I__656 (
            .O(N__7781),
            .I(N__7777));
    CascadeMux I__655 (
            .O(N__7780),
            .I(N__7771));
    Span12Mux_v I__654 (
            .O(N__7777),
            .I(N__7767));
    InMux I__653 (
            .O(N__7776),
            .I(N__7764));
    InMux I__652 (
            .O(N__7775),
            .I(N__7759));
    InMux I__651 (
            .O(N__7774),
            .I(N__7759));
    InMux I__650 (
            .O(N__7771),
            .I(N__7754));
    InMux I__649 (
            .O(N__7770),
            .I(N__7754));
    Odrv12 I__648 (
            .O(N__7767),
            .I(debug_c_0));
    LocalMux I__647 (
            .O(N__7764),
            .I(debug_c_0));
    LocalMux I__646 (
            .O(N__7759),
            .I(debug_c_0));
    LocalMux I__645 (
            .O(N__7754),
            .I(debug_c_0));
    IoInMux I__644 (
            .O(N__7745),
            .I(N__7742));
    LocalMux I__643 (
            .O(N__7742),
            .I(N__7739));
    IoSpan4Mux I__642 (
            .O(N__7739),
            .I(N__7735));
    InMux I__641 (
            .O(N__7738),
            .I(N__7732));
    Span4Mux_s3_h I__640 (
            .O(N__7735),
            .I(N__7727));
    LocalMux I__639 (
            .O(N__7732),
            .I(N__7727));
    Odrv4 I__638 (
            .O(N__7727),
            .I(rgb_c_2));
    InMux I__637 (
            .O(N__7724),
            .I(N__7716));
    InMux I__636 (
            .O(N__7723),
            .I(N__7713));
    InMux I__635 (
            .O(N__7722),
            .I(N__7708));
    InMux I__634 (
            .O(N__7721),
            .I(N__7708));
    InMux I__633 (
            .O(N__7720),
            .I(N__7703));
    InMux I__632 (
            .O(N__7719),
            .I(N__7703));
    LocalMux I__631 (
            .O(N__7716),
            .I(M_hcounter_q_esr_RNIH8GJ4_9));
    LocalMux I__630 (
            .O(N__7713),
            .I(M_hcounter_q_esr_RNIH8GJ4_9));
    LocalMux I__629 (
            .O(N__7708),
            .I(M_hcounter_q_esr_RNIH8GJ4_9));
    LocalMux I__628 (
            .O(N__7703),
            .I(M_hcounter_q_esr_RNIH8GJ4_9));
    InMux I__627 (
            .O(N__7694),
            .I(N__7691));
    LocalMux I__626 (
            .O(N__7691),
            .I(\this_vga_signals.new_pixel_1Z0Z_1 ));
    InMux I__625 (
            .O(N__7688),
            .I(\this_vga_signals.new_pixel_1_cry_0 ));
    InMux I__624 (
            .O(N__7685),
            .I(N__7682));
    LocalMux I__623 (
            .O(N__7682),
            .I(\this_vga_signals.new_pixel_1_2 ));
    InMux I__622 (
            .O(N__7679),
            .I(\this_vga_signals.new_pixel_1_cry_1 ));
    CascadeMux I__621 (
            .O(N__7676),
            .I(N__7673));
    InMux I__620 (
            .O(N__7673),
            .I(N__7670));
    LocalMux I__619 (
            .O(N__7670),
            .I(N__7667));
    Odrv4 I__618 (
            .O(N__7667),
            .I(\this_vga_signals.new_pixel_1_3 ));
    InMux I__617 (
            .O(N__7664),
            .I(\this_vga_signals.new_pixel_1_cry_2 ));
    InMux I__616 (
            .O(N__7661),
            .I(N__7658));
    LocalMux I__615 (
            .O(N__7658),
            .I(\this_vga_signals.new_pixel_1_4 ));
    InMux I__614 (
            .O(N__7655),
            .I(\this_vga_signals.new_pixel_1_cry_3 ));
    CascadeMux I__613 (
            .O(N__7652),
            .I(\this_vga_signals.new_pixel_1_1_cascade_ ));
    CascadeMux I__612 (
            .O(N__7649),
            .I(debug_c_0_cascade_));
    IoInMux I__611 (
            .O(N__7646),
            .I(N__7643));
    LocalMux I__610 (
            .O(N__7643),
            .I(N__7640));
    Span4Mux_s2_h I__609 (
            .O(N__7640),
            .I(N__7637));
    Span4Mux_v I__608 (
            .O(N__7637),
            .I(N__7633));
    InMux I__607 (
            .O(N__7636),
            .I(N__7630));
    Odrv4 I__606 (
            .O(N__7633),
            .I(rgb_c_3));
    LocalMux I__605 (
            .O(N__7630),
            .I(rgb_c_3));
    InMux I__604 (
            .O(N__7625),
            .I(N__7622));
    LocalMux I__603 (
            .O(N__7622),
            .I(N__7619));
    Odrv4 I__602 (
            .O(N__7619),
            .I(N_37));
    IoInMux I__601 (
            .O(N__7616),
            .I(N__7613));
    LocalMux I__600 (
            .O(N__7613),
            .I(N__7610));
    IoSpan4Mux I__599 (
            .O(N__7610),
            .I(N__7607));
    Span4Mux_s3_v I__598 (
            .O(N__7607),
            .I(N__7604));
    Span4Mux_v I__597 (
            .O(N__7604),
            .I(N__7600));
    CascadeMux I__596 (
            .O(N__7603),
            .I(N__7597));
    Span4Mux_v I__595 (
            .O(N__7600),
            .I(N__7594));
    InMux I__594 (
            .O(N__7597),
            .I(N__7591));
    Odrv4 I__593 (
            .O(N__7594),
            .I(rgb_c_4));
    LocalMux I__592 (
            .O(N__7591),
            .I(rgb_c_4));
    CascadeMux I__591 (
            .O(N__7586),
            .I(\this_vga_signals.new_pixel_1_3_1_cascade_ ));
    InMux I__590 (
            .O(N__7583),
            .I(N__7580));
    LocalMux I__589 (
            .O(N__7580),
            .I(\this_vga_signals.new_pixel_sx_0 ));
    IoInMux I__588 (
            .O(N__7577),
            .I(N__7574));
    LocalMux I__587 (
            .O(N__7574),
            .I(N__7571));
    Odrv12 I__586 (
            .O(N__7571),
            .I(this_vga_signals_vvisibility_i));
    InMux I__585 (
            .O(N__7568),
            .I(N__7565));
    LocalMux I__584 (
            .O(N__7565),
            .I(N_60));
    InMux I__583 (
            .O(N__7562),
            .I(N__7559));
    LocalMux I__582 (
            .O(N__7559),
            .I(N__7556));
    Odrv4 I__581 (
            .O(N__7556),
            .I(i7_mux));
    IoInMux I__580 (
            .O(N__7553),
            .I(N__7550));
    LocalMux I__579 (
            .O(N__7550),
            .I(N__7547));
    Span12Mux_s3_h I__578 (
            .O(N__7547),
            .I(N__7544));
    Odrv12 I__577 (
            .O(N__7544),
            .I(port_nmib_0_i));
    InMux I__576 (
            .O(N__7541),
            .I(N__7538));
    LocalMux I__575 (
            .O(N__7538),
            .I(N__7535));
    Odrv12 I__574 (
            .O(N__7535),
            .I(port_clk_c));
    InMux I__573 (
            .O(N__7532),
            .I(N__7529));
    LocalMux I__572 (
            .O(N__7529),
            .I(\this_delay_clk.M_pipe_qZ0Z_0 ));
    IoInMux I__571 (
            .O(N__7526),
            .I(N__7523));
    LocalMux I__570 (
            .O(N__7523),
            .I(N__7520));
    Span4Mux_s0_h I__569 (
            .O(N__7520),
            .I(N__7517));
    Span4Mux_h I__568 (
            .O(N__7517),
            .I(N__7514));
    Sp12to4 I__567 (
            .O(N__7514),
            .I(N__7511));
    Span12Mux_v I__566 (
            .O(N__7511),
            .I(N__7507));
    InMux I__565 (
            .O(N__7510),
            .I(N__7504));
    Odrv12 I__564 (
            .O(N__7507),
            .I(rgb_c_0));
    LocalMux I__563 (
            .O(N__7504),
            .I(rgb_c_0));
    InMux I__562 (
            .O(N__7499),
            .I(N__7496));
    LocalMux I__561 (
            .O(N__7496),
            .I(i7_mux_0));
    IoInMux I__560 (
            .O(N__7493),
            .I(N__7490));
    LocalMux I__559 (
            .O(N__7490),
            .I(N__7487));
    IoSpan4Mux I__558 (
            .O(N__7487),
            .I(N__7483));
    CascadeMux I__557 (
            .O(N__7486),
            .I(N__7480));
    Span4Mux_s2_h I__556 (
            .O(N__7483),
            .I(N__7477));
    InMux I__555 (
            .O(N__7480),
            .I(N__7474));
    Odrv4 I__554 (
            .O(N__7477),
            .I(rgb_c_1));
    LocalMux I__553 (
            .O(N__7474),
            .I(rgb_c_1));
    InMux I__552 (
            .O(N__7469),
            .I(N__7466));
    LocalMux I__551 (
            .O(N__7466),
            .I(N__7463));
    Odrv4 I__550 (
            .O(N__7463),
            .I(N_28_0));
    IoInMux I__549 (
            .O(N__7460),
            .I(N__7457));
    LocalMux I__548 (
            .O(N__7457),
            .I(N__7454));
    IoSpan4Mux I__547 (
            .O(N__7454),
            .I(N__7450));
    CascadeMux I__546 (
            .O(N__7453),
            .I(N__7447));
    IoSpan4Mux I__545 (
            .O(N__7450),
            .I(N__7444));
    InMux I__544 (
            .O(N__7447),
            .I(N__7441));
    Span4Mux_s3_h I__543 (
            .O(N__7444),
            .I(N__7438));
    LocalMux I__542 (
            .O(N__7441),
            .I(N__7435));
    Odrv4 I__541 (
            .O(N__7438),
            .I(rgb_c_5));
    Odrv4 I__540 (
            .O(N__7435),
            .I(rgb_c_5));
    IoInMux I__539 (
            .O(N__7430),
            .I(N__7427));
    LocalMux I__538 (
            .O(N__7427),
            .I(N_377_i));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_6_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_21_0_));
    defparam IN_MUX_bfv_6_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_22_0_ (
            .carryinitin(\this_vga_signals.new_pixel_1_cry_7 ),
            .carryinitout(bfn_6_22_0_));
    defparam IN_MUX_bfv_30_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_30_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_30_23_0_));
    defparam IN_MUX_bfv_30_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_30_24_0_ (
            .carryinitin(un1_M_this_external_address_q_cry_7),
            .carryinitout(bfn_30_24_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_20_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_21_0_));
    defparam IN_MUX_bfv_20_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_22_0_ (
            .carryinitin(un1_M_this_internal_address_q_cry_7),
            .carryinitout(bfn_20_22_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_16_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_24_0_ (
            .carryinitin(un1_M_this_data_count_q_cry_7),
            .carryinitout(bfn_16_24_0_));
    defparam IN_MUX_bfv_16_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_25_0_ (
            .carryinitin(un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO),
            .carryinitout(bfn_16_25_0_));
    ICE_GB \this_vga_signals.M_hcounter_q_esr_RNIUKG82_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__8027),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_583_g ));
    ICE_GB \this_reset_cond.M_stage_q_RNI6VB7_3  (
            .USERSIGNALTOGLOBALBUFFER(N__15770),
            .GLOBALBUFFEROUTPUT(M_this_state_q_nss_g_0));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_start_data_delay.N_377_i_LC_1_22_0 .C_ON=1'b0;
    defparam \this_start_data_delay.N_377_i_LC_1_22_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.N_377_i_LC_1_22_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \this_start_data_delay.N_377_i_LC_1_22_0  (
            .in0(N__14874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15907),
            .lcout(N_377_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNILC1D4_9_LC_4_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILC1D4_9_LC_4_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNILC1D4_9_LC_4_20_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNILC1D4_9_LC_4_20_3  (
            .in0(N__14878),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11988),
            .lcout(port_nmib_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_0_LC_4_20_4 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_0_LC_4_20_4 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_0_LC_4_20_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_delay_clk.M_pipe_q_0_LC_4_20_4  (
            .in0(N__7541),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21642),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_1_LC_4_20_6 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_1_LC_4_20_6 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_1_LC_4_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_1_LC_4_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7532),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21642),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.m27_LC_5_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.m27_LC_5_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.m27_LC_5_19_0 .LUT_INIT=16'b0001110100100101;
    LogicCell40 \this_vga_signals.m27_LC_5_19_0  (
            .in0(N__18460),
            .in1(N__17926),
            .in2(N__18417),
            .in3(N__18308),
            .lcout(N_28_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.m36_LC_5_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.m36_LC_5_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.m36_LC_5_19_4 .LUT_INIT=16'b0010110101110001;
    LogicCell40 \this_vga_signals.m36_LC_5_19_4  (
            .in0(N__18459),
            .in1(N__17925),
            .in2(N__18418),
            .in3(N__18309),
            .lcout(N_37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.m55_LC_5_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.m55_LC_5_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.m55_LC_5_19_7 .LUT_INIT=16'b0000001111101111;
    LogicCell40 \this_vga_signals.m55_LC_5_19_7  (
            .in0(N__18310),
            .in1(N__18461),
            .in2(N__17930),
            .in3(N__18412),
            .lcout(i7_mux_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_pixel_data_q_0_LC_5_20_1.C_ON=1'b0;
    defparam M_this_pixel_data_q_0_LC_5_20_1.SEQ_MODE=4'b1000;
    defparam M_this_pixel_data_q_0_LC_5_20_1.LUT_INIT=16'b0011001000000010;
    LogicCell40 M_this_pixel_data_q_0_LC_5_20_1 (
            .in0(N__7510),
            .in1(N__7720),
            .in2(N__7780),
            .in3(N__7568),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21639),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_pixel_data_q_1_LC_5_20_4.C_ON=1'b0;
    defparam M_this_pixel_data_q_1_LC_5_20_4.SEQ_MODE=4'b1000;
    defparam M_this_pixel_data_q_1_LC_5_20_4.LUT_INIT=16'b0001000101010000;
    LogicCell40 M_this_pixel_data_q_1_LC_5_20_4 (
            .in0(N__7719),
            .in1(N__7499),
            .in2(N__7486),
            .in3(N__7770),
            .lcout(rgb_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21639),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_pixel_data_q_5_LC_5_21_0.C_ON=1'b0;
    defparam M_this_pixel_data_q_5_LC_5_21_0.SEQ_MODE=4'b1000;
    defparam M_this_pixel_data_q_5_LC_5_21_0.LUT_INIT=16'b0001000101010000;
    LogicCell40 M_this_pixel_data_q_5_LC_5_21_0 (
            .in0(N__7722),
            .in1(N__7469),
            .in2(N__7453),
            .in3(N__7775),
            .lcout(rgb_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21643),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_2_c_RNIIU2M1G_LC_5_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.new_pixel_1_cry_2_c_RNIIU2M1G_LC_5_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_2_c_RNIIU2M1G_LC_5_21_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_2_c_RNIIU2M1G_LC_5_21_3  (
            .in0(N__7661),
            .in1(N__7859),
            .in2(N__7676),
            .in3(N__7850),
            .lcout(),
            .ltout(\this_vga_signals.new_pixel_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_9_c_RNIKG4BDR1_LC_5_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.new_pixel_1_cry_9_c_RNIKG4BDR1_LC_5_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_9_c_RNIKG4BDR1_LC_5_21_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_9_c_RNIKG4BDR1_LC_5_21_4  (
            .in0(N__7583),
            .in1(N__7841),
            .in2(N__7652),
            .in3(N__7829),
            .lcout(debug_c_0),
            .ltout(debug_c_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_pixel_data_q_3_LC_5_21_5.C_ON=1'b0;
    defparam M_this_pixel_data_q_3_LC_5_21_5.SEQ_MODE=4'b1000;
    defparam M_this_pixel_data_q_3_LC_5_21_5.LUT_INIT=16'b0000000001011100;
    LogicCell40 M_this_pixel_data_q_3_LC_5_21_5 (
            .in0(N__7562),
            .in1(N__7636),
            .in2(N__7649),
            .in3(N__7721),
            .lcout(rgb_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21643),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_pixel_data_q_4_LC_5_21_6.C_ON=1'b0;
    defparam M_this_pixel_data_q_4_LC_5_21_6.SEQ_MODE=4'b1000;
    defparam M_this_pixel_data_q_4_LC_5_21_6.LUT_INIT=16'b0001000100110000;
    LogicCell40 M_this_pixel_data_q_4_LC_5_21_6 (
            .in0(N__7625),
            .in1(N__7724),
            .in2(N__7603),
            .in3(N__7774),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21643),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_1_c_RNI7QR2DF2_LC_5_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.new_pixel_1_cry_1_c_RNI7QR2DF2_LC_5_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_1_c_RNI7QR2DF2_LC_5_22_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_1_c_RNI7QR2DF2_LC_5_22_1  (
            .in0(N__7694),
            .in1(N__7685),
            .in2(_gnd_net_),
            .in3(N__7895),
            .lcout(),
            .ltout(\this_vga_signals.new_pixel_1_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_5_c_RNIG1FT9B1_LC_5_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.new_pixel_1_cry_5_c_RNIG1FT9B1_LC_5_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_5_c_RNIG1FT9B1_LC_5_22_2 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_5_c_RNIG1FT9B1_LC_5_22_2  (
            .in0(N__7904),
            .in1(N__7886),
            .in2(N__7586),
            .in3(N__7868),
            .lcout(\this_vga_signals.new_pixel_sx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR31O3_0_9_LC_5_25_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR31O3_0_9_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR31O3_0_9_LC_5_25_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIR31O3_0_9_LC_5_25_3  (
            .in0(N__11993),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(this_vga_signals_vvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.m59_LC_6_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.m59_LC_6_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.m59_LC_6_19_3 .LUT_INIT=16'b0000111101010000;
    LogicCell40 \this_vga_signals.m59_LC_6_19_3  (
            .in0(N__17923),
            .in1(_gnd_net_),
            .in2(N__18467),
            .in3(N__18306),
            .lcout(N_60),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.m43_LC_6_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.m43_LC_6_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.m43_LC_6_19_4 .LUT_INIT=16'b0110000100110111;
    LogicCell40 \this_vga_signals.m43_LC_6_19_4  (
            .in0(N__18307),
            .in1(N__17922),
            .in2(N__18413),
            .in3(N__18462),
            .lcout(i7_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIFBM6_7_LC_6_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIFBM6_7_LC_6_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIFBM6_7_LC_6_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIFBM6_7_LC_6_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14111),
            .lcout(\this_vga_signals.M_hcounter_q_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUTFM_6_LC_6_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUTFM_6_LC_6_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUTFM_6_LC_6_20_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIUTFM_6_LC_6_20_3  (
            .in0(N__10931),
            .in1(N__14789),
            .in2(_gnd_net_),
            .in3(N__14606),
            .lcout(\this_vga_signals.un4_hsynclt8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.m49_LC_6_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.m49_LC_6_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.m49_LC_6_20_5 .LUT_INIT=16'b0000011101100111;
    LogicCell40 \this_vga_signals.m49_LC_6_20_5  (
            .in0(N__17924),
            .in1(N__18466),
            .in2(N__18419),
            .in3(N__18317),
            .lcout(),
            .ltout(N_50_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_pixel_data_q_2_LC_6_20_6.C_ON=1'b0;
    defparam M_this_pixel_data_q_2_LC_6_20_6.SEQ_MODE=4'b1000;
    defparam M_this_pixel_data_q_2_LC_6_20_6.LUT_INIT=16'b0000001100100010;
    LogicCell40 M_this_pixel_data_q_2_LC_6_20_6 (
            .in0(N__7738),
            .in1(N__7723),
            .in2(N__7796),
            .in3(N__7776),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21637),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIH8GJ4_9_LC_6_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIH8GJ4_9_LC_6_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIH8GJ4_9_LC_6_20_7 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIH8GJ4_9_LC_6_20_7  (
            .in0(N__11601),
            .in1(N__21390),
            .in2(_gnd_net_),
            .in3(N__11989),
            .lcout(M_hcounter_q_esr_RNIH8GJ4_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_0_c_LC_6_21_0 .C_ON=1'b1;
    defparam \this_vga_signals.new_pixel_1_cry_0_c_LC_6_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_0_c_LC_6_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_0_c_LC_6_21_0  (
            .in0(_gnd_net_),
            .in1(N__7958),
            .in2(N__9858),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_21_0_),
            .carryout(\this_vga_signals.new_pixel_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_0_c_RNIA47RND_LC_6_21_1 .C_ON=1'b1;
    defparam \this_vga_signals.new_pixel_1_cry_0_c_RNIA47RND_LC_6_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_0_c_RNIA47RND_LC_6_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_0_c_RNIA47RND_LC_6_21_1  (
            .in0(_gnd_net_),
            .in1(N__7964),
            .in2(N__11555),
            .in3(N__7688),
            .lcout(\this_vga_signals.new_pixel_1Z0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.new_pixel_1_cry_0 ),
            .carryout(\this_vga_signals.new_pixel_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_1_c_RNIRL8DV02_LC_6_21_2 .C_ON=1'b1;
    defparam \this_vga_signals.new_pixel_1_cry_1_c_RNIRL8DV02_LC_6_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_1_c_RNIRL8DV02_LC_6_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_1_c_RNIRL8DV02_LC_6_21_2  (
            .in0(_gnd_net_),
            .in1(N__8345),
            .in2(N__11480),
            .in3(N__7679),
            .lcout(\this_vga_signals.new_pixel_1_2 ),
            .ltout(),
            .carryin(\this_vga_signals.new_pixel_1_cry_1 ),
            .carryout(\this_vga_signals.new_pixel_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_2_c_RNIFPSJ9D_LC_6_21_3 .C_ON=1'b1;
    defparam \this_vga_signals.new_pixel_1_cry_2_c_RNIFPSJ9D_LC_6_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_2_c_RNIFPSJ9D_LC_6_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_2_c_RNIFPSJ9D_LC_6_21_3  (
            .in0(_gnd_net_),
            .in1(N__8303),
            .in2(N__11150),
            .in3(N__7664),
            .lcout(\this_vga_signals.new_pixel_1_3 ),
            .ltout(),
            .carryin(\this_vga_signals.new_pixel_1_cry_2 ),
            .carryout(\this_vga_signals.new_pixel_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_3_c_RNITQA682_LC_6_21_4 .C_ON=1'b1;
    defparam \this_vga_signals.new_pixel_1_cry_3_c_RNITQA682_LC_6_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_3_c_RNITQA682_LC_6_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_3_c_RNITQA682_LC_6_21_4  (
            .in0(_gnd_net_),
            .in1(N__8276),
            .in2(N__10997),
            .in3(N__7655),
            .lcout(\this_vga_signals.new_pixel_1_4 ),
            .ltout(),
            .carryin(\this_vga_signals.new_pixel_1_cry_3 ),
            .carryout(\this_vga_signals.new_pixel_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_4_c_RNI20CQL_LC_6_21_5 .C_ON=1'b1;
    defparam \this_vga_signals.new_pixel_1_cry_4_c_RNI20CQL_LC_6_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_4_c_RNI20CQL_LC_6_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_4_c_RNI20CQL_LC_6_21_5  (
            .in0(_gnd_net_),
            .in1(N__8261),
            .in2(N__14815),
            .in3(N__7889),
            .lcout(\this_vga_signals.new_pixel_1_5 ),
            .ltout(),
            .carryin(\this_vga_signals.new_pixel_1_cry_4 ),
            .carryout(\this_vga_signals.new_pixel_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_5_c_RNIJ8OH7_LC_6_21_6 .C_ON=1'b1;
    defparam \this_vga_signals.new_pixel_1_cry_5_c_RNIJ8OH7_LC_6_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_5_c_RNIJ8OH7_LC_6_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_5_c_RNIJ8OH7_LC_6_21_6  (
            .in0(_gnd_net_),
            .in1(N__8372),
            .in2(N__14607),
            .in3(N__7880),
            .lcout(\this_vga_signals.new_pixel_1_6 ),
            .ltout(),
            .carryin(\this_vga_signals.new_pixel_1_cry_5 ),
            .carryout(\this_vga_signals.new_pixel_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_6_c_RNI6UM51_LC_6_21_7 .C_ON=1'b1;
    defparam \this_vga_signals.new_pixel_1_cry_6_c_RNI6UM51_LC_6_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_6_c_RNI6UM51_LC_6_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_6_c_RNI6UM51_LC_6_21_7  (
            .in0(_gnd_net_),
            .in1(N__8435),
            .in2(N__7877),
            .in3(N__7862),
            .lcout(\this_vga_signals.new_pixel_1_7 ),
            .ltout(),
            .carryin(\this_vga_signals.new_pixel_1_cry_6 ),
            .carryout(\this_vga_signals.new_pixel_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_7_c_RNI22G7F_LC_6_22_0 .C_ON=1'b1;
    defparam \this_vga_signals.new_pixel_1_cry_7_c_RNI22G7F_LC_6_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_7_c_RNI22G7F_LC_6_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_7_c_RNI22G7F_LC_6_22_0  (
            .in0(_gnd_net_),
            .in1(N__8420),
            .in2(N__8399),
            .in3(N__7853),
            .lcout(\this_vga_signals.new_pixel_1_8 ),
            .ltout(),
            .carryin(bfn_6_22_0_),
            .carryout(\this_vga_signals.new_pixel_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_8_c_RNI48BK_LC_6_22_1 .C_ON=1'b1;
    defparam \this_vga_signals.new_pixel_1_cry_8_c_RNI48BK_LC_6_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_8_c_RNI48BK_LC_6_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_8_c_RNI48BK_LC_6_22_1  (
            .in0(_gnd_net_),
            .in1(N__7952),
            .in2(N__20356),
            .in3(N__7844),
            .lcout(\this_vga_signals.new_pixel_1_9 ),
            .ltout(),
            .carryin(\this_vga_signals.new_pixel_1_cry_8 ),
            .carryout(\this_vga_signals.new_pixel_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_9_c_RNI5ACK_LC_6_22_2 .C_ON=1'b1;
    defparam \this_vga_signals.new_pixel_1_cry_9_c_RNI5ACK_LC_6_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_9_c_RNI5ACK_LC_6_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_9_c_RNI5ACK_LC_6_22_2  (
            .in0(_gnd_net_),
            .in1(N__20312),
            .in2(N__7919),
            .in3(N__7835),
            .lcout(\this_vga_signals.new_pixel_1_10 ),
            .ltout(),
            .carryin(\this_vga_signals.new_pixel_1_cry_9 ),
            .carryout(\this_vga_signals.new_pixel_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_10_c_RNID6631_LC_6_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.new_pixel_1_cry_10_c_RNID6631_LC_6_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_10_c_RNID6631_LC_6_22_3 .LUT_INIT=16'b0000000111111110;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_10_c_RNID6631_LC_6_22_3  (
            .in0(N__14112),
            .in1(N__14298),
            .in2(N__14483),
            .in3(N__7832),
            .lcout(\this_vga_signals.new_pixel_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC1312_9_LC_6_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC1312_9_LC_6_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC1312_9_LC_6_22_4 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIC1312_9_LC_6_22_4  (
            .in0(N__7823),
            .in1(N__7910),
            .in2(N__14303),
            .in3(N__14476),
            .lcout(this_vga_signals_hsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_2_9_LC_6_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_2_9_LC_6_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_2_9_LC_6_24_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIG53K_2_9_LC_6_24_6  (
            .in0(N__11602),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(debug_c_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clock.M_counter_q_0_LC_7_19_0 .C_ON=1'b0;
    defparam \this_pixel_clock.M_counter_q_0_LC_7_19_0 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clock.M_counter_q_0_LC_7_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_pixel_clock.M_counter_q_0_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8054),
            .lcout(this_pixel_clock_M_counter_q_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21632),
            .ce(),
            .sr(N__21349));
    defparam \this_vga_signals.M_hcounter_q_0_LC_7_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_7_20_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_7_20_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(N__12853),
            .in2(_gnd_net_),
            .in3(N__9840),
            .lcout(\this_vga_signals.new_pixel_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21634),
            .ce(),
            .sr(N__11341));
    defparam \this_vga_signals.M_hcounter_q_1_LC_7_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_7_20_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_7_20_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_7_20_4  (
            .in0(N__9839),
            .in1(_gnd_net_),
            .in2(N__12883),
            .in3(N__11513),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21634),
            .ce(),
            .sr(N__11341));
    defparam \this_pixel_clock.M_counter_q_1_LC_7_21_1 .C_ON=1'b0;
    defparam \this_pixel_clock.M_counter_q_1_LC_7_21_1 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clock.M_counter_q_1_LC_7_21_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_pixel_clock.M_counter_q_1_LC_7_21_1  (
            .in0(N__8077),
            .in1(N__8059),
            .in2(_gnd_net_),
            .in3(N__21386),
            .lcout(this_pixel_clock_M_counter_q_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21638),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_1_9_LC_7_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_1_9_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_1_9_LC_7_21_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIG53K_1_9_LC_7_21_2  (
            .in0(N__14437),
            .in1(N__14283),
            .in2(_gnd_net_),
            .in3(N__14114),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNIG53K_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.G_296_LC_7_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.G_296_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.G_296_LC_7_21_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.G_296_LC_7_21_3  (
            .in0(N__8076),
            .in1(N__8058),
            .in2(_gnd_net_),
            .in3(N__21385),
            .lcout(\this_vga_signals.GZ0Z_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNID96T_6_LC_7_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNID96T_6_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNID96T_6_LC_7_21_4 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNID96T_6_LC_7_21_4  (
            .in0(N__14591),
            .in1(N__10996),
            .in2(N__14816),
            .in3(N__14115),
            .lcout(\this_vga_signals.un3_hsynclt8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIG043KR2_0_LC_7_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIG043KR2_0_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIG043KR2_0_LC_7_22_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIG043KR2_0_LC_7_22_0  (
            .in0(N__9559),
            .in1(N__9850),
            .in2(N__9593),
            .in3(N__9614),
            .lcout(\this_vga_signals.new_pixel_1_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIUA42ND_1_LC_7_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIUA42ND_1_LC_7_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIUA42ND_1_LC_7_22_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIUA42ND_1_LC_7_22_4  (
            .in0(N__11528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8819),
            .lcout(\this_vga_signals.M_hcounter_q_RNIUA42NDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_cry_0_c_RNO_LC_7_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.new_pixel_1_cry_0_c_RNO_LC_7_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_cry_0_c_RNO_LC_7_22_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.new_pixel_1_cry_0_c_RNO_LC_7_22_5  (
            .in0(N__9613),
            .in1(N__9589),
            .in2(N__9859),
            .in3(N__9558),
            .lcout(\this_vga_signals.new_pixel_1_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_9_LC_7_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_9_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_9_LC_7_22_6 .LUT_INIT=16'b1010101010011001;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIG53K_9_LC_7_22_6  (
            .in0(N__14470),
            .in1(N__14296),
            .in2(_gnd_net_),
            .in3(N__14113),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNIG53KZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_6_LC_9_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_6_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_6_LC_9_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_6_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11273),
            .lcout(\this_vga_signals.M_hcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21603),
            .ce(N__9062),
            .sr(N__11339));
    defparam \this_vga_signals.un4_haddress_g0_6_LC_9_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_6_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_6_LC_9_17_0 .LUT_INIT=16'b0110101111010111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_6_LC_9_17_0  (
            .in0(N__14198),
            .in1(N__14000),
            .in2(N__14397),
            .in3(N__14532),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_5_LC_9_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_5_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_5_LC_9_17_1 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_5_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7946),
            .in3(N__14750),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_2_LC_9_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_2_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_2_LC_9_17_2 .LUT_INIT=16'b0001000100010111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_2_LC_9_17_2  (
            .in0(N__11124),
            .in1(N__10974),
            .in2(N__7943),
            .in3(N__8554),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_9_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_9_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_9_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_9_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11180),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21613),
            .ce(N__9068),
            .sr(N__11336));
    defparam \this_vga_signals.un4_haddress_g0_25_LC_9_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_25_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_25_LC_9_17_4 .LUT_INIT=16'b0110101111010111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_25_LC_9_17_4  (
            .in0(N__14199),
            .in1(N__14001),
            .in2(N__14398),
            .in3(N__14533),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_23_LC_9_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_23_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_23_LC_9_17_5 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_23_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7940),
            .in3(N__14751),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHGHF3_9_LC_9_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHGHF3_9_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIHGHF3_9_LC_9_18_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIHGHF3_9_LC_9_18_1  (
            .in0(N__12895),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11345),
            .lcout(\this_vga_signals.N_550_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_30_LC_9_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_30_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_30_LC_9_18_4 .LUT_INIT=16'b0111100110011111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_30_LC_9_18_4  (
            .in0(N__13999),
            .in1(N__9144),
            .in2(N__14219),
            .in3(N__9187),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_28_LC_9_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_28_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_28_LC_9_18_5 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_28_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7997),
            .in3(N__14745),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_13_N_3L3_x0_LC_9_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_13_N_3L3_x0_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_13_N_3L3_x0_LC_9_19_0 .LUT_INIT=16'b1110000110100101;
    LogicCell40 \this_vga_signals.un4_haddress_g0_13_N_3L3_x0_LC_9_19_0  (
            .in0(N__7991),
            .in1(N__10161),
            .in2(N__10991),
            .in3(N__10032),
            .lcout(),
            .ltout(\this_vga_signals.g0_13_N_3L3_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_13_N_3L3_ns_LC_9_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_13_N_3L3_ns_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_13_N_3L3_ns_LC_9_19_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \this_vga_signals.un4_haddress_g0_13_N_3L3_ns_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__7973),
            .in2(N__7994),
            .in3(N__10246),
            .lcout(\this_vga_signals.g0_13_N_3L3_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_13_N_3L3_x1_LC_9_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_13_N_3L3_x1_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_13_N_3L3_x1_LC_9_19_2 .LUT_INIT=16'b1111000011100001;
    LogicCell40 \this_vga_signals.un4_haddress_g0_13_N_3L3_x1_LC_9_19_2  (
            .in0(N__10026),
            .in1(N__7990),
            .in2(N__10990),
            .in3(N__10160),
            .lcout(\this_vga_signals.g0_13_N_3L3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_9_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_9_19_4 .LUT_INIT=16'b0010110101001011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_9_19_4  (
            .in0(N__10965),
            .in1(N__14746),
            .in2(N__10051),
            .in3(N__10159),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_0 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_axb_4_l_fx_LC_9_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un1_haddress_0_axb_4_l_fx_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_axb_4_l_fx_LC_9_19_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un1_haddress_0_axb_4_l_fx_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__8677),
            .in2(N__7967),
            .in3(N__9794),
            .lcout(\this_vga_signals.un1_haddress_0_axb_4_l_fxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_9_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_9_19_6 .LUT_INIT=16'b0000000100010101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_9_19_6  (
            .in0(N__10093),
            .in1(N__10162),
            .in2(N__10255),
            .in3(N__10033),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_address_buffer_q_esr_3_LC_9_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_3_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_3_LC_9_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_3_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__8784),
            .in2(N__8201),
            .in3(N__9795),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21623),
            .ce(N__15307),
            .sr(N__15218));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIAV2K_6_LC_9_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIAV2K_6_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIAV2K_6_LC_9_20_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIAV2K_6_LC_9_20_0  (
            .in0(N__14741),
            .in1(N__14092),
            .in2(_gnd_net_),
            .in3(N__14564),
            .lcout(),
            .ltout(\this_vga_signals.M_hcounter_d6lt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIBPF11_9_LC_9_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIBPF11_9_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIBPF11_9_LC_9_20_1 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIBPF11_9_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__14408),
            .in2(N__8087),
            .in3(N__14271),
            .lcout(\this_vga_signals.M_hcounter_d6_0 ),
            .ltout(\this_vga_signals.M_hcounter_d6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUKG82_9_LC_9_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUKG82_9_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUKG82_9_LC_9_20_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIUKG82_9_LC_9_20_2  (
            .in0(N__8084),
            .in1(N__8060),
            .in2(N__8030),
            .in3(N__21384),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNIUKG82Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_1_sx_LC_9_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_1_sx_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_1_sx_LC_9_20_3 .LUT_INIT=16'b0000111101101111;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_1_sx_LC_9_20_3  (
            .in0(N__11092),
            .in1(N__8620),
            .in2(N__11467),
            .in3(N__8598),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_ac0_1_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_1_LC_9_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_1_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_1_LC_9_20_4 .LUT_INIT=16'b0000011100001101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_1_LC_9_20_4  (
            .in0(N__8599),
            .in1(N__11093),
            .in2(N__8003),
            .in3(N__8676),
            .lcout(\this_vga_signals.mult1_un75_sum_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_5_LC_9_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_5_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_5_LC_9_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_5_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11303),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21628),
            .ce(N__9069),
            .sr(N__11340));
    defparam \this_vga_signals.un4_haddress_if_m2_0_LC_9_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m2_0_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m2_0_LC_9_20_6 .LUT_INIT=16'b0100100000010010;
    LogicCell40 \this_vga_signals.un4_haddress_if_m2_0_LC_9_20_6  (
            .in0(N__10932),
            .in1(N__14717),
            .in2(N__11123),
            .in3(N__10163),
            .lcout(\this_vga_signals.if_m2_0 ),
            .ltout(\this_vga_signals.if_m2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_x0_LC_9_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_x0_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_x0_LC_9_20_7 .LUT_INIT=16'b0101011010101001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_x0_LC_9_20_7  (
            .in0(N__8630),
            .in1(N__8619),
            .in2(N__8000),
            .in3(N__8774),
            .lcout(\this_vga_signals.mult1_un75_sum_axb2_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_1_9_LC_9_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_1_9_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_1_9_LC_9_21_1 .LUT_INIT=16'b0010110011001010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_1_9_LC_9_21_1  (
            .in0(N__14565),
            .in1(N__14267),
            .in2(N__14449),
            .in3(N__14093),
            .lcout(\this_vga_signals.un1_haddress_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_3_LC_9_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_3_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_3_LC_9_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_3_LC_9_21_2  (
            .in0(N__8573),
            .in1(N__10983),
            .in2(N__11143),
            .in3(N__9792),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_axb2_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_N_4_i_1_LC_9_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_N_4_i_1_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_N_4_i_1_LC_9_21_3 .LUT_INIT=16'b0000111011000100;
    LogicCell40 \this_vga_signals.un4_haddress_N_4_i_1_LC_9_21_3  (
            .in0(N__9536),
            .in1(N__9722),
            .in2(N__8228),
            .in3(N__9509),
            .lcout(),
            .ltout(\this_vga_signals.N_4_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_N_4_i_LC_9_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_N_4_i_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_N_4_i_LC_9_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_N_4_i_LC_9_21_4  (
            .in0(N__14770),
            .in1(N__8225),
            .in2(N__8216),
            .in3(N__10208),
            .lcout(\this_vga_signals.N_4_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_i_3_LC_9_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_i_3_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_i_3_LC_9_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_i_3_LC_9_21_6  (
            .in0(N__8786),
            .in1(N__8507),
            .in2(_gnd_net_),
            .in3(N__9793),
            .lcout(\this_vga_signals.mult1_un68_sum_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_1_LC_9_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_1_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_1_LC_9_22_0 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_1_LC_9_22_0  (
            .in0(N__11470),
            .in1(N__10439),
            .in2(N__11550),
            .in3(N__10396),
            .lcout(\this_vga_signals.mult1_un82_sum_ac0_1 ),
            .ltout(\this_vga_signals.mult1_un82_sum_ac0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_9_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_9_22_1 .LUT_INIT=16'b0010001111011100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_LC_9_22_1  (
            .in0(N__10647),
            .in1(N__10580),
            .in2(N__8213),
            .in3(N__10670),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un82_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_axb_2_l_ofx_LC_9_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.un1_haddress_0_axb_2_l_ofx_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_axb_2_l_ofx_LC_9_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un1_haddress_0_axb_2_l_ofx_LC_9_22_2  (
            .in0(N__8210),
            .in1(N__10440),
            .in2(N__8204),
            .in3(N__10397),
            .lcout(\this_vga_signals.un1_haddress_0_axb_2_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_i_3_LC_9_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_i_3_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_i_3_LC_9_22_3 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_i_3_LC_9_22_3  (
            .in0(N__10398),
            .in1(_gnd_net_),
            .in2(N__10448),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.mult1_un75_sum_i_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_axb_3_l_fx_LC_9_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un1_haddress_0_axb_3_l_fx_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_axb_3_l_fx_LC_9_22_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un1_haddress_0_axb_3_l_fx_LC_9_22_4  (
            .in0(N__10446),
            .in1(N__9281),
            .in2(N__8320),
            .in3(N__10399),
            .lcout(\this_vga_signals.un1_haddress_0_axb_3_l_fxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGF3C6_9_LC_9_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGF3C6_9_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGF3C6_9_LC_9_22_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIGF3C6_9_LC_9_22_5  (
            .in0(N__8800),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8708),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNIGF3C6Z0Z_9 ),
            .ltout(\this_vga_signals.M_hcounter_q_esr_RNIGF3C6Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TA7_LC_9_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TA7_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TA7_LC_9_22_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TA7_LC_9_22_6  (
            .in0(N__8237),
            .in1(_gnd_net_),
            .in2(N__8375),
            .in3(N__8710),
            .lcout(\this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TAZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TA7_0_LC_9_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TA7_0_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TA7_0_LC_9_22_7 .LUT_INIT=16'b0001111111011111;
    LogicCell40 \this_vga_signals.un1_haddress_0_cry_5_c_RNIK1TA7_0_LC_9_22_7  (
            .in0(N__8709),
            .in1(N__8804),
            .in2(N__8452),
            .in3(N__8236),
            .lcout(\this_vga_signals.un1_haddress_0_cry_7_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_cry_1_c_LC_9_23_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_haddress_0_cry_1_c_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_cry_1_c_LC_9_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_haddress_0_cry_1_c_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__8970),
            .in2(N__8951),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\this_vga_signals.un1_haddress_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_cry_1_c_RNIDP44V02_LC_9_23_1 .C_ON=1'b1;
    defparam \this_vga_signals.un1_haddress_0_cry_1_c_RNIDP44V02_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_cry_1_c_RNIDP44V02_LC_9_23_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un1_haddress_0_cry_1_c_RNIDP44V02_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__8360),
            .in2(N__8354),
            .in3(N__8333),
            .lcout(\this_vga_signals.un1_haddress_0_cry_1_c_RNIDP44VZ0Z02 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_haddress_0_cry_1 ),
            .carryout(\this_vga_signals.un1_haddress_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_cry_2_c_RNIVPNA9D_LC_9_23_2 .C_ON=1'b1;
    defparam \this_vga_signals.un1_haddress_0_cry_2_c_RNIVPNA9D_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_cry_2_c_RNIVPNA9D_LC_9_23_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un1_haddress_0_cry_2_c_RNIVPNA9D_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__8330),
            .in2(N__8324),
            .in3(N__8291),
            .lcout(\this_vga_signals.un1_haddress_0_cry_2_c_RNIVPNA9DZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_haddress_0_cry_2 ),
            .carryout(\this_vga_signals.un1_haddress_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_cry_3_c_RNIBO4T72_LC_9_23_3 .C_ON=1'b1;
    defparam \this_vga_signals.un1_haddress_0_cry_3_c_RNIBO4T72_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_cry_3_c_RNIBO4T72_LC_9_23_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un1_haddress_0_cry_3_c_RNIBO4T72_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__8686),
            .in2(N__8288),
            .in3(N__8264),
            .lcout(\this_vga_signals.un1_haddress_0_cry_3_c_RNIBO4TZ0Z72 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_haddress_0_cry_3 ),
            .carryout(\this_vga_signals.un1_haddress_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_cry_4_c_RNI5SHJL_LC_9_23_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_haddress_0_cry_4_c_RNI5SHJL_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_cry_4_c_RNI5SHJL_LC_9_23_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un1_haddress_0_cry_4_c_RNI5SHJL_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__10222),
            .in2(N__8690),
            .in3(N__8249),
            .lcout(\this_vga_signals.un1_haddress_0_cry_4_c_RNI5SHJLZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_haddress_0_cry_4 ),
            .carryout(\this_vga_signals.un1_haddress_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_cry_5_THRU_LUT4_0_LC_9_23_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_haddress_0_cry_5_THRU_LUT4_0_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_cry_5_THRU_LUT4_0_LC_9_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.un1_haddress_0_cry_5_THRU_LUT4_0_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(N__8711),
            .in2(N__8246),
            .in3(N__8456),
            .lcout(\this_vga_signals.un1_haddress_0_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\this_vga_signals.un1_haddress_0_cry_5 ),
            .carryout(\this_vga_signals.un1_haddress_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_cry_6_c_RNI5KQU_LC_9_23_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_haddress_0_cry_6_c_RNI5KQU_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_cry_6_c_RNI5KQU_LC_9_23_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un1_haddress_0_cry_6_c_RNI5KQU_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(N__8453),
            .in2(_gnd_net_),
            .in3(N__8423),
            .lcout(\this_vga_signals.un1_haddress_0_cry_6_c_RNI5KQUZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_haddress_0_cry_6 ),
            .carryout(\this_vga_signals.un1_haddress_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_cry_7_c_RNIRVBS7_LC_9_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.un1_haddress_0_cry_7_c_RNIRVBS7_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_cry_7_c_RNIRVBS7_LC_9_23_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un1_haddress_0_cry_7_c_RNIRVBS7_LC_9_23_7  (
            .in0(N__14292),
            .in1(N__14116),
            .in2(N__8419),
            .in3(N__8402),
            .lcout(\this_vga_signals.un1_haddress_0_cry_7_c_RNIRVBSZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI0EQT_6_LC_10_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI0EQT_6_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI0EQT_6_LC_10_16_1 .LUT_INIT=16'b1111010011111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNI0EQT_6_LC_10_16_1  (
            .in0(N__9245),
            .in1(N__8882),
            .in2(N__9424),
            .in3(N__9224),
            .lcout(\this_vga_signals.m8_0_1_tz ),
            .ltout(\this_vga_signals.m8_0_1_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGQG41_8_LC_10_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGQG41_8_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGQG41_8_LC_10_16_2 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIGQG41_8_LC_10_16_2  (
            .in0(N__14177),
            .in1(_gnd_net_),
            .in2(N__8384),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\this_vga_signals.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_LC_10_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_LC_10_16_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \this_vga_signals.un4_haddress_g1_LC_10_16_3  (
            .in0(N__14790),
            .in1(N__9011),
            .in2(N__8381),
            .in3(N__9398),
            .lcout(),
            .ltout(\this_vga_signals.g1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_0_LC_10_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_0_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_0_LC_10_16_4 .LUT_INIT=16'b1110110010000000;
    LogicCell40 \this_vga_signals.un4_haddress_g1_0_LC_10_16_4  (
            .in0(N__10975),
            .in1(N__10052),
            .in2(N__8378),
            .in3(N__10199),
            .lcout(\this_vga_signals.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_7_LC_10_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_7_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_7_LC_10_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_7_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11242),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21596),
            .ce(N__9076),
            .sr(N__11334));
    defparam \this_vga_signals.M_hcounter_q_esr_8_LC_10_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_8_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_8_LC_10_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_8_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11219),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21596),
            .ce(N__9076),
            .sr(N__11334));
    defparam \this_vga_signals.M_hcounter_q_9_rep1_esr_LC_10_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_9_rep1_esr_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_9_rep1_esr_LC_10_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_9_rep1_esr_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11179),
            .lcout(\this_vga_signals.M_hcounter_q_9_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21596),
            .ce(N__9076),
            .sr(N__11334));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIN6RR_7_LC_10_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIN6RR_7_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIN6RR_7_LC_10_17_6 .LUT_INIT=16'b1111110011111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNIN6RR_7_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__9133),
            .in2(N__9231),
            .in3(N__9179),
            .lcout(\this_vga_signals.M_hcounter_q_fast_esr_RNIN6RRZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_7_LC_10_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_7_LC_10_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_7_LC_10_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_7_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11243),
            .lcout(\this_vga_signals.M_hcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21596),
            .ce(N__9076),
            .sr(N__11334));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIPO3M_7_LC_10_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIPO3M_7_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIPO3M_7_LC_10_18_1 .LUT_INIT=16'b0101111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNIPO3M_7_LC_10_18_1  (
            .in0(N__9358),
            .in1(_gnd_net_),
            .in2(N__9232),
            .in3(N__9135),
            .lcout(\this_vga_signals.N_75 ),
            .ltout(\this_vga_signals.N_75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_x1_1_LC_10_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_x1_1_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_x1_1_LC_10_18_2 .LUT_INIT=16'b0011100111001001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_x1_1_LC_10_18_2  (
            .in0(N__14530),
            .in1(N__8885),
            .in2(N__8483),
            .in3(N__8480),
            .lcout(\this_vga_signals.mult1_un54_sum_m_x1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_1_1_LC_10_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_1_1_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_1_1_LC_10_18_3 .LUT_INIT=16'b0000010000101011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_1_1_LC_10_18_3  (
            .in0(N__9357),
            .in1(N__9134),
            .in2(N__8913),
            .in3(N__9180),
            .lcout(\this_vga_signals.mult1_un54_sum_m_1_1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_m_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_x0_1_LC_10_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_x0_1_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_x0_1_LC_10_18_4 .LUT_INIT=16'b0011110001100110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_x0_1_LC_10_18_4  (
            .in0(N__14531),
            .in1(N__8886),
            .in2(N__8474),
            .in3(N__8471),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_m_x0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_ns_1_LC_10_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_ns_1_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_ns_1_LC_10_18_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_m_ns_1_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__8924),
            .in2(N__8465),
            .in3(N__8462),
            .lcout(\this_vga_signals.mult1_un54_sum_m_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_6_LC_10_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_6_LC_10_18_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_6_LC_10_18_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_6_LC_10_18_6  (
            .in0(N__11272),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21605),
            .ce(N__9054),
            .sr(N__11337));
    defparam \this_vga_signals.M_hcounter_q_6_rep1_esr_LC_10_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_6_rep1_esr_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_rep1_esr_LC_10_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_rep1_esr_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11271),
            .lcout(\this_vga_signals.M_hcounter_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21605),
            .ce(N__9054),
            .sr(N__11337));
    defparam \this_vga_signals.M_hcounter_q_7_rep1_esr_RNIJOM71_LC_10_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_7_rep1_esr_RNIJOM71_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_7_rep1_esr_RNIJOM71_LC_10_19_0 .LUT_INIT=16'b0111100100001001;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_rep1_esr_RNIJOM71_LC_10_19_0  (
            .in0(N__9145),
            .in1(N__8914),
            .in2(N__9188),
            .in3(N__8887),
            .lcout(),
            .ltout(\this_vga_signals.M_hcounter_q_7_rep1_esr_RNIJOMZ0Z71_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_8_rep1_esr_RNI1Q1C1_LC_10_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_8_rep1_esr_RNI1Q1C1_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_8_rep1_esr_RNI1Q1C1_LC_10_19_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_rep1_esr_RNI1Q1C1_LC_10_19_1  (
            .in0(N__20360),
            .in1(_gnd_net_),
            .in2(N__8522),
            .in3(N__9369),
            .lcout(\this_vga_signals.m8_0_2 ),
            .ltout(\this_vga_signals.m8_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_1_LC_10_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_1_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_1_LC_10_19_2 .LUT_INIT=16'b0010100010001000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_1_LC_10_19_2  (
            .in0(N__10963),
            .in1(N__8888),
            .in2(N__8519),
            .in3(N__9335),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_10_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_10_19_3 .LUT_INIT=16'b1111111011101100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_10_19_3  (
            .in0(N__10027),
            .in1(N__10086),
            .in2(N__8516),
            .in3(N__10164),
            .lcout(\this_vga_signals.mult1_un61_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_8_rep1_esr_RNIKFGM4_LC_10_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_8_rep1_esr_RNIKFGM4_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_8_rep1_esr_RNIKFGM4_LC_10_19_4 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_rep1_esr_RNIKFGM4_LC_10_19_4  (
            .in0(N__9370),
            .in1(N__9393),
            .in2(N__8942),
            .in3(N__9005),
            .lcout(\this_vga_signals.mult1_un54_sum_i_0_3 ),
            .ltout(\this_vga_signals.mult1_un54_sum_i_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_31_LC_10_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_31_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_31_LC_10_19_5 .LUT_INIT=16'b1010111111110101;
    LogicCell40 \this_vga_signals.un4_haddress_g0_31_LC_10_19_5  (
            .in0(N__14740),
            .in1(_gnd_net_),
            .in2(N__8513),
            .in3(N__10964),
            .lcout(\this_vga_signals.g1_6_0 ),
            .ltout(\this_vga_signals.g1_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_13_N_2L1_LC_10_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_13_N_2L1_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_13_N_2L1_LC_10_19_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un4_haddress_g0_13_N_2L1_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8510),
            .in3(N__10028),
            .lcout(),
            .ltout(\this_vga_signals.g0_13_N_2L1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_13_N_4L5_LC_10_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_13_N_4L5_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_13_N_4L5_LC_10_19_7 .LUT_INIT=16'b0010000100010010;
    LogicCell40 \this_vga_signals.un4_haddress_g0_13_N_4L5_LC_10_19_7  (
            .in0(N__8503),
            .in1(N__8492),
            .in2(N__8486),
            .in3(N__9779),
            .lcout(\this_vga_signals.g0_13_N_4L5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_10_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_10_20_0 .LUT_INIT=16'b1111011000001001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_10_20_0  (
            .in0(N__8663),
            .in1(N__8621),
            .in2(N__8600),
            .in3(N__8776),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_x1_LC_10_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_x1_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_x1_LC_10_20_1 .LUT_INIT=16'b0101011010010101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_x1_LC_10_20_1  (
            .in0(N__11088),
            .in1(N__8777),
            .in2(N__10992),
            .in3(N__8664),
            .lcout(\this_vga_signals.mult1_un75_sum_ac0_3_0_1_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_0_0_LC_10_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_0_0_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_0_0_LC_10_20_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_0_0_LC_10_20_2  (
            .in0(N__10924),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11087),
            .lcout(\this_vga_signals.mult1_un75_sum_axb2_0_0 ),
            .ltout(\this_vga_signals.mult1_un75_sum_axb2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_x1_LC_10_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_x1_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_x1_LC_10_20_3 .LUT_INIT=16'b1001011010100101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_x1_LC_10_20_3  (
            .in0(N__8775),
            .in1(N__8593),
            .in2(N__8624),
            .in3(N__8618),
            .lcout(\this_vga_signals.mult1_un75_sum_axb2_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI43A65_5_LC_10_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI43A65_5_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI43A65_5_LC_10_20_4 .LUT_INIT=16'b0110100110100101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI43A65_5_LC_10_20_4  (
            .in0(N__14752),
            .in1(N__9006),
            .in2(N__10972),
            .in3(N__9334),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5 ),
            .ltout(\this_vga_signals.M_hcounter_q_esr_RNI43A65Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_3_LC_10_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_3_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_3_LC_10_20_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_3_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(N__8594),
            .in2(N__8576),
            .in3(N__8662),
            .lcout(\this_vga_signals.mult1_un68_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_10_3_0_a2_0_0_LC_10_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_10_3_0_a2_0_0_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_10_3_0_a2_0_0_LC_10_20_6 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \this_vga_signals.un4_haddress_g0_10_3_0_a2_0_0_LC_10_20_6  (
            .in0(N__14753),
            .in1(N__10201),
            .in2(N__10973),
            .in3(N__10060),
            .lcout(\this_vga_signals.g0_10_3_0_a2_0_0 ),
            .ltout(\this_vga_signals.g0_10_3_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_1_3_a2_LC_10_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_1_3_a2_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_1_3_a2_LC_10_20_7 .LUT_INIT=16'b1110000100011110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_1_3_a2_LC_10_20_7  (
            .in0(N__8567),
            .in1(N__8555),
            .in2(N__8540),
            .in3(N__9780),
            .lcout(\this_vga_signals.mult1_un68_sum_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_10_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_10_21_0 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_10_21_0  (
            .in0(N__11131),
            .in1(_gnd_net_),
            .in2(N__9796),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.mult1_un75_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_ns_LC_10_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_ns_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_ns_LC_10_21_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb2_ns_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__8537),
            .in2(N__8531),
            .in3(N__8678),
            .lcout(\this_vga_signals.mult1_un75_sum_axb2_i ),
            .ltout(\this_vga_signals.mult1_un75_sum_axb2_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc2_LC_10_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc2_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc2_LC_10_21_3 .LUT_INIT=16'b1111000000101101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc2_LC_10_21_3  (
            .in0(N__9271),
            .in1(N__11132),
            .in2(N__8789),
            .in3(N__8734),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_x0_LC_10_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_x0_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_x0_LC_10_21_4 .LUT_INIT=16'b0100101100101101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_x0_LC_10_21_4  (
            .in0(N__10982),
            .in1(N__8785),
            .in2(N__11144),
            .in3(N__8679),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_ac0_3_0_1_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_ns_LC_10_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_ns_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_ns_LC_10_21_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_1_ns_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(N__8744),
            .in2(N__8738),
            .in3(N__9781),
            .lcout(\this_vga_signals.mult1_un75_sum_ac0_3_0_1 ),
            .ltout(\this_vga_signals.mult1_un75_sum_ac0_3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_LC_10_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_LC_10_21_6 .LUT_INIT=16'b0000001111101011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_ac0_3_0_LC_10_21_6  (
            .in0(N__8735),
            .in1(N__9272),
            .in2(N__8726),
            .in3(N__8723),
            .lcout(\this_vga_signals.mult1_un75_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_10_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_10_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__10445),
            .in2(N__10411),
            .in3(N__8717),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_0_9_LC_10_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_0_9_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_0_9_LC_10_22_1 .LUT_INIT=16'b0110101100101000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_0_9_LC_10_22_1  (
            .in0(N__14266),
            .in1(N__14077),
            .in2(N__14472),
            .in3(N__14578),
            .lcout(\this_vga_signals.N_510_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axb2_LC_10_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axb2_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axb2_LC_10_22_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axb2_LC_10_22_2  (
            .in0(N__8851),
            .in1(N__11469),
            .in2(N__10410),
            .in3(N__10444),
            .lcout(\this_vga_signals.mult1_un82_sum_axb2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_1_0_LC_10_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_1_0_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_1_0_LC_10_22_3 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_1_0_LC_10_22_3  (
            .in0(N__11148),
            .in1(N__10980),
            .in2(_gnd_net_),
            .in3(N__8680),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_10_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_10_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_10_22_4  (
            .in0(N__14801),
            .in1(N__9277),
            .in2(N__8633),
            .in3(N__10202),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_1_i ),
            .ltout(\this_vga_signals.mult1_un75_sum_axbxc3_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_0_0_LC_10_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_0_0_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_0_0_LC_10_22_5 .LUT_INIT=16'b0100011001100100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_0_0_LC_10_22_5  (
            .in0(N__11468),
            .in1(N__8852),
            .in2(N__8843),
            .in3(N__10400),
            .lcout(\this_vga_signals.mult1_un82_sum_ac0_3_0_0 ),
            .ltout(\this_vga_signals.mult1_un82_sum_ac0_3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_i_3_LC_10_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_i_3_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_i_3_LC_10_22_6 .LUT_INIT=16'b1100011011000011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_i_3_LC_10_22_6  (
            .in0(N__10651),
            .in1(N__10671),
            .in2(N__8840),
            .in3(N__10611),
            .lcout(\this_vga_signals.un1_haddress_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI5HOBQC_1_LC_10_22_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI5HOBQC_1_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI5HOBQC_1_LC_10_22_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI5HOBQC_1_LC_10_22_7  (
            .in0(N__10672),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11541),
            .lcout(\this_vga_signals.M_hcounter_q_RNI5HOBQCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIPIQRNR_2_LC_10_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIPIQRNR_2_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIPIQRNR_2_LC_10_23_0 .LUT_INIT=16'b0011111110010110;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIPIQRNR_2_LC_10_23_0  (
            .in0(N__11476),
            .in1(N__10649),
            .in2(N__10586),
            .in3(N__10612),
            .lcout(\this_vga_signals.M_hcounter_q_RNIPIQRNRZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.new_pixel_1_axb_1_N_4L5_x1_LC_10_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.new_pixel_1_axb_1_N_4L5_x1_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.new_pixel_1_axb_1_N_4L5_x1_LC_10_23_1 .LUT_INIT=16'b0111011110011001;
    LogicCell40 \this_vga_signals.new_pixel_1_axb_1_N_4L5_x1_LC_10_23_1  (
            .in0(N__10650),
            .in1(N__10584),
            .in2(_gnd_net_),
            .in3(N__10610),
            .lcout(),
            .ltout(\this_vga_signals.new_pixel_1_axb_1_N_4L5_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI8TTVN32_2_LC_10_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI8TTVN32_2_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI8TTVN32_2_LC_10_23_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI8TTVN32_2_LC_10_23_2  (
            .in0(N__9466),
            .in1(_gnd_net_),
            .in2(N__8837),
            .in3(N__8834),
            .lcout(),
            .ltout(\this_vga_signals.M_hcounter_q_RNI8TTVN32Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIU31PMD_1_LC_10_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIU31PMD_1_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIU31PMD_1_LC_10_23_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIU31PMD_1_LC_10_23_3  (
            .in0(N__8828),
            .in1(N__8971),
            .in2(N__8822),
            .in3(N__9582),
            .lcout(\this_vga_signals.new_pixel_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_9_LC_10_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_9_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_9_LC_10_23_4 .LUT_INIT=16'b1001010011010111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_9_LC_10_23_4  (
            .in0(N__14265),
            .in1(N__14076),
            .in2(N__14471),
            .in3(N__14577),
            .lcout(),
            .ltout(\this_vga_signals.N_510_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIIV9H5_9_LC_10_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIIV9H5_9_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIIV9H5_9_LC_10_23_5 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIIV9H5_9_LC_10_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8807),
            .in3(N__10221),
            .lcout(\this_vga_signals.un1_haddress_0_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_4_LC_10_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_4_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_4_LC_10_23_6 .LUT_INIT=16'b1010101101010100;
    LogicCell40 \this_vga_signals.un4_haddress_g0_4_LC_10_23_6  (
            .in0(N__10609),
            .in1(N__11475),
            .in2(N__9467),
            .in3(N__10648),
            .lcout(\this_vga_signals.mult1_un89_sum_axbxc3_0 ),
            .ltout(\this_vga_signals.mult1_un89_sum_axbxc3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_haddress_0_cry_1_c_RNO_LC_10_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.un1_haddress_0_cry_1_c_RNO_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_haddress_0_cry_1_c_RNO_LC_10_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un1_haddress_0_cry_1_c_RNO_LC_10_23_7  (
            .in0(N__8972),
            .in1(N__9581),
            .in2(N__8954),
            .in3(N__9549),
            .lcout(\this_vga_signals.un1_haddress_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGQG41_0_8_LC_11_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGQG41_0_8_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGQG41_0_8_LC_11_16_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIGQG41_0_8_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__8938),
            .in2(_gnd_net_),
            .in3(N__14178),
            .lcout(\this_vga_signals.g1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI58601_7_LC_11_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI58601_7_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI58601_7_LC_11_17_0 .LUT_INIT=16'b0010101100100000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNI58601_7_LC_11_17_0  (
            .in0(N__9367),
            .in1(N__9142),
            .in2(N__9233),
            .in3(N__9185),
            .lcout(\this_vga_signals.ANC2_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_8_rep1_esr_LC_11_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_8_rep1_esr_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_rep1_esr_LC_11_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_rep1_esr_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11218),
            .lcout(\this_vga_signals.M_hcounter_q_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21590),
            .ce(N__9077),
            .sr(N__11333));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_2_LC_11_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_2_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_2_LC_11_17_2 .LUT_INIT=16'b0110101111010111;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_2_LC_11_17_2  (
            .in0(N__9368),
            .in1(N__9143),
            .in2(N__8915),
            .in3(N__9186),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_LC_11_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_LC_11_17_3 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_LC_11_17_3  (
            .in0(N__8884),
            .in1(_gnd_net_),
            .in2(N__8918),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_7_rep1_esr_LC_11_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_7_rep1_esr_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_rep1_esr_LC_11_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_rep1_esr_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11241),
            .lcout(\this_vga_signals.M_hcounter_q_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21590),
            .ce(N__9077),
            .sr(N__11333));
    defparam \this_vga_signals.M_hcounter_q_5_rep1_esr_LC_11_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_5_rep1_esr_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_rep1_esr_LC_11_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_rep1_esr_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11302),
            .lcout(\this_vga_signals.M_hcounter_q_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21590),
            .ce(N__9077),
            .sr(N__11333));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI52HL_9_LC_11_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI52HL_9_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI52HL_9_LC_11_17_6 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNI52HL_9_LC_11_17_6  (
            .in0(N__9244),
            .in1(N__8883),
            .in2(_gnd_net_),
            .in3(N__9222),
            .lcout(\this_vga_signals.M_hcounter_q_fast_esr_RNI52HLZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_9_LC_11_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_9_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_9_LC_11_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_9_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11178),
            .lcout(\this_vga_signals.M_hcounter_q_fastZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21590),
            .ce(N__9077),
            .sr(N__11333));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIHH441_5_LC_11_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIHH441_5_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIHH441_5_LC_11_18_0 .LUT_INIT=16'b1111101101001011;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNIHH441_5_LC_11_18_0  (
            .in0(N__9223),
            .in1(N__9181),
            .in2(N__9146),
            .in3(N__9089),
            .lcout(),
            .ltout(\this_vga_signals.M_hcounter_q_fast_esr_RNIHH441Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI56982_8_LC_11_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI56982_8_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI56982_8_LC_11_18_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNI56982_8_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__9083),
            .in2(N__9098),
            .in3(N__9095),
            .lcout(\this_vga_signals.m8_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_5_LC_11_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_5_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_5_LC_11_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_5_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11301),
            .lcout(\this_vga_signals.M_hcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21597),
            .ce(N__9058),
            .sr(N__11335));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_8_LC_11_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_8_LC_11_18_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_8_LC_11_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_8_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11217),
            .lcout(\this_vga_signals.M_hcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21597),
            .ce(N__9058),
            .sr(N__11335));
    defparam \this_vga_signals.un4_haddress_g0_17_LC_11_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_17_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_17_LC_11_19_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_vga_signals.un4_haddress_g0_17_LC_11_19_0  (
            .in0(N__9392),
            .in1(N__9010),
            .in2(N__14813),
            .in3(N__8984),
            .lcout(\this_vga_signals.g1_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g4_1_1_LC_11_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g4_1_1_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g4_1_1_LC_11_19_1 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \this_vga_signals.un4_haddress_g4_1_1_LC_11_19_1  (
            .in0(N__10049),
            .in1(N__10171),
            .in2(_gnd_net_),
            .in3(N__10251),
            .lcout(),
            .ltout(\this_vga_signals.g4_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g4_1_LC_11_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g4_1_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g4_1_LC_11_19_2 .LUT_INIT=16'b1110000000011111;
    LogicCell40 \this_vga_signals.un4_haddress_g4_1_LC_11_19_2  (
            .in0(N__14798),
            .in1(N__9323),
            .in2(N__8975),
            .in3(N__10907),
            .lcout(\this_vga_signals.g4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_8_LC_11_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_8_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_8_LC_11_19_3 .LUT_INIT=16'b0110101111010111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_8_LC_11_19_3  (
            .in0(N__14263),
            .in1(N__14038),
            .in2(N__14479),
            .in3(N__14534),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_0_a2_0_0_LC_11_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_0_a2_0_0_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_0_a2_0_0_LC_11_19_4 .LUT_INIT=16'b1001101001011001;
    LogicCell40 \this_vga_signals.un4_haddress_g1_0_a2_0_0_LC_11_19_4  (
            .in0(N__10050),
            .in1(N__10908),
            .in2(N__10200),
            .in3(N__14799),
            .lcout(\this_vga_signals.g1_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIJLEA3_6_LC_11_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIJLEA3_6_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIJLEA3_6_LC_11_19_6 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNIJLEA3_6_LC_11_19_6  (
            .in0(N__9428),
            .in1(N__9407),
            .in2(N__9397),
            .in3(N__9371),
            .lcout(\this_vga_signals.m8_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_16_LC_11_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_16_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_16_LC_11_19_7 .LUT_INIT=16'b0110101111010111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_16_LC_11_19_7  (
            .in0(N__14264),
            .in1(N__14039),
            .in2(N__14480),
            .in3(N__14535),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_14_LC_11_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_14_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_14_LC_11_20_0 .LUT_INIT=16'b1110101010000000;
    LogicCell40 \this_vga_signals.un4_haddress_g0_14_LC_11_20_0  (
            .in0(N__10170),
            .in1(N__10909),
            .in2(N__9317),
            .in3(N__10055),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_21_LC_11_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_21_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_21_LC_11_20_1 .LUT_INIT=16'b0000000100110111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_21_LC_11_20_1  (
            .in0(N__9308),
            .in1(N__11116),
            .in2(N__9296),
            .in3(N__10945),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_0_a2_0_LC_11_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_0_a2_0_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_0_a2_0_LC_11_20_2 .LUT_INIT=16'b0010010011011011;
    LogicCell40 \this_vga_signals.un4_haddress_g1_0_a2_0_LC_11_20_2  (
            .in0(N__10168),
            .in1(N__14754),
            .in2(N__10979),
            .in3(N__10054),
            .lcout(\this_vga_signals.N_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_29_LC_11_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_29_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_29_LC_11_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_29_LC_11_20_3  (
            .in0(N__10056),
            .in1(N__9293),
            .in2(N__10793),
            .in3(N__9791),
            .lcout(\this_vga_signals.mult1_un75_sum_axb2_i_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g4_LC_11_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g4_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g4_LC_11_20_4 .LUT_INIT=16'b0000000011010010;
    LogicCell40 \this_vga_signals.un4_haddress_g4_LC_11_20_4  (
            .in0(N__9287),
            .in1(N__9273),
            .in2(N__11142),
            .in3(N__9507),
            .lcout(\this_vga_signals.g4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_9_LC_11_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_9_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_9_LC_11_20_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.un4_haddress_g0_9_LC_11_20_5  (
            .in0(N__11418),
            .in1(N__11117),
            .in2(_gnd_net_),
            .in3(N__9790),
            .lcout(\this_vga_signals.mult1_un75_sum_ac0_1_1 ),
            .ltout(\this_vga_signals.mult1_un75_sum_ac0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_13_LC_11_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_13_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_13_LC_11_20_6 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_13_LC_11_20_6  (
            .in0(N__11118),
            .in1(N__9524),
            .in2(N__9518),
            .in3(N__9506),
            .lcout(\this_vga_signals.g1_1_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_1_LC_11_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_1_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_1_LC_11_20_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \this_vga_signals.un4_haddress_g1_1_LC_11_20_7  (
            .in0(N__10053),
            .in1(N__10250),
            .in2(_gnd_net_),
            .in3(N__10169),
            .lcout(\this_vga_signals.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_0_2_LC_11_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_0_2_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_0_2_LC_11_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_0_2_LC_11_21_0  (
            .in0(N__9515),
            .in1(N__10215),
            .in2(N__14814),
            .in3(N__9508),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_12_LC_11_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_12_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_12_LC_11_21_1 .LUT_INIT=16'b0010110101111000;
    LogicCell40 \this_vga_signals.un4_haddress_g0_12_LC_11_21_1  (
            .in0(N__9488),
            .in1(N__9482),
            .in2(N__9476),
            .in3(N__9473),
            .lcout(\this_vga_signals.N_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_7_LC_11_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_7_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_7_LC_11_21_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.un4_haddress_g0_7_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(N__9452),
            .in2(_gnd_net_),
            .in3(N__14800),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0 ),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_2_0_a2_LC_11_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_2_0_a2_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_2_0_a2_LC_11_21_3 .LUT_INIT=16'b1010100101010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_2_0_a2_LC_11_21_3  (
            .in0(N__9730),
            .in1(N__9655),
            .in2(N__9443),
            .in3(N__9786),
            .lcout(\this_vga_signals.mult1_un68_sum_0_3 ),
            .ltout(\this_vga_signals.mult1_un68_sum_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g1_0_a2_LC_11_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g1_0_a2_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g1_0_a2_LC_11_21_4 .LUT_INIT=16'b1011101001000101;
    LogicCell40 \this_vga_signals.un4_haddress_g1_0_a2_LC_11_21_4  (
            .in0(N__9707),
            .in1(N__11110),
            .in2(N__9440),
            .in3(N__9437),
            .lcout(\this_vga_signals.g1_0_a2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_11_LC_11_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_11_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_11_LC_11_21_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.un4_haddress_g0_11_LC_11_21_5  (
            .in0(N__11471),
            .in1(N__11085),
            .in2(_gnd_net_),
            .in3(N__9785),
            .lcout(\this_vga_signals.mult1_un75_sum_ac0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_12_0_a2_LC_11_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_12_0_a2_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_12_0_a2_LC_11_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_12_0_a2_LC_11_21_6  (
            .in0(N__11086),
            .in1(N__10981),
            .in2(N__9797),
            .in3(N__9731),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_axb2_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_1_LC_11_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_1_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_1_LC_11_21_7 .LUT_INIT=16'b0001111100011001;
    LogicCell40 \this_vga_signals.un4_haddress_g0_1_LC_11_21_7  (
            .in0(N__9721),
            .in1(N__9633),
            .in2(N__9710),
            .in3(N__9706),
            .lcout(\this_vga_signals.mult1_un75_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_x2_0_0_a2_3_LC_11_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_x2_0_0_a2_3_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_x2_0_0_a2_3_LC_11_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_x2_0_0_a2_3_LC_11_22_0  (
            .in0(N__9644),
            .in1(N__10220),
            .in2(N__9677),
            .in3(N__9635),
            .lcout(),
            .ltout(\this_vga_signals.g0_i_x2_0_0_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_LC_11_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_LC_11_22_1 .LUT_INIT=16'b0110000000000110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_LC_11_22_1  (
            .in0(N__11549),
            .in1(N__9854),
            .in2(N__9698),
            .in3(N__9694),
            .lcout(),
            .ltout(\this_vga_signals.if_i4_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_LC_11_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_LC_11_22_2 .LUT_INIT=16'b0000011011110110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_LC_11_22_2  (
            .in0(N__9695),
            .in1(N__9620),
            .in2(N__9686),
            .in3(N__9683),
            .lcout(\this_vga_signals.mult1_un89_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_i_x2_0_0_a2_0_LC_11_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_i_x2_0_0_a2_0_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_i_x2_0_0_a2_0_LC_11_22_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un4_haddress_g0_i_x2_0_0_a2_0_LC_11_22_4  (
            .in0(N__11445),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14802),
            .lcout(\this_vga_signals.g0_i_x2_0_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_10_LC_11_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_10_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_10_LC_11_22_5 .LUT_INIT=16'b0001000100010111;
    LogicCell40 \this_vga_signals.un4_haddress_g0_10_LC_11_22_5  (
            .in0(N__11149),
            .in1(N__10923),
            .in2(N__9668),
            .in3(N__9659),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_0 ),
            .ltout(\this_vga_signals.mult1_un75_sum_axbxc3_1_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_0_a2_4_LC_11_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_0_a2_4_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_0_a2_4_LC_11_22_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_0_a2_4_LC_11_22_6  (
            .in0(N__11378),
            .in1(N__10219),
            .in2(N__9638),
            .in3(N__9634),
            .lcout(\this_vga_signals.g0_0_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_address_buffer_q_esr_0_LC_11_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_0_LC_11_23_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_0_LC_11_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_0_LC_11_23_1  (
            .in0(N__9607),
            .in1(N__9588),
            .in2(_gnd_net_),
            .in3(N__9563),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21629),
            .ce(N__15292),
            .sr(N__15204));
    defparam \this_vga_signals.M_address_buffer_q_esr_1_LC_11_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_1_LC_11_23_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_1_LC_11_23_2 .LUT_INIT=16'b1010101001100101;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_1_LC_11_23_2  (
            .in0(N__10673),
            .in1(N__10652),
            .in2(N__10622),
            .in3(N__10585),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21629),
            .ce(N__15292),
            .sr(N__15204));
    defparam \this_vga_signals.M_address_buffer_q_esr_2_LC_11_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_2_LC_11_23_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_2_LC_11_23_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_2_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(N__10447),
            .in2(_gnd_net_),
            .in3(N__10412),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21629),
            .ce(N__15292),
            .sr(N__15204));
    defparam \this_vga_signals.M_address_buffer_q_esr_4_LC_11_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_4_LC_11_24_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_4_LC_11_24_0 .LUT_INIT=16'b1111111011111000;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_4_LC_11_24_0  (
            .in0(N__10259),
            .in1(N__10223),
            .in2(N__10094),
            .in3(N__10061),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21633),
            .ce(N__15306),
            .sr(N__15197));
    defparam \this_vga_signals.M_address_buffer_q_esr_12_LC_12_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_12_LC_12_19_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_12_LC_12_19_1 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_12_LC_12_19_1  (
            .in0(N__11789),
            .in1(N__11822),
            .in2(N__11807),
            .in3(N__11774),
            .lcout(M_this_vga_signals_address_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21598),
            .ce(N__15268),
            .sr(N__15179));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_20_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__9860),
            .in2(N__11554),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_12_20_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_12_20_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_12_20_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_12_20_1  (
            .in0(N__12921),
            .in1(N__11441),
            .in2(_gnd_net_),
            .in3(N__9806),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__21606),
            .ce(),
            .sr(N__11338));
    defparam \this_vga_signals.M_hcounter_q_3_LC_12_20_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_12_20_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_12_20_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_12_20_2  (
            .in0(N__12896),
            .in1(N__11122),
            .in2(_gnd_net_),
            .in3(N__9803),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__21606),
            .ce(),
            .sr(N__11338));
    defparam \this_vga_signals.M_hcounter_q_4_LC_12_20_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_12_20_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_12_20_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_12_20_3  (
            .in0(N__12922),
            .in1(N__10910),
            .in2(_gnd_net_),
            .in3(N__9800),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__21606),
            .ce(),
            .sr(N__11338));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRD_LC_12_20_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRD_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRD_LC_12_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRD_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(N__14758),
            .in2(_gnd_net_),
            .in3(N__11276),
            .lcout(\this_vga_signals.un1_M_hcounter_d_cry_4_c_RNICHRDZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSD_LC_12_20_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSD_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSD_LC_12_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSD_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(N__14602),
            .in2(_gnd_net_),
            .in3(N__11246),
            .lcout(\this_vga_signals.un1_M_hcounter_d_cry_5_c_RNIEKSDZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTD_LC_12_20_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTD_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTD_LC_12_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTD_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(N__14098),
            .in2(_gnd_net_),
            .in3(N__11222),
            .lcout(\this_vga_signals.un1_M_hcounter_d_cry_6_c_RNIGNTDZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUD_LC_12_20_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUD_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUD_LC_12_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUD_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(N__14279),
            .in2(_gnd_net_),
            .in3(N__11186),
            .lcout(\this_vga_signals.un1_M_hcounter_d_cry_7_c_RNIIQUDZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVD_LC_12_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVD_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVD_LC_12_21_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVD_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(N__14463),
            .in2(_gnd_net_),
            .in3(N__11183),
            .lcout(\this_vga_signals.un1_M_hcounter_d_cry_8_c_RNIKTVDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU45J5_9_LC_12_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU45J5_9_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU45J5_9_LC_12_21_1 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU45J5_9_LC_12_21_1  (
            .in0(N__11573),
            .in1(N__12884),
            .in2(_gnd_net_),
            .in3(N__11972),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNIU45J5Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIH06Q6_9_LC_12_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIH06Q6_9_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIH06Q6_9_LC_12_21_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIH06Q6_9_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(N__12885),
            .in2(_gnd_net_),
            .in3(N__15126),
            .lcout(\this_vga_signals.N_550_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_4_0_LC_12_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_4_0_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_4_0_LC_12_21_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un4_haddress_g0_4_0_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(N__11084),
            .in2(_gnd_net_),
            .in3(N__10906),
            .lcout(\this_vga_signals.g0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_0_9_LC_12_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_0_9_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIG53K_0_9_LC_12_21_7 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIG53K_0_9_LC_12_21_7  (
            .in0(N__14462),
            .in1(N__14278),
            .in2(_gnd_net_),
            .in3(N__14097),
            .lcout(debug_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_g0_0_a2_1_LC_12_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_g0_0_a2_1_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_g0_0_a2_1_LC_12_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un4_haddress_g0_0_a2_1_LC_12_22_5  (
            .in0(N__11548),
            .in1(N__11446),
            .in2(_gnd_net_),
            .in3(N__14791),
            .lcout(\this_vga_signals.g0_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_3_LC_12_22_6 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_3_LC_12_22_6 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_3_LC_12_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_3_LC_12_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11357),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21617),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_2_LC_12_22_7 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_2_LC_12_22_7 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_2_LC_12_22_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_delay_clk.M_pipe_q_2_LC_12_22_7  (
            .in0(N__11372),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21617),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_13_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_13_18_4 .LUT_INIT=16'b0001111000101101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_13_18_4  (
            .in0(N__13036),
            .in1(N__13453),
            .in2(N__13289),
            .in3(N__13222),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_0_0 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m7_0_o4_LC_13_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m7_0_o4_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m7_0_o4_LC_13_18_5 .LUT_INIT=16'b1000111011101000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m7_0_o4_LC_13_18_5  (
            .in0(N__13114),
            .in1(N__13199),
            .in2(N__11351),
            .in3(N__11837),
            .lcout(\this_vga_signals.if_N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_LC_13_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_LC_13_19_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_LC_13_19_0  (
            .in0(N__11896),
            .in1(N__11871),
            .in2(_gnd_net_),
            .in3(N__11931),
            .lcout(\this_vga_signals.mult1_un40_sum_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_4_LC_13_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_4_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_4_LC_13_19_1 .LUT_INIT=16'b0100100010000100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_4_LC_13_19_1  (
            .in0(N__11932),
            .in1(N__12809),
            .in2(N__11878),
            .in3(N__11897),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_13_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_13_19_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__11911),
            .in2(_gnd_net_),
            .in3(N__11918),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3 ),
            .ltout(\this_vga_signals.mult1_un47_sum_ac0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_LC_13_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_LC_13_19_3 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_LC_13_19_3  (
            .in0(N__11802),
            .in1(N__11821),
            .in2(N__11348),
            .in3(N__11772),
            .lcout(\this_vga_signals.mult1_un47_sum_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_2_LC_13_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_2_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_2_LC_13_19_5 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_2_LC_13_19_5  (
            .in0(N__11933),
            .in1(_gnd_net_),
            .in2(N__11879),
            .in3(N__12808),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_1_2 ),
            .ltout(\this_vga_signals.mult1_un47_sum_axbxc3_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_0_LC_13_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_0_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_0_LC_13_19_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_0_LC_13_19_6  (
            .in0(N__13021),
            .in1(_gnd_net_),
            .in2(N__11810),
            .in3(N__13452),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_axb1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_13_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_13_19_7 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_13_19_7  (
            .in0(N__11803),
            .in1(N__11788),
            .in2(N__11777),
            .in3(N__11773),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_13_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_13_20_7 .LUT_INIT=16'b0000000101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_13_20_7  (
            .in0(N__13025),
            .in1(N__13198),
            .in2(N__12718),
            .in3(N__13121),
            .lcout(\this_vga_signals.un2_vsynclt8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI6CLG4_5_LC_13_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI6CLG4_5_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI6CLG4_5_LC_13_21_3 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI6CLG4_5_LC_13_21_3  (
            .in0(N__13454),
            .in1(N__11945),
            .in2(N__11759),
            .in3(N__13739),
            .lcout(this_vga_signals_vsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_address_buffer_q_esr_6_LC_13_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_6_LC_13_22_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_6_LC_13_22_2 .LUT_INIT=16'b0001010110111000;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_6_LC_13_22_2  (
            .in0(N__14302),
            .in1(N__14117),
            .in2(N__14615),
            .in3(N__14478),
            .lcout(M_this_vga_signals_address_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21615),
            .ce(N__15299),
            .sr(N__15183));
    defparam \this_vga_signals.un5_vaddress_if_m7_0_m2_LC_14_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m7_0_m2_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m7_0_m2_LC_14_17_1 .LUT_INIT=16'b0110000011111001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m7_0_m2_LC_14_17_1  (
            .in0(N__13033),
            .in1(N__12490),
            .in2(N__13124),
            .in3(N__11621),
            .lcout(\this_vga_signals.if_N_10 ),
            .ltout(\this_vga_signals.if_N_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_14_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_14_17_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_14_17_2  (
            .in0(N__12330),
            .in1(N__12346),
            .in2(N__11615),
            .in3(N__12186),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_0_0 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_c2_LC_14_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_c2_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_c2_LC_14_17_3 .LUT_INIT=16'b1111010101010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_c2_LC_14_17_3  (
            .in0(N__13202),
            .in1(_gnd_net_),
            .in2(N__11612),
            .in3(N__12713),
            .lcout(\this_vga_signals.mult1_un75_sum_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_14_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_14_17_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_14_17_4  (
            .in0(N__13120),
            .in1(N__13200),
            .in2(_gnd_net_),
            .in3(N__12187),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_ns_1_LC_14_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_ns_1_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_ns_1_LC_14_17_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_ns_1_LC_14_17_7  (
            .in0(N__13201),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12147),
            .lcout(\this_vga_signals.mult1_un82_sum_c3_0_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_14_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_14_18_0 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_14_18_0  (
            .in0(N__11836),
            .in1(_gnd_net_),
            .in2(N__13037),
            .in3(N__12487),
            .lcout(\this_vga_signals.mult1_un61_sum_axb2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_14_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_14_18_2 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_14_18_2  (
            .in0(N__13026),
            .in1(N__13445),
            .in2(_gnd_net_),
            .in3(N__13220),
            .lcout(\this_vga_signals.mult1_un54_sum_c2 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_14_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_14_18_3 .LUT_INIT=16'b1011110101000010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_14_18_3  (
            .in0(N__13221),
            .in1(N__13281),
            .in2(N__11846),
            .in3(N__13258),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_14_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_14_18_4 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_14_18_4  (
            .in0(N__13028),
            .in1(_gnd_net_),
            .in2(N__11843),
            .in3(N__13115),
            .lcout(\this_vga_signals.mult1_un61_sum_c2 ),
            .ltout(\this_vga_signals.mult1_un61_sum_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_14_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_14_18_5 .LUT_INIT=16'b0110110011001001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_14_18_5  (
            .in0(N__12488),
            .in1(N__12502),
            .in2(N__11840),
            .in3(N__12520),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_0_LC_14_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_0_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_0_LC_14_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_0_LC_14_18_6  (
            .in0(N__13032),
            .in1(N__13116),
            .in2(_gnd_net_),
            .in3(N__12489),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_14_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_14_18_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__13027),
            .in2(_gnd_net_),
            .in3(N__11835),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI48605_9_LC_14_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI48605_9_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI48605_9_LC_14_19_1 .LUT_INIT=16'b0011111110011101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI48605_9_LC_14_19_1  (
            .in0(N__13335),
            .in1(N__13817),
            .in2(N__11870),
            .in3(N__12004),
            .lcout(\this_vga_signals.SUM_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_0_3_LC_14_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_0_3_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_0_3_LC_14_19_2 .LUT_INIT=16'b1000111110011111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_0_3_LC_14_19_2  (
            .in0(N__15070),
            .in1(N__15456),
            .in2(N__12776),
            .in3(N__13805),
            .lcout(\this_vga_signals.mult1_un47_sum_axb2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_14_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_14_19_3 .LUT_INIT=16'b0110011100001110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_14_19_3  (
            .in0(N__13018),
            .in1(N__13428),
            .in2(N__12807),
            .in3(N__15071),
            .lcout(\this_vga_signals.mult1_un47_sum_c2 ),
            .ltout(\this_vga_signals.mult1_un47_sum_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_0_LC_14_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_0_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_0_LC_14_19_4 .LUT_INIT=16'b0111100000111100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_0_LC_14_19_4  (
            .in0(N__11885),
            .in1(N__11912),
            .in2(N__11900),
            .in3(N__15457),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI87V41_6_LC_14_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI87V41_6_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI87V41_6_LC_14_19_5 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI87V41_6_LC_14_19_5  (
            .in0(N__13017),
            .in1(N__15069),
            .in2(_gnd_net_),
            .in3(N__13427),
            .lcout(\this_vga_signals.vaddress_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_4_tz_LC_14_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_4_tz_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_4_tz_LC_14_19_6 .LUT_INIT=16'b1101111111110111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_4_tz_LC_14_19_6  (
            .in0(N__15072),
            .in1(N__13806),
            .in2(N__13738),
            .in3(N__13336),
            .lcout(\this_vga_signals.mult1_un47_sum_axb2_3_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI94581_6_LC_14_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI94581_6_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI94581_6_LC_14_20_1 .LUT_INIT=16'b1110110000010011;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNI94581_6_LC_14_20_1  (
            .in0(N__13425),
            .in1(N__15391),
            .in2(N__13034),
            .in3(N__13722),
            .lcout(\this_vga_signals.vaddress_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_1_6_LC_14_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_1_6_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_1_6_LC_14_20_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_1_6_LC_14_20_2  (
            .in0(N__13721),
            .in1(N__15447),
            .in2(N__15068),
            .in3(N__13794),
            .lcout(\this_vga_signals.vaddress_c5_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_20_3 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_14_20_3  (
            .in0(N__12742),
            .in1(N__13080),
            .in2(N__12712),
            .in3(N__13192),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_d7lt8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBJQP3_6_LC_14_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBJQP3_6_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBJQP3_6_LC_14_20_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIBJQP3_6_LC_14_20_4  (
            .in0(N__15050),
            .in1(N__12014),
            .in2(N__11849),
            .in3(N__13795),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_d7lt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI8MOD6_9_LC_14_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI8MOD6_9_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI8MOD6_9_LC_14_20_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI8MOD6_9_LC_14_20_5  (
            .in0(N__12916),
            .in1(N__13337),
            .in2(N__12017),
            .in3(N__12765),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNI8MOD6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI0IM71_5_LC_14_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI0IM71_5_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI0IM71_5_LC_14_20_7 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI0IM71_5_LC_14_20_7  (
            .in0(N__13426),
            .in1(_gnd_net_),
            .in2(N__13035),
            .in3(N__13723),
            .lcout(\this_vga_signals.M_vcounter_d7lto8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_0_6_LC_14_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_0_6_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_0_6_LC_14_21_2 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_0_6_LC_14_21_2  (
            .in0(N__15458),
            .in1(N__13796),
            .in2(N__15083),
            .in3(N__13727),
            .lcout(),
            .ltout(\this_vga_signals.un6_vvisibilitylt9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR31O3_9_LC_14_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR31O3_9_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR31O3_9_LC_14_21_3 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIR31O3_9_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__13329),
            .in2(N__12008),
            .in3(N__12005),
            .lcout(\this_vga_signals.vvisibility ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_a5_1_0_LC_14_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_a5_1_0_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_a5_1_0_LC_14_21_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_a5_1_0_LC_14_21_4  (
            .in0(N__13330),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13797),
            .lcout(),
            .ltout(\this_vga_signals.vsync_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIP8HU1_6_LC_14_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIP8HU1_6_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIP8HU1_6_LC_14_21_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIP8HU1_6_LC_14_21_5  (
            .in0(N__13181),
            .in1(N__15082),
            .in2(N__11948),
            .in3(N__13010),
            .lcout(\this_vga_signals.vsync_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIRHPK7_9_LC_14_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIRHPK7_9_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIRHPK7_9_LC_14_21_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIRHPK7_9_LC_14_21_6  (
            .in0(N__14931),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12917),
            .lcout(\this_vga_signals.N_550_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_14_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_14_22_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_14_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_4_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13370),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21607),
            .ce(N__14990),
            .sr(N__14957));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_ns_LC_15_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_ns_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_ns_LC_15_17_2 .LUT_INIT=16'b1110100000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_ns_LC_15_17_2  (
            .in0(N__12743),
            .in1(N__12353),
            .in2(N__12719),
            .in3(N__11939),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_address_buffer_q_esr_7_LC_15_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_7_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_7_LC_15_17_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_7_LC_15_17_3  (
            .in0(N__12656),
            .in1(N__12527),
            .in2(N__12650),
            .in3(N__12191),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21579),
            .ce(N__15329),
            .sr(N__15216));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_ac0_3_0_LC_15_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_ac0_3_0_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_ac0_3_0_LC_15_17_5 .LUT_INIT=16'b1100010011011100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_ac0_3_0_LC_15_17_5  (
            .in0(N__13196),
            .in1(N__12536),
            .in2(N__12717),
            .in3(N__12148),
            .lcout(\this_vga_signals.mult1_un75_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un75_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_i_1_3_LC_15_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_i_1_3_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_i_1_3_LC_15_17_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_i_1_3_LC_15_17_6  (
            .in0(N__13113),
            .in1(N__13197),
            .in2(N__12530),
            .in3(N__12164),
            .lcout(\this_vga_signals.mult1_un82_sum_i_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_address_buffer_q_esr_10_LC_15_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_10_LC_15_18_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_10_LC_15_18_0 .LUT_INIT=16'b1000011100011110;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_10_LC_15_18_0  (
            .in0(N__12521),
            .in1(N__12331),
            .in2(N__12509),
            .in3(N__12491),
            .lcout(M_this_vga_signals_address_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21582),
            .ce(N__15327),
            .sr(N__15193));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_bm_LC_15_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_bm_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_bm_LC_15_18_2 .LUT_INIT=16'b0110110011001001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_c3_0_bm_LC_15_18_2  (
            .in0(N__13194),
            .in1(N__12199),
            .in2(N__13122),
            .in3(N__12188),
            .lcout(\this_vga_signals.mult1_un82_sum_c3_0_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_address_buffer_q_esr_9_LC_15_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_9_LC_15_18_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_9_LC_15_18_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_9_LC_15_18_3  (
            .in0(N__12190),
            .in1(N__12347),
            .in2(N__12335),
            .in3(N__12317),
            .lcout(M_this_vga_signals_address_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21582),
            .ce(N__15327),
            .sr(N__15193));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_LC_15_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_LC_15_18_4 .LUT_INIT=16'b0110001100111001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc2_LC_15_18_4  (
            .in0(N__13195),
            .in1(N__12200),
            .in2(N__13123),
            .in3(N__12189),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc2 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_address_buffer_q_esr_8_LC_15_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_8_LC_15_18_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_8_LC_15_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_8_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__12158),
            .in2(N__12152),
            .in3(N__12149),
            .lcout(M_this_vga_signals_address_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21582),
            .ce(N__15327),
            .sr(N__15193));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_15_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_15_19_0 .LUT_INIT=16'b1111111100011000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_15_19_0  (
            .in0(N__15445),
            .in1(N__15384),
            .in2(N__15409),
            .in3(N__15340),
            .lcout(\this_vga_signals.mult1_un40_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un40_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_15_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_15_19_1 .LUT_INIT=16'b0101101001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_15_19_1  (
            .in0(N__15073),
            .in1(N__13019),
            .in2(N__12785),
            .in3(N__13424),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_15_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_15_19_2 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_15_19_2  (
            .in0(N__13717),
            .in1(N__13332),
            .in2(N__13808),
            .in3(N__15383),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_x0_LC_15_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_x0_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_x0_LC_15_19_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_x0_LC_15_19_3  (
            .in0(N__15382),
            .in1(N__13799),
            .in2(_gnd_net_),
            .in3(N__13716),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a2_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_ns_LC_15_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_ns_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_ns_LC_15_19_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_ns_LC_15_19_4  (
            .in0(N__13423),
            .in1(_gnd_net_),
            .in2(N__12782),
            .in3(N__13664),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a2_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_3_LC_15_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_3_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_3_LC_15_19_5 .LUT_INIT=16'b1111001011110100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_3_LC_15_19_5  (
            .in0(N__13333),
            .in1(N__13803),
            .in2(N__12779),
            .in3(N__13718),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_0_3_1_1_LC_15_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_0_3_1_1_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_0_3_1_1_LC_15_19_7 .LUT_INIT=16'b0100010010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axb2_0_3_1_1_LC_15_19_7  (
            .in0(N__13334),
            .in1(N__13804),
            .in2(_gnd_net_),
            .in3(N__13719),
            .lcout(\this_vga_signals.mult1_un47_sum_axb2_0_3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_15_20_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_0_LC_15_20_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_15_20_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_15_20_0  (
            .in0(N__12919),
            .in1(N__12738),
            .in2(N__12767),
            .in3(N__12766),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .clk(N__21588),
            .ce(),
            .sr(N__14932));
    defparam \this_vga_signals.M_vcounter_q_1_LC_15_20_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_1_LC_15_20_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_15_20_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_15_20_1  (
            .in0(N__12923),
            .in1(N__12690),
            .in2(_gnd_net_),
            .in3(N__12659),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .clk(N__21588),
            .ce(),
            .sr(N__14932));
    defparam \this_vga_signals.M_vcounter_q_2_LC_15_20_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_2_LC_15_20_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_15_20_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_15_20_2  (
            .in0(N__12920),
            .in1(N__13193),
            .in2(_gnd_net_),
            .in3(N__13127),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .clk(N__21588),
            .ce(),
            .sr(N__14932));
    defparam \this_vga_signals.M_vcounter_q_3_LC_15_20_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_3_LC_15_20_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_15_20_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_15_20_3  (
            .in0(N__12924),
            .in1(N__13086),
            .in2(_gnd_net_),
            .in3(N__13040),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .clk(N__21588),
            .ce(),
            .sr(N__14932));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_15_20_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_15_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(N__13020),
            .in2(_gnd_net_),
            .in3(N__12938),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_LC_15_20_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_5_LC_15_20_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_LC_15_20_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_LC_15_20_5  (
            .in0(N__12925),
            .in1(N__13438),
            .in2(_gnd_net_),
            .in3(N__12935),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .clk(N__21588),
            .ce(),
            .sr(N__14932));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_15_20_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_15_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__15067),
            .in2(_gnd_net_),
            .in3(N__12932),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_LC_15_20_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_7_LC_15_20_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_LC_15_20_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_LC_15_20_7  (
            .in0(N__12926),
            .in1(N__13728),
            .in2(_gnd_net_),
            .in3(N__12929),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .clk(N__21588),
            .ce(),
            .sr(N__14932));
    defparam \this_vga_signals.M_vcounter_q_8_LC_15_21_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_8_LC_15_21_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_LC_15_21_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_LC_15_21_0  (
            .in0(N__12918),
            .in1(N__13798),
            .in2(_gnd_net_),
            .in3(N__12812),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .clk(N__21591),
            .ce(),
            .sr(N__14936));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_0_LC_15_21_1 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_0_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_0_LC_15_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_0_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__20255),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_1_LC_15_21_2 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_1_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_1_LC_15_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_1_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__20316),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_0_THRU_CO ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_2_LC_15_21_3 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_2_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_2_LC_15_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_2_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__20259),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_1_THRU_CO ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_3_LC_15_21_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_3_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_3_LC_15_21_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_3_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__20317),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_2_THRU_CO ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_4_LC_15_21_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_4_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_4_LC_15_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_4_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__20263),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_3_THRU_CO ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_5_LC_15_21_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_5_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_5_LC_15_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_5_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__20318),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_4_THRU_CO ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_6_LC_15_21_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_6_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_6_LC_15_21_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_THRU_CRY_6_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__20267),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_5_THRU_CO ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_15_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_15_22_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_15_22_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_9_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__13331),
            .in2(_gnd_net_),
            .in3(N__13340),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21599),
            .ce(N__15003),
            .sr(N__14965));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_2_9_LC_16_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_2_9_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_2_9_LC_16_17_0 .LUT_INIT=16'b0101101101111000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIUFPQ_2_9_LC_16_17_0  (
            .in0(N__14258),
            .in1(N__14102),
            .in2(N__14481),
            .in3(N__14608),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNIUFPQ_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_address_buffer_q_esr_11_LC_16_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_11_LC_16_18_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_11_LC_16_18_6 .LUT_INIT=16'b0011011010010011;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_11_LC_16_18_6  (
            .in0(N__13282),
            .in1(N__13262),
            .in2(N__13241),
            .in3(N__13229),
            .lcout(M_this_vga_signals_address_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21578),
            .ce(N__15328),
            .sr(N__15217));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_6_LC_16_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_6_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_6_LC_16_19_0 .LUT_INIT=16'b1100110011001001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIUQ9M1_6_LC_16_19_0  (
            .in0(N__15435),
            .in1(N__13807),
            .in2(N__15051),
            .in3(N__13720),
            .lcout(\this_vga_signals.vaddress_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_x1_LC_16_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_x1_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_x1_LC_16_20_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a2_x1_LC_16_20_5  (
            .in0(N__13354),
            .in1(N__13790),
            .in2(N__15381),
            .in3(N__13715),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a2_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam port_dmab_c_sbtinv_LC_16_20_6.C_ON=1'b0;
    defparam port_dmab_c_sbtinv_LC_16_20_6.SEQ_MODE=4'b0000;
    defparam port_dmab_c_sbtinv_LC_16_20_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 port_dmab_c_sbtinv_LC_16_20_6 (
            .in0(N__14861),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(port_dmab_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIP3JE_4_LC_16_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIP3JE_4_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIP3JE_4_LC_16_20_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIP3JE_4_LC_16_20_7  (
            .in0(N__13355),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13422),
            .lcout(\this_vga_signals.vaddress_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_16_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_16_21_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_16_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_6_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15097),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21587),
            .ce(N__15007),
            .sr(N__14966));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_16_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_16_21_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_16_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_4_LC_16_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13366),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21587),
            .ce(N__15007),
            .sr(N__14966));
    defparam M_this_data_count_q_0_LC_16_23_0.C_ON=1'b1;
    defparam M_this_data_count_q_0_LC_16_23_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_0_LC_16_23_0.LUT_INIT=16'b0011110000111100;
    LogicCell40 M_this_data_count_q_0_LC_16_23_0 (
            .in0(_gnd_net_),
            .in1(N__15641),
            .in2(N__20047),
            .in3(_gnd_net_),
            .lcout(M_this_data_count_qZ0Z_0),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(un1_M_this_data_count_q_cry_0),
            .clk(N__21595),
            .ce(),
            .sr(N__15482));
    defparam M_this_data_count_q_1_LC_16_23_1.C_ON=1'b1;
    defparam M_this_data_count_q_1_LC_16_23_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_1_LC_16_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_1_LC_16_23_1 (
            .in0(_gnd_net_),
            .in1(N__20011),
            .in2(N__15701),
            .in3(N__13346),
            .lcout(M_this_data_count_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_0),
            .carryout(un1_M_this_data_count_q_cry_1),
            .clk(N__21595),
            .ce(),
            .sr(N__15482));
    defparam M_this_data_count_q_2_LC_16_23_2.C_ON=1'b1;
    defparam M_this_data_count_q_2_LC_16_23_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_2_LC_16_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_2_LC_16_23_2 (
            .in0(_gnd_net_),
            .in1(N__15671),
            .in2(N__20048),
            .in3(N__13343),
            .lcout(M_this_data_count_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_1),
            .carryout(un1_M_this_data_count_q_cry_2),
            .clk(N__21595),
            .ce(),
            .sr(N__15482));
    defparam M_this_data_count_q_3_LC_16_23_3.C_ON=1'b1;
    defparam M_this_data_count_q_3_LC_16_23_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_3_LC_16_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_3_LC_16_23_3 (
            .in0(_gnd_net_),
            .in1(N__20015),
            .in2(N__15716),
            .in3(N__13847),
            .lcout(M_this_data_count_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_2),
            .carryout(un1_M_this_data_count_q_cry_3),
            .clk(N__21595),
            .ce(),
            .sr(N__15482));
    defparam M_this_data_count_q_4_LC_16_23_4.C_ON=1'b1;
    defparam M_this_data_count_q_4_LC_16_23_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_4_LC_16_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_4_LC_16_23_4 (
            .in0(_gnd_net_),
            .in1(N__15557),
            .in2(N__20049),
            .in3(N__13844),
            .lcout(M_this_data_count_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_3),
            .carryout(un1_M_this_data_count_q_cry_4),
            .clk(N__21595),
            .ce(),
            .sr(N__15482));
    defparam M_this_data_count_q_5_LC_16_23_5.C_ON=1'b1;
    defparam M_this_data_count_q_5_LC_16_23_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_5_LC_16_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_5_LC_16_23_5 (
            .in0(_gnd_net_),
            .in1(N__20019),
            .in2(N__15590),
            .in3(N__13841),
            .lcout(M_this_data_count_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_4),
            .carryout(un1_M_this_data_count_q_cry_5),
            .clk(N__21595),
            .ce(),
            .sr(N__15482));
    defparam M_this_data_count_q_6_LC_16_23_6.C_ON=1'b1;
    defparam M_this_data_count_q_6_LC_16_23_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_6_LC_16_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_6_LC_16_23_6 (
            .in0(_gnd_net_),
            .in1(N__15602),
            .in2(N__20050),
            .in3(N__13838),
            .lcout(M_this_data_count_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_5),
            .carryout(un1_M_this_data_count_q_cry_6),
            .clk(N__21595),
            .ce(),
            .sr(N__15482));
    defparam M_this_data_count_q_7_LC_16_23_7.C_ON=1'b1;
    defparam M_this_data_count_q_7_LC_16_23_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_7_LC_16_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_7_LC_16_23_7 (
            .in0(_gnd_net_),
            .in1(N__20023),
            .in2(N__15575),
            .in3(N__13835),
            .lcout(M_this_data_count_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_6),
            .carryout(un1_M_this_data_count_q_cry_7),
            .clk(N__21595),
            .ce(),
            .sr(N__15482));
    defparam M_this_data_count_q_8_LC_16_24_0.C_ON=1'b1;
    defparam M_this_data_count_q_8_LC_16_24_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_8_LC_16_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_8_LC_16_24_0 (
            .in0(_gnd_net_),
            .in1(N__15527),
            .in2(N__20051),
            .in3(N__13832),
            .lcout(M_this_data_count_qZ0Z_8),
            .ltout(),
            .carryin(bfn_16_24_0_),
            .carryout(un1_M_this_data_count_q_cry_8),
            .clk(N__21604),
            .ce(),
            .sr(N__15478));
    defparam M_this_data_count_q_9_LC_16_24_1.C_ON=1'b1;
    defparam M_this_data_count_q_9_LC_16_24_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_9_LC_16_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_9_LC_16_24_1 (
            .in0(_gnd_net_),
            .in1(N__15500),
            .in2(N__20054),
            .in3(N__13829),
            .lcout(M_this_data_count_qZ0Z_9),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_8),
            .carryout(un1_M_this_data_count_q_cry_9),
            .clk(N__21604),
            .ce(),
            .sr(N__15478));
    defparam M_this_data_count_q_10_LC_16_24_2.C_ON=1'b1;
    defparam M_this_data_count_q_10_LC_16_24_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_10_LC_16_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_10_LC_16_24_2 (
            .in0(_gnd_net_),
            .in1(N__15539),
            .in2(N__20052),
            .in3(N__13826),
            .lcout(M_this_data_count_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_9),
            .carryout(un1_M_this_data_count_q_cry_10),
            .clk(N__21604),
            .ce(),
            .sr(N__15478));
    defparam M_this_data_count_q_11_LC_16_24_3.C_ON=1'b1;
    defparam M_this_data_count_q_11_LC_16_24_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_11_LC_16_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_11_LC_16_24_3 (
            .in0(_gnd_net_),
            .in1(N__15514),
            .in2(N__20055),
            .in3(N__13823),
            .lcout(M_this_data_count_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_10),
            .carryout(un1_M_this_data_count_q_cry_11),
            .clk(N__21604),
            .ce(),
            .sr(N__15478));
    defparam M_this_data_count_q_12_LC_16_24_4.C_ON=1'b1;
    defparam M_this_data_count_q_12_LC_16_24_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_12_LC_16_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_12_LC_16_24_4 (
            .in0(_gnd_net_),
            .in1(N__15685),
            .in2(N__20053),
            .in3(N__13820),
            .lcout(M_this_data_count_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_11),
            .carryout(un1_M_this_data_count_q_cry_12),
            .clk(N__21604),
            .ce(),
            .sr(N__15478));
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_16_24_5.C_ON=1'b1;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_16_24_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_16_24_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_16_24_5 (
            .in0(_gnd_net_),
            .in1(N__20131),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_12),
            .carryout(un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_16_24_6.C_ON=1'b1;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_16_24_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_16_24_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_16_24_6 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__20181),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO),
            .carryout(un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_16_24_7.C_ON=1'b1;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_16_24_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_16_24_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_16_24_7 (
            .in0(_gnd_net_),
            .in1(N__20135),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO),
            .carryout(un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_13_LC_16_25_0.C_ON=1'b0;
    defparam M_this_data_count_q_13_LC_16_25_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_13_LC_16_25_0.LUT_INIT=16'b1110101110111110;
    LogicCell40 M_this_data_count_q_13_LC_16_25_0 (
            .in0(N__21761),
            .in1(N__20040),
            .in2(N__15659),
            .in3(N__14822),
            .lcout(M_this_data_count_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21614),
            .ce(),
            .sr(N__21340));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_1_c2_1_LC_17_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_1_c2_1_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_1_c2_1_LC_17_17_4 .LUT_INIT=16'b0101101101111000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_1_c2_1_LC_17_17_4  (
            .in0(N__14259),
            .in1(N__14118),
            .in2(N__14482),
            .in3(N__14609),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_1_c2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_1_c2_LC_17_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_1_c2_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_1_c2_LC_17_17_5 .LUT_INIT=16'b0101111100000101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_1_c2_LC_17_17_5  (
            .in0(N__14610),
            .in1(_gnd_net_),
            .in2(N__14819),
            .in3(N__14812),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_1_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum1_i_1_3_LC_17_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum1_i_1_3_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum1_i_1_3_LC_17_17_6 .LUT_INIT=16'b0100001000101011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum1_i_1_3_LC_17_17_6  (
            .in0(N__14627),
            .in1(N__14119),
            .in2(N__14618),
            .in3(N__14611),
            .lcout(\this_vga_signals.mult1_un54_sum1_i_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_address_buffer_q_esr_5_LC_17_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_5_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_5_LC_17_18_1 .LUT_INIT=16'b1011001001001101;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_5_LC_17_18_1  (
            .in0(N__14477),
            .in1(N__14297),
            .in2(N__14126),
            .in3(N__13961),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21583),
            .ce(N__15317),
            .sr(N__15211));
    defparam \this_vga_signals.M_address_buffer_q_esr_13_LC_17_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_address_buffer_q_esr_13_LC_17_19_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_address_buffer_q_esr_13_LC_17_19_7 .LUT_INIT=16'b1111111100100100;
    LogicCell40 \this_vga_signals.M_address_buffer_q_esr_13_LC_17_19_7  (
            .in0(N__15446),
            .in1(N__15410),
            .in2(N__15392),
            .in3(N__15344),
            .lcout(M_this_vga_signals_address_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21584),
            .ce(N__15316),
            .sr(N__15215));
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_17_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_17_20_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_17_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_6_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15098),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21589),
            .ce(N__15011),
            .sr(N__14958));
    defparam \this_start_data_delay.M_last_q_RNI9P6N1_LC_17_21_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI9P6N1_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI9P6N1_LC_17_21_4 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \this_start_data_delay.M_last_q_RNI9P6N1_LC_17_21_4  (
            .in0(N__15978),
            .in1(N__21395),
            .in2(N__15740),
            .in3(N__19023),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_state_q_srsts_i_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_2_LC_17_21_5.C_ON=1'b0;
    defparam M_this_state_q_2_LC_17_21_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_2_LC_17_21_5.LUT_INIT=16'b0100000001110000;
    LogicCell40 M_this_state_q_2_LC_17_21_5 (
            .in0(N__15620),
            .in1(N__15979),
            .in2(N__14900),
            .in3(N__18771),
            .lcout(M_this_state_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21592),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_1_LC_17_22_0.C_ON=1'b0;
    defparam M_this_state_q_1_LC_17_22_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_1_LC_17_22_0.LUT_INIT=16'b0000000001001111;
    LogicCell40 M_this_state_q_1_LC_17_22_0 (
            .in0(N__15616),
            .in1(N__15739),
            .in2(N__14897),
            .in3(N__21389),
            .lcout(M_this_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21600),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_0_1_1_LC_17_22_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_0_1_1_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_0_1_1_LC_17_22_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_i_a2_0_1_1_LC_17_22_4  (
            .in0(N__21747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19996),
            .lcout(\this_start_data_delay.N_389_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.dma_i_a2_LC_17_22_5 .C_ON=1'b0;
    defparam \this_start_data_delay.dma_i_a2_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.dma_i_a2_LC_17_22_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_start_data_delay.dma_i_a2_LC_17_22_5  (
            .in0(N__19995),
            .in1(N__15975),
            .in2(_gnd_net_),
            .in3(N__19014),
            .lcout(port_dmab_c),
            .ltout(port_dmab_c_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI7S6U1_LC_17_22_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI7S6U1_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI7S6U1_LC_17_22_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI7S6U1_LC_17_22_6  (
            .in0(N__21746),
            .in1(N__21387),
            .in2(N__14828),
            .in3(N__18740),
            .lcout(),
            .ltout(\this_start_data_delay.N_385_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNINC2J4_LC_17_22_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNINC2J4_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNINC2J4_LC_17_22_7 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \this_start_data_delay.M_last_q_RNINC2J4_LC_17_22_7  (
            .in0(N__21388),
            .in1(N__15976),
            .in2(N__14825),
            .in3(N__15615),
            .lcout(\this_start_data_delay.M_this_state_q_srsts_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_9_1_LC_17_23_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_9_1_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_9_1_LC_17_23_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_i_a2_1_9_1_LC_17_23_0  (
            .in0(N__15712),
            .in1(N__15697),
            .in2(N__15686),
            .in3(N__15670),
            .lcout(\this_start_data_delay.M_this_state_q_srsts_i_a2_1_9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_6_1_LC_17_23_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_6_1_LC_17_23_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_6_1_LC_17_23_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_i_a2_1_6_1_LC_17_23_2  (
            .in0(_gnd_net_),
            .in1(N__15658),
            .in2(_gnd_net_),
            .in3(N__15640),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_state_q_srsts_i_a2_1_6Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_1_LC_17_23_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_1_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_1_LC_17_23_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_i_a2_1_1_LC_17_23_3  (
            .in0(N__15629),
            .in1(N__15545),
            .in2(N__15623),
            .in3(N__15488),
            .lcout(\this_start_data_delay.N_413 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_8_1_LC_17_23_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_8_1_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_8_1_LC_17_23_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_i_a2_1_8_1_LC_17_23_6  (
            .in0(N__15601),
            .in1(N__15586),
            .in2(N__15574),
            .in3(N__15556),
            .lcout(\this_start_data_delay.M_this_state_q_srsts_i_a2_1_8Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_7_1_LC_17_24_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_7_1_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_a2_1_7_1_LC_17_24_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_i_a2_1_7_1_LC_17_24_1  (
            .in0(N__15538),
            .in1(N__15526),
            .in2(N__15515),
            .in3(N__15499),
            .lcout(\this_start_data_delay.M_this_state_q_srsts_i_a2_1_7Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI20CE_0_LC_17_24_2.C_ON=1'b0;
    defparam M_this_state_q_RNI20CE_0_LC_17_24_2.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI20CE_0_LC_17_24_2.LUT_INIT=16'b1111111110101010;
    LogicCell40 M_this_state_q_RNI20CE_0_LC_17_24_2 (
            .in0(N__21727),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21393),
            .lcout(M_this_state_q_RNI20CEZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_17_25_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_17_25_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_17_25_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_17_25_0  (
            .in0(_gnd_net_),
            .in1(N__15798),
            .in2(_gnd_net_),
            .in3(N__15776),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21618),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_17_25_1 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_17_25_1 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_17_25_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_17_25_1  (
            .in0(N__15799),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15464),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21618),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_17_25_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_17_25_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_17_25_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_17_25_2  (
            .in0(_gnd_net_),
            .in1(N__15800),
            .in2(_gnd_net_),
            .in3(N__15806),
            .lcout(M_this_state_q_nss_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21618),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_17_25_3 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_17_25_3 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_17_25_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_17_25_3  (
            .in0(N__15797),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21618),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_0_LC_17_25_5.C_ON=1'b0;
    defparam M_this_state_q_0_LC_17_25_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_0_LC_17_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_state_q_0_LC_17_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15766),
            .lcout(M_this_state_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21618),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_11_LC_18_21_5.C_ON=1'b0;
    defparam M_this_internal_address_q_11_LC_18_21_5.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_11_LC_18_21_5.LUT_INIT=16'b0101001101010000;
    LogicCell40 M_this_internal_address_q_11_LC_18_21_5 (
            .in0(N__15722),
            .in1(N__21782),
            .in2(N__18051),
            .in3(N__17471),
            .lcout(M_this_internal_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21601),
            .ce(),
            .sr(N__21342));
    defparam \this_start_data_delay.M_this_state_q_srsts_0_a2_1_0_4_LC_18_22_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_a2_1_0_4_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_a2_1_0_4_LC_18_22_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_0_a2_1_0_4_LC_18_22_0  (
            .in0(N__15946),
            .in1(N__21394),
            .in2(N__20039),
            .in3(N__19015),
            .lcout(\this_start_data_delay.M_this_state_q_srsts_0_a2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_4_LC_18_22_1 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_4_LC_18_22_1 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_4_LC_18_22_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_delay_clk.M_pipe_q_4_LC_18_22_1  (
            .in0(_gnd_net_),
            .in1(N__15749),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_delay_clk_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21608),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI8LQ11_LC_18_22_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI8LQ11_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI8LQ11_LC_18_22_2 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI8LQ11_LC_18_22_2  (
            .in0(N__15853),
            .in1(N__15876),
            .in2(N__15839),
            .in3(N__15977),
            .lcout(\this_start_data_delay.N_353_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_LC_18_22_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_LC_18_22_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_LC_18_22_3 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIBJQQ_LC_18_22_3  (
            .in0(N__15877),
            .in1(N__15834),
            .in2(_gnd_net_),
            .in3(N__15851),
            .lcout(M_this_start_data_delay_out_0),
            .ltout(M_this_start_data_delay_out_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_11_LC_18_22_4 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_11_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_11_LC_18_22_4 .LUT_INIT=16'b0100000001111111;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_11_LC_18_22_4  (
            .in0(N__18938),
            .in1(N__17737),
            .in2(N__15725),
            .in3(N__20634),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNICHCU_LC_18_22_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNICHCU_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNICHCU_LC_18_22_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_start_data_delay.M_last_q_RNICHCU_LC_18_22_5  (
            .in0(N__15878),
            .in1(N__15835),
            .in2(N__15920),
            .in3(N__15852),
            .lcout(\this_start_data_delay.N_352_0 ),
            .ltout(\this_start_data_delay.N_352_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_4_LC_18_22_6.C_ON=1'b0;
    defparam M_this_state_q_4_LC_18_22_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_4_LC_18_22_6.LUT_INIT=16'b1000110011111111;
    LogicCell40 M_this_state_q_4_LC_18_22_6 (
            .in0(N__16073),
            .in1(N__15896),
            .in2(N__15890),
            .in3(N__15887),
            .lcout(M_this_state_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21608),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_LC_18_22_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_LC_18_22_7 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.M_last_q_LC_18_22_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.M_last_q_LC_18_22_7  (
            .in0(N__15875),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15854),
            .lcout(\this_start_data_delay.M_last_qZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21608),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIILOC1_LC_18_23_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIILOC1_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIILOC1_LC_18_23_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIILOC1_LC_18_23_3  (
            .in0(N__15824),
            .in1(N__15945),
            .in2(_gnd_net_),
            .in3(N__21391),
            .lcout(\this_start_data_delay.N_398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_4_LC_18_23_4 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_4_LC_18_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_4_LC_18_23_4 .LUT_INIT=16'b0100011101010101;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_4_LC_18_23_4  (
            .in0(N__16896),
            .in1(N__17722),
            .in2(N__18937),
            .in3(N__18761),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_1_LC_18_24_2 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_1_LC_18_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_1_LC_18_24_2 .LUT_INIT=16'b0000001011011111;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_1_LC_18_24_2  (
            .in0(N__18791),
            .in1(N__17721),
            .in2(N__18270),
            .in3(N__16290),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIHI621_LC_18_24_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIHI621_LC_18_24_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIHI621_LC_18_24_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_start_data_delay.M_last_q_RNIHI621_LC_18_24_5  (
            .in0(_gnd_net_),
            .in1(N__21392),
            .in2(_gnd_net_),
            .in3(N__18790),
            .lcout(\this_start_data_delay.N_407 ),
            .ltout(\this_start_data_delay.N_407_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_6_LC_18_24_6.C_ON=1'b0;
    defparam M_this_state_q_6_LC_18_24_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_6_LC_18_24_6.LUT_INIT=16'b1110101011000000;
    LogicCell40 M_this_state_q_6_LC_18_24_6 (
            .in0(N__16001),
            .in1(N__15995),
            .in2(N__15818),
            .in3(N__16092),
            .lcout(M_this_state_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21619),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_1_LC_18_25_0.C_ON=1'b0;
    defparam M_this_internal_address_q_1_LC_18_25_0.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_1_LC_18_25_0.LUT_INIT=16'b0001110100001100;
    LogicCell40 M_this_internal_address_q_1_LC_18_25_0 (
            .in0(N__21718),
            .in1(N__18013),
            .in2(N__15815),
            .in3(N__16271),
            .lcout(M_this_internal_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21624),
            .ce(),
            .sr(N__21341));
    defparam \this_start_data_delay.M_this_internal_address_q_3s2_LC_18_25_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_internal_address_q_3s2_LC_18_25_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_internal_address_q_3s2_LC_18_25_7 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \this_start_data_delay.M_this_internal_address_q_3s2_LC_18_25_7  (
            .in0(N__15994),
            .in1(N__17726),
            .in2(_gnd_net_),
            .in3(N__21717),
            .lcout(M_this_internal_address_q_3_sm0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_5_LC_19_20_2 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_5_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_5_LC_19_20_2 .LUT_INIT=16'b0000001011011111;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_5_LC_19_20_2  (
            .in0(N__18793),
            .in1(N__17746),
            .in2(N__18226),
            .in3(N__16765),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_7_LC_19_20_3 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_7_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_7_LC_19_20_3 .LUT_INIT=16'b0001101100110011;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_7_LC_19_20_3  (
            .in0(N__17748),
            .in1(N__16632),
            .in2(N__18980),
            .in3(N__18794),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_3_LC_19_20_7 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_3_LC_19_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_3_LC_19_20_7 .LUT_INIT=16'b0010011100110011;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_3_LC_19_20_7  (
            .in0(N__17747),
            .in1(N__17035),
            .in2(N__19520),
            .in3(N__18792),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_13_LC_19_21_0 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_13_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_13_LC_19_21_0 .LUT_INIT=16'b0001101100110011;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_13_LC_19_21_0  (
            .in0(N__17734),
            .in1(N__20550),
            .in2(N__20942),
            .in3(N__18738),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_12_LC_19_21_2 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_12_LC_19_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_12_LC_19_21_2 .LUT_INIT=16'b0001101100110011;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_12_LC_19_21_2  (
            .in0(N__17735),
            .in1(N__20730),
            .in2(N__18227),
            .in3(N__18737),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI95RM1_LC_19_21_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI95RM1_LC_19_21_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI95RM1_LC_19_21_4 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \this_start_data_delay.M_last_q_RNI95RM1_LC_19_21_4  (
            .in0(N__15983),
            .in1(N__18683),
            .in2(N__15947),
            .in3(N__18736),
            .lcout(N_346_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_9_LC_19_21_6 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_9_LC_19_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_9_LC_19_21_6 .LUT_INIT=16'b0001101100110011;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_9_LC_19_21_6  (
            .in0(N__17736),
            .in1(N__16497),
            .in2(N__20977),
            .in3(N__18739),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_4_LC_19_22_3.C_ON=1'b0;
    defparam M_this_internal_address_q_4_LC_19_22_3.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_4_LC_19_22_3.LUT_INIT=16'b0011010100110000;
    LogicCell40 M_this_internal_address_q_4_LC_19_22_3 (
            .in0(N__21836),
            .in1(N__15926),
            .in2(N__18082),
            .in3(N__16877),
            .lcout(M_this_internal_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21616),
            .ce(),
            .sr(N__21343));
    defparam M_this_internal_address_q_2_LC_19_22_4.C_ON=1'b0;
    defparam M_this_internal_address_q_2_LC_19_22_4.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_2_LC_19_22_4.LUT_INIT=16'b0101010100110000;
    LogicCell40 M_this_internal_address_q_2_LC_19_22_4 (
            .in0(N__16112),
            .in1(N__21838),
            .in2(N__16133),
            .in3(N__18069),
            .lcout(M_this_internal_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21616),
            .ce(),
            .sr(N__21343));
    defparam M_this_internal_address_q_9_LC_19_22_7.C_ON=1'b0;
    defparam M_this_internal_address_q_9_LC_19_22_7.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_9_LC_19_22_7.LUT_INIT=16'b0011010100110000;
    LogicCell40 M_this_internal_address_q_9_LC_19_22_7 (
            .in0(N__21837),
            .in1(N__16118),
            .in2(N__18083),
            .in3(N__16478),
            .lcout(M_this_internal_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21616),
            .ce(),
            .sr(N__21343));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_10_LC_19_23_0 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_10_LC_19_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_10_LC_19_23_0 .LUT_INIT=16'b0001101100110011;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_10_LC_19_23_0  (
            .in0(N__17719),
            .in1(N__17196),
            .in2(N__19519),
            .in3(N__18762),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_2_LC_19_23_2 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_2_LC_19_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_2_LC_19_23_2 .LUT_INIT=16'b0010011100110011;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_2_LC_19_23_2  (
            .in0(N__17720),
            .in1(N__16152),
            .in2(N__20984),
            .in3(N__18763),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_5_LC_19_24_2.C_ON=1'b0;
    defparam M_this_state_q_5_LC_19_24_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_5_LC_19_24_2.LUT_INIT=16'b1110101011000000;
    LogicCell40 M_this_state_q_5_LC_19_24_2 (
            .in0(N__16061),
            .in1(N__16105),
            .in2(N__17745),
            .in3(N__16093),
            .lcout(M_this_state_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21625),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_7_LC_19_24_6.C_ON=1'b0;
    defparam M_this_state_q_7_LC_19_24_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_7_LC_19_24_6.LUT_INIT=16'b1110110010100000;
    LogicCell40 M_this_state_q_7_LC_19_24_6 (
            .in0(N__16106),
            .in1(N__16094),
            .in2(N__19053),
            .in3(N__16079),
            .lcout(M_this_state_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21625),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_d29_LC_19_25_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_d29_LC_19_25_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_d29_LC_19_25_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_start_data_delay.M_this_state_d29_LC_19_25_0  (
            .in0(N__17491),
            .in1(N__16023),
            .in2(N__16055),
            .in3(N__21201),
            .lcout(\this_start_data_delay.M_this_state_dZ0Z29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_0_a2_3_4_LC_19_25_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_a2_3_4_LC_19_25_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_a2_3_4_LC_19_25_1 .LUT_INIT=16'b1000111111111111;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_0_a2_3_4_LC_19_25_1  (
            .in0(N__16053),
            .in1(N__16025),
            .in2(N__21206),
            .in3(N__17492),
            .lcout(\this_start_data_delay.N_396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_d27_LC_19_25_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_d27_LC_19_25_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_d27_LC_19_25_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_start_data_delay.M_this_state_d27_LC_19_25_6  (
            .in0(N__17489),
            .in1(N__16022),
            .in2(N__16054),
            .in3(N__21197),
            .lcout(\this_start_data_delay.M_this_state_dZ0Z27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_d28_LC_19_25_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_d28_LC_19_25_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_d28_LC_19_25_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_start_data_delay.M_this_state_d28_LC_19_25_7  (
            .in0(N__16052),
            .in1(N__16024),
            .in2(N__21205),
            .in3(N__17490),
            .lcout(\this_start_data_delay.M_this_state_dZ0Z28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_13_LC_20_19_0 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_13_LC_20_19_0 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_13_LC_20_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vram.mem_radreg_13_LC_20_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16466),
            .lcout(\this_vram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21602),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_12_LC_20_19_4 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_12_LC_20_19_4 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_12_LC_20_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vram.mem_radreg_12_LC_20_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16457),
            .lcout(\this_vram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21602),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_5_LC_20_20_2.C_ON=1'b0;
    defparam M_this_internal_address_q_5_LC_20_20_2.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_5_LC_20_20_2.LUT_INIT=16'b0101001101010000;
    LogicCell40 M_this_internal_address_q_5_LC_20_20_2 (
            .in0(N__16445),
            .in1(N__21857),
            .in2(N__18073),
            .in3(N__16745),
            .lcout(M_this_internal_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21609),
            .ce(),
            .sr(N__21346));
    defparam M_this_internal_address_q_3_LC_20_20_5.C_ON=1'b0;
    defparam M_this_internal_address_q_3_LC_20_20_5.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_3_LC_20_20_5.LUT_INIT=16'b0011001101010000;
    LogicCell40 M_this_internal_address_q_3_LC_20_20_5 (
            .in0(N__21856),
            .in1(N__16439),
            .in2(N__17012),
            .in3(N__18046),
            .lcout(M_this_internal_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21609),
            .ce(),
            .sr(N__21346));
    defparam M_this_internal_address_q_7_LC_20_20_6.C_ON=1'b0;
    defparam M_this_internal_address_q_7_LC_20_20_6.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_7_LC_20_20_6.LUT_INIT=16'b0001101100001010;
    LogicCell40 M_this_internal_address_q_7_LC_20_20_6 (
            .in0(N__18045),
            .in1(N__21858),
            .in2(N__16433),
            .in3(N__16613),
            .lcout(M_this_internal_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21609),
            .ce(),
            .sr(N__21346));
    defparam M_this_internal_address_q_0_LC_20_20_7.C_ON=1'b0;
    defparam M_this_internal_address_q_0_LC_20_20_7.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_0_LC_20_20_7.LUT_INIT=16'b0000111101000100;
    LogicCell40 M_this_internal_address_q_0_LC_20_20_7 (
            .in0(N__21855),
            .in1(N__16406),
            .in2(N__17324),
            .in3(N__18050),
            .lcout(M_this_internal_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21609),
            .ce(),
            .sr(N__21346));
    defparam M_this_internal_address_q_RNI6EA12_0_LC_20_21_0.C_ON=1'b1;
    defparam M_this_internal_address_q_RNI6EA12_0_LC_20_21_0.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNI6EA12_0_LC_20_21_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNI6EA12_0_LC_20_21_0 (
            .in0(_gnd_net_),
            .in1(N__17343),
            .in2(N__16421),
            .in3(N__16420),
            .lcout(M_this_internal_address_q_RNI6EA12Z0Z_0),
            .ltout(),
            .carryin(bfn_20_21_0_),
            .carryout(un1_M_this_internal_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_0_c_RNI4MQI_LC_20_21_1.C_ON=1'b1;
    defparam un1_M_this_internal_address_q_cry_0_c_RNI4MQI_LC_20_21_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_0_c_RNI4MQI_LC_20_21_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_internal_address_q_cry_0_c_RNI4MQI_LC_20_21_1 (
            .in0(_gnd_net_),
            .in1(N__16303),
            .in2(_gnd_net_),
            .in3(N__16259),
            .lcout(un1_M_this_internal_address_q_cry_0_c_RNI4MQIZ0),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_0),
            .carryout(un1_M_this_internal_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_1_c_RNI6PRI_LC_20_21_2.C_ON=1'b1;
    defparam un1_M_this_internal_address_q_cry_1_c_RNI6PRI_LC_20_21_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_1_c_RNI6PRI_LC_20_21_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_internal_address_q_cry_1_c_RNI6PRI_LC_20_21_2 (
            .in0(_gnd_net_),
            .in1(N__16153),
            .in2(_gnd_net_),
            .in3(N__16121),
            .lcout(un1_M_this_internal_address_q_cry_1_c_RNI6PRIZ0),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_1),
            .carryout(un1_M_this_internal_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_2_c_RNI8SSI_LC_20_21_3.C_ON=1'b1;
    defparam un1_M_this_internal_address_q_cry_2_c_RNI8SSI_LC_20_21_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_2_c_RNI8SSI_LC_20_21_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_internal_address_q_cry_2_c_RNI8SSI_LC_20_21_3 (
            .in0(_gnd_net_),
            .in1(N__17031),
            .in2(_gnd_net_),
            .in3(N__17003),
            .lcout(un1_M_this_internal_address_q_cry_2_c_RNI8SSIZ0),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_2),
            .carryout(un1_M_this_internal_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_3_c_RNIAVTI_LC_20_21_4.C_ON=1'b1;
    defparam un1_M_this_internal_address_q_cry_3_c_RNIAVTI_LC_20_21_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_3_c_RNIAVTI_LC_20_21_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_internal_address_q_cry_3_c_RNIAVTI_LC_20_21_4 (
            .in0(_gnd_net_),
            .in1(N__16897),
            .in2(_gnd_net_),
            .in3(N__16871),
            .lcout(un1_M_this_internal_address_q_cry_3_c_RNIAVTIZ0),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_3),
            .carryout(un1_M_this_internal_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_4_c_RNIC2VI_LC_20_21_5.C_ON=1'b1;
    defparam un1_M_this_internal_address_q_cry_4_c_RNIC2VI_LC_20_21_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_4_c_RNIC2VI_LC_20_21_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_internal_address_q_cry_4_c_RNIC2VI_LC_20_21_5 (
            .in0(_gnd_net_),
            .in1(N__16764),
            .in2(_gnd_net_),
            .in3(N__16739),
            .lcout(un1_M_this_internal_address_q_cry_4_c_RNIC2VIZ0),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_4),
            .carryout(un1_M_this_internal_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_5_c_RNIE50J_LC_20_21_6.C_ON=1'b1;
    defparam un1_M_this_internal_address_q_cry_5_c_RNIE50J_LC_20_21_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_5_c_RNIE50J_LC_20_21_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_internal_address_q_cry_5_c_RNIE50J_LC_20_21_6 (
            .in0(_gnd_net_),
            .in1(N__17775),
            .in2(_gnd_net_),
            .in3(N__16736),
            .lcout(un1_M_this_internal_address_q_cry_5_c_RNIE50JZ0),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_5),
            .carryout(un1_M_this_internal_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_6_c_RNIG81J_LC_20_21_7.C_ON=1'b1;
    defparam un1_M_this_internal_address_q_cry_6_c_RNIG81J_LC_20_21_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_6_c_RNIG81J_LC_20_21_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_internal_address_q_cry_6_c_RNIG81J_LC_20_21_7 (
            .in0(_gnd_net_),
            .in1(N__16633),
            .in2(_gnd_net_),
            .in3(N__16607),
            .lcout(un1_M_this_internal_address_q_cry_6_c_RNIG81JZ0),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_6),
            .carryout(un1_M_this_internal_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_7_c_RNIIB2J_LC_20_22_0.C_ON=1'b1;
    defparam un1_M_this_internal_address_q_cry_7_c_RNIIB2J_LC_20_22_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_7_c_RNIIB2J_LC_20_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_internal_address_q_cry_7_c_RNIIB2J_LC_20_22_0 (
            .in0(_gnd_net_),
            .in1(N__17539),
            .in2(_gnd_net_),
            .in3(N__16604),
            .lcout(un1_M_this_internal_address_q_cry_7_c_RNIIB2JZ0),
            .ltout(),
            .carryin(bfn_20_22_0_),
            .carryout(un1_M_this_internal_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_8_c_RNIKE3J_LC_20_22_1.C_ON=1'b1;
    defparam un1_M_this_internal_address_q_cry_8_c_RNIKE3J_LC_20_22_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_8_c_RNIKE3J_LC_20_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_internal_address_q_cry_8_c_RNIKE3J_LC_20_22_1 (
            .in0(_gnd_net_),
            .in1(N__16498),
            .in2(_gnd_net_),
            .in3(N__16472),
            .lcout(un1_M_this_internal_address_q_cry_8_c_RNIKE3JZ0),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_8),
            .carryout(un1_M_this_internal_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_9_c_RNITQCI_LC_20_22_2.C_ON=1'b1;
    defparam un1_M_this_internal_address_q_cry_9_c_RNITQCI_LC_20_22_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_9_c_RNITQCI_LC_20_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_internal_address_q_cry_9_c_RNITQCI_LC_20_22_2 (
            .in0(_gnd_net_),
            .in1(N__17197),
            .in2(_gnd_net_),
            .in3(N__16469),
            .lcout(un1_M_this_internal_address_q_cry_9_c_RNITQCIZ0),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_9),
            .carryout(un1_M_this_internal_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_10_c_RNI6I0D_LC_20_22_3.C_ON=1'b1;
    defparam un1_M_this_internal_address_q_cry_10_c_RNI6I0D_LC_20_22_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_10_c_RNI6I0D_LC_20_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_internal_address_q_cry_10_c_RNI6I0D_LC_20_22_3 (
            .in0(_gnd_net_),
            .in1(N__20663),
            .in2(_gnd_net_),
            .in3(N__17459),
            .lcout(un1_M_this_internal_address_q_cry_10_c_RNI6I0DZ0),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_10),
            .carryout(un1_M_this_internal_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_11_c_RNI8L1D_LC_20_22_4.C_ON=1'b1;
    defparam un1_M_this_internal_address_q_cry_11_c_RNI8L1D_LC_20_22_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_11_c_RNI8L1D_LC_20_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_internal_address_q_cry_11_c_RNI8L1D_LC_20_22_4 (
            .in0(_gnd_net_),
            .in1(N__20712),
            .in2(_gnd_net_),
            .in3(N__17456),
            .lcout(un1_M_this_internal_address_q_cry_11_c_RNI8L1DZ0),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_11),
            .carryout(un1_M_this_internal_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_internal_address_q_cry_12_c_RNIAO2D_LC_20_22_5.C_ON=1'b0;
    defparam un1_M_this_internal_address_q_cry_12_c_RNIAO2D_LC_20_22_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_internal_address_q_cry_12_c_RNIAO2D_LC_20_22_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_M_this_internal_address_q_cry_12_c_RNIAO2D_LC_20_22_5 (
            .in0(_gnd_net_),
            .in1(N__20526),
            .in2(_gnd_net_),
            .in3(N__17453),
            .lcout(un1_M_this_internal_address_q_cry_12_c_RNIAO2DZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_0_LC_20_22_6 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_0_LC_20_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_0_LC_20_22_6 .LUT_INIT=16'b0001101100001111;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_0_LC_20_22_6  (
            .in0(N__17741),
            .in1(N__18975),
            .in2(N__17356),
            .in3(N__18783),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_10_LC_20_23_5.C_ON=1'b0;
    defparam M_this_internal_address_q_10_LC_20_23_5.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_10_LC_20_23_5.LUT_INIT=16'b0101001101010000;
    LogicCell40 M_this_internal_address_q_10_LC_20_23_5 (
            .in0(N__17312),
            .in1(N__21835),
            .in2(N__18080),
            .in3(N__17306),
            .lcout(M_this_internal_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21626),
            .ce(),
            .sr(N__21344));
    defparam M_this_internal_address_q_12_LC_21_21_1.C_ON=1'b0;
    defparam M_this_internal_address_q_12_LC_21_21_1.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_12_LC_21_21_1.LUT_INIT=16'b0101001101010000;
    LogicCell40 M_this_internal_address_q_12_LC_21_21_1 (
            .in0(N__17177),
            .in1(N__21859),
            .in2(N__18085),
            .in3(N__17168),
            .lcout(M_this_internal_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21620),
            .ce(),
            .sr(N__21347));
    defparam M_this_internal_address_q_6_LC_21_21_5.C_ON=1'b0;
    defparam M_this_internal_address_q_6_LC_21_21_5.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_6_LC_21_21_5.LUT_INIT=16'b0101001101010000;
    LogicCell40 M_this_internal_address_q_6_LC_21_21_5 (
            .in0(N__17756),
            .in1(N__21860),
            .in2(N__18086),
            .in3(N__17162),
            .lcout(M_this_internal_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21620),
            .ce(),
            .sr(N__21347));
    defparam M_this_internal_address_q_13_LC_21_22_0.C_ON=1'b0;
    defparam M_this_internal_address_q_13_LC_21_22_0.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_13_LC_21_22_0.LUT_INIT=16'b0101001101010000;
    LogicCell40 M_this_internal_address_q_13_LC_21_22_0 (
            .in0(N__17156),
            .in1(N__21820),
            .in2(N__18081),
            .in3(N__17144),
            .lcout(M_this_internal_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21627),
            .ce(),
            .sr(N__21345));
    defparam M_this_internal_address_q_8_LC_21_22_1.C_ON=1'b0;
    defparam M_this_internal_address_q_8_LC_21_22_1.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_8_LC_21_22_1.LUT_INIT=16'b0000010011110100;
    LogicCell40 M_this_internal_address_q_8_LC_21_22_1 (
            .in0(N__21819),
            .in1(N__17138),
            .in2(N__18084),
            .in3(N__17519),
            .lcout(M_this_internal_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21627),
            .ce(),
            .sr(N__21345));
    defparam M_this_state_q_3_LC_21_22_3.C_ON=1'b0;
    defparam M_this_state_q_3_LC_21_22_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_3_LC_21_22_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 M_this_state_q_3_LC_21_22_3 (
            .in0(_gnd_net_),
            .in1(N__19030),
            .in2(_gnd_net_),
            .in3(N__18798),
            .lcout(M_this_state_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21627),
            .ce(),
            .sr(N__21345));
    defparam \this_vram.mem_mem_0_0_RNIQOI11_0_LC_22_17_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_0_LC_22_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_0_LC_22_17_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_0_0_RNIQOI11_0_LC_22_17_1  (
            .in0(N__19618),
            .in1(N__17972),
            .in2(_gnd_net_),
            .in3(N__17963),
            .lcout(),
            .ltout(\this_vram.mem_mem_0_0_RNIQOI11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI95PB2_11_LC_22_17_2 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI95PB2_11_LC_22_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI95PB2_11_LC_22_17_2 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \this_vram.mem_radreg_RNI95PB2_11_LC_22_17_2  (
            .in0(N__18363),
            .in1(N__19212),
            .in2(N__17948),
            .in3(N__18512),
            .lcout(\this_vram.mem_DOUT_7_i_m2_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_11_LC_22_18_3 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_11_LC_22_18_3 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_11_LC_22_18_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_vram.mem_radreg_11_LC_22_18_3  (
            .in0(_gnd_net_),
            .in1(N__17945),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21610),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIDSEJ4_11_LC_22_18_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIDSEJ4_11_LC_22_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIDSEJ4_11_LC_22_18_6 .LUT_INIT=16'b1010000011001111;
    LogicCell40 \this_vram.mem_radreg_RNIDSEJ4_11_LC_22_18_6  (
            .in0(N__19775),
            .in1(N__18473),
            .in2(N__18365),
            .in3(N__17936),
            .lcout(M_this_vram_read_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_6_LC_22_21_7 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_6_LC_22_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_6_LC_22_21_7 .LUT_INIT=16'b0010011100110011;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_6_LC_22_21_7  (
            .in0(N__17749),
            .in1(N__17776),
            .in2(N__20938),
            .in3(N__18800),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.M_this_internal_address_q_3_ns_1_8_LC_22_22_6 .C_ON=1'b0;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_8_LC_22_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.M_this_internal_address_q_3_ns_1_8_LC_22_22_6 .LUT_INIT=16'b0001101100110011;
    LogicCell40 \this_vram.M_this_internal_address_q_3_ns_1_8_LC_22_22_6  (
            .in0(N__17750),
            .in1(N__17538),
            .in2(N__18278),
            .in3(N__18797),
            .lcout(\this_vram.M_this_internal_address_q_3_ns_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_d27_2_LC_22_28_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_d27_2_LC_22_28_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_d27_2_LC_22_28_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_start_data_delay.M_this_state_d27_2_LC_22_28_5  (
            .in0(N__17513),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17501),
            .lcout(\this_start_data_delay.M_this_state_d27Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_wclke_3_LC_23_16_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_wclke_3_LC_23_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_wclke_3_LC_23_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vram.mem_mem_0_0_wclke_3_LC_23_16_0  (
            .in0(N__20759),
            .in1(N__20685),
            .in2(N__20595),
            .in3(N__20502),
            .lcout(\this_vram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_RNIU0N11_0_LC_23_17_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_0_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_0_LC_23_17_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_2_0_RNIU0N11_0_LC_23_17_3  (
            .in0(N__19619),
            .in1(N__18542),
            .in2(_gnd_net_),
            .in3(N__18527),
            .lcout(\this_vram.mem_mem_2_0_RNIU0N11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_RNI05P11_0_LC_23_18_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_RNI05P11_0_LC_23_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_RNI05P11_0_LC_23_18_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_3_0_RNI05P11_0_LC_23_18_3  (
            .in0(N__18506),
            .in1(N__18488),
            .in2(_gnd_net_),
            .in3(N__19628),
            .lcout(\this_vram.mem_mem_3_0_RNI05P11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIKREJ4_11_LC_23_18_5 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIKREJ4_11_LC_23_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIKREJ4_11_LC_23_18_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_radreg_RNIKREJ4_11_LC_23_18_5  (
            .in0(N__18351),
            .in1(N__19160),
            .in2(_gnd_net_),
            .in3(N__19277),
            .lcout(M_this_vram_read_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI95PB2_0_11_LC_23_18_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI95PB2_0_11_LC_23_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI95PB2_0_11_LC_23_18_6 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \this_vram.mem_radreg_RNI95PB2_0_11_LC_23_18_6  (
            .in0(N__19211),
            .in1(N__19097),
            .in2(N__19133),
            .in3(N__18350),
            .lcout(\this_vram.mem_DOUT_7_i_m2_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNID5PB2_11_LC_23_19_0 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNID5PB2_11_LC_23_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNID5PB2_11_LC_23_19_0 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \this_vram.mem_radreg_RNID5PB2_11_LC_23_19_0  (
            .in0(N__19199),
            .in1(N__19340),
            .in2(N__19637),
            .in3(N__18355),
            .lcout(),
            .ltout(\this_vram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNILSEJ4_11_LC_23_19_1 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNILSEJ4_11_LC_23_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNILSEJ4_11_LC_23_19_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_vram.mem_radreg_RNILSEJ4_11_LC_23_19_1  (
            .in0(N__18359),
            .in1(N__19706),
            .in2(N__18422),
            .in3(N__19739),
            .lcout(M_this_vram_read_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIDSEJ4_0_11_LC_23_19_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIDSEJ4_0_11_LC_23_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIDSEJ4_0_11_LC_23_19_7 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \this_vram.mem_radreg_RNIDSEJ4_0_11_LC_23_19_7  (
            .in0(N__19670),
            .in1(N__19526),
            .in2(N__18364),
            .in3(N__18323),
            .lcout(M_this_vram_read_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIIUD53_LC_23_21_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIIUD53_LC_23_21_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIIUD53_LC_23_21_0 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIIUD53_LC_23_21_0  (
            .in0(N__18274),
            .in1(N__20901),
            .in2(N__18219),
            .in3(N__20879),
            .lcout(M_this_vram_write_data_0_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un23_i_o2_LC_23_21_2 .C_ON=1'b0;
    defparam \this_start_data_delay.un23_i_o2_LC_23_21_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un23_i_o2_LC_23_21_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_start_data_delay.un23_i_o2_LC_23_21_2  (
            .in0(_gnd_net_),
            .in1(N__19054),
            .in2(_gnd_net_),
            .in3(N__19019),
            .lcout(\this_start_data_delay.N_351_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIDVQ81_LC_23_21_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIDVQ81_LC_23_21_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIDVQ81_LC_23_21_7 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \this_start_data_delay.M_last_q_RNIDVQ81_LC_23_21_7  (
            .in0(N__19055),
            .in1(N__19965),
            .in2(_gnd_net_),
            .in3(N__18799),
            .lcout(\this_start_data_delay.un1_M_this_state_q_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI9MQ11_LC_23_22_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI9MQ11_LC_23_22_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI9MQ11_LC_23_22_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI9MQ11_LC_23_22_1  (
            .in0(_gnd_net_),
            .in1(N__19031),
            .in2(_gnd_net_),
            .in3(N__18795),
            .lcout(M_this_vram_write_data_0_sqmuxa),
            .ltout(M_this_vram_write_data_0_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIGSD53_LC_23_22_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIGSD53_LC_23_22_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIGSD53_LC_23_22_2 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIGSD53_LC_23_22_2  (
            .in0(N__18979),
            .in1(N__18933),
            .in2(N__18890),
            .in3(N__20876),
            .lcout(M_this_vram_write_data_0_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIB2RF1_LC_23_22_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIB2RF1_LC_23_22_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIB2RF1_LC_23_22_4 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \this_start_data_delay.M_last_q_RNIB2RF1_LC_23_22_4  (
            .in0(N__18796),
            .in1(N__19943),
            .in2(_gnd_net_),
            .in3(N__18682),
            .lcout(M_this_vram_write_en_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_wclke_3_LC_24_16_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_wclke_3_LC_24_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_wclke_3_LC_24_16_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_vram.mem_mem_3_0_wclke_3_LC_24_16_2  (
            .in0(N__20762),
            .in1(N__20681),
            .in2(N__20597),
            .in3(N__20513),
            .lcout(\this_vram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_0_wclke_3_LC_24_16_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_wclke_3_LC_24_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_wclke_3_LC_24_16_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vram.mem_mem_1_0_wclke_3_LC_24_16_4  (
            .in0(N__20760),
            .in1(N__20680),
            .in2(N__20596),
            .in3(N__20511),
            .lcout(\this_vram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_wclke_3_LC_24_16_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_wclke_3_LC_24_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_wclke_3_LC_24_16_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vram.mem_mem_2_0_wclke_3_LC_24_16_5  (
            .in0(N__20512),
            .in1(N__20590),
            .in2(N__20687),
            .in3(N__20761),
            .lcout(\this_vram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_1_RNISOI11_LC_24_16_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_1_RNISOI11_LC_24_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_1_RNISOI11_LC_24_16_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_0_1_RNISOI11_LC_24_16_6  (
            .in0(N__19622),
            .in1(N__18602),
            .in2(_gnd_net_),
            .in3(N__18590),
            .lcout(\this_vram.mem_mem_0_1_RNISOIZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_1_RNI7JS51_LC_24_17_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_1_RNI7JS51_LC_24_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_1_RNI7JS51_LC_24_17_2 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \this_vram.mem_mem_1_1_RNI7JS51_LC_24_17_2  (
            .in0(N__19616),
            .in1(N__19331),
            .in2(N__19213),
            .in3(N__19319),
            .lcout(),
            .ltout(\this_vram.mem_DOUT_6_i_m2_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_1_RNI8NL72_LC_24_17_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_1_RNI8NL72_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_1_RNI8NL72_LC_24_17_3 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \this_vram.mem_mem_3_1_RNI8NL72_LC_24_17_3  (
            .in0(N__19304),
            .in1(N__19295),
            .in2(N__19280),
            .in3(N__19209),
            .lcout(\this_vram.mem_N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_1_RNI5FQ51_LC_24_17_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_1_RNI5FQ51_LC_24_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_1_RNI5FQ51_LC_24_17_4 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \this_vram.mem_mem_0_1_RNI5FQ51_LC_24_17_4  (
            .in0(N__19617),
            .in1(N__19271),
            .in2(N__19214),
            .in3(N__19259),
            .lcout(),
            .ltout(\this_vram.mem_DOUT_3_i_m2_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_1_RNI4FH72_LC_24_17_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_1_RNI4FH72_LC_24_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_1_RNI4FH72_LC_24_17_5 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \this_vram.mem_mem_2_1_RNI4FH72_LC_24_17_5  (
            .in0(N__19244),
            .in1(N__19229),
            .in2(N__19217),
            .in3(N__19210),
            .lcout(\this_vram.mem_N_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_RNIQOI11_LC_24_17_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_LC_24_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_RNIQOI11_LC_24_17_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_0_0_RNIQOI11_LC_24_17_7  (
            .in0(N__19154),
            .in1(N__19615),
            .in2(_gnd_net_),
            .in3(N__19139),
            .lcout(\this_vram.mem_mem_0_0_RNIQOIZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_RNIU0N11_LC_24_18_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_LC_24_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_RNIU0N11_LC_24_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_2_0_RNIU0N11_LC_24_18_0  (
            .in0(N__19620),
            .in1(N__19124),
            .in2(_gnd_net_),
            .in3(N__19112),
            .lcout(\this_vram.mem_mem_2_0_RNIU0NZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_4_0_wclke_3_LC_24_18_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_4_0_wclke_3_LC_24_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_4_0_wclke_3_LC_24_18_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_vram.mem_mem_4_0_wclke_3_LC_24_18_4  (
            .in0(N__20679),
            .in1(N__20751),
            .in2(N__20594),
            .in3(N__20510),
            .lcout(\this_vram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_18_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_18_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_18_5  (
            .in0(N__19070),
            .in1(N__19784),
            .in2(_gnd_net_),
            .in3(N__19621),
            .lcout(\this_vram.mem_mem_1_0_RNISSK11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_1_RNIUSK11_LC_24_19_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_1_RNIUSK11_LC_24_19_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_1_1_RNIUSK11_LC_24_19_1  (
            .in0(N__19626),
            .in1(N__19766),
            .in2(_gnd_net_),
            .in3(N__19754),
            .lcout(\this_vram.mem_mem_1_1_RNIUSKZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_1_RNI25P11_LC_24_19_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_1_RNI25P11_LC_24_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_1_RNI25P11_LC_24_19_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_3_1_RNI25P11_LC_24_19_3  (
            .in0(N__19627),
            .in1(N__19733),
            .in2(_gnd_net_),
            .in3(N__19718),
            .lcout(\this_vram.mem_mem_3_1_RNI25PZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_RNI05P11_LC_24_19_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_RNI05P11_LC_24_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_RNI05P11_LC_24_19_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_3_0_RNI05P11_LC_24_19_4  (
            .in0(N__19700),
            .in1(N__19685),
            .in2(_gnd_net_),
            .in3(N__19625),
            .lcout(\this_vram.mem_mem_3_0_RNI05PZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_1_RNI01N11_LC_24_19_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_1_RNI01N11_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_1_RNI01N11_LC_24_19_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \this_vram.mem_mem_2_1_RNI01N11_LC_24_19_6  (
            .in0(N__19664),
            .in1(_gnd_net_),
            .in2(N__19652),
            .in3(N__19623),
            .lcout(\this_vram.mem_mem_2_1_RNI01NZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_0_RNISSK11_LC_24_19_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_RNISSK11_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_RNISSK11_LC_24_19_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_1_0_RNISSK11_LC_24_19_7  (
            .in0(N__19624),
            .in1(N__19553),
            .in2(_gnd_net_),
            .in3(N__19544),
            .lcout(\this_vram.mem_mem_1_0_RNISSKZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIM2E53_LC_24_20_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIM2E53_LC_24_20_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIM2E53_LC_24_20_7 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIM2E53_LC_24_20_7  (
            .in0(N__19506),
            .in1(N__20878),
            .in2(N__19463),
            .in3(N__20902),
            .lcout(M_this_vram_write_data_0_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_5_0_wclke_3_LC_24_21_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_5_0_wclke_3_LC_24_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_5_0_wclke_3_LC_24_21_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_vram.mem_mem_5_0_wclke_3_LC_24_21_0  (
            .in0(N__20734),
            .in1(N__20567),
            .in2(N__20664),
            .in3(N__20489),
            .lcout(\this_vram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIK0E53_LC_24_21_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIK0E53_LC_24_21_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIK0E53_LC_24_21_3 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIK0E53_LC_24_21_3  (
            .in0(N__20970),
            .in1(N__20920),
            .in2(N__20903),
            .in3(N__20877),
            .lcout(M_this_vram_write_data_0_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_7_0_wclke_3_LC_24_22_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_7_0_wclke_3_LC_24_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_7_0_wclke_3_LC_24_22_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vram.mem_mem_7_0_wclke_3_LC_24_22_3  (
            .in0(N__20488),
            .in1(N__20554),
            .in2(N__20686),
            .in3(N__20750),
            .lcout(\this_vram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_6_0_wclke_3_LC_24_22_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_6_0_wclke_3_LC_24_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_6_0_wclke_3_LC_24_22_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_vram.mem_mem_6_0_wclke_3_LC_24_22_6  (
            .in0(N__20749),
            .in1(N__20675),
            .in2(N__20566),
            .in3(N__20487),
            .lcout(\this_vram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_24_24_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_24_24_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_24_24_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_24_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_0_LC_30_23_0.C_ON=1'b1;
    defparam M_this_external_address_q_0_LC_30_23_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_0_LC_30_23_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_0_LC_30_23_0 (
            .in0(N__21843),
            .in1(N__19888),
            .in2(N__20060),
            .in3(N__20059),
            .lcout(M_this_external_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_30_23_0_),
            .carryout(un1_M_this_external_address_q_cry_0),
            .clk(N__21648),
            .ce(),
            .sr(N__21350));
    defparam M_this_external_address_q_1_LC_30_23_1.C_ON=1'b1;
    defparam M_this_external_address_q_1_LC_30_23_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_1_LC_30_23_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_1_LC_30_23_1 (
            .in0(N__21851),
            .in1(N__19867),
            .in2(_gnd_net_),
            .in3(N__19856),
            .lcout(M_this_external_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_0),
            .carryout(un1_M_this_external_address_q_cry_1),
            .clk(N__21648),
            .ce(),
            .sr(N__21350));
    defparam M_this_external_address_q_2_LC_30_23_2.C_ON=1'b1;
    defparam M_this_external_address_q_2_LC_30_23_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_2_LC_30_23_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_2_LC_30_23_2 (
            .in0(N__21844),
            .in1(N__19837),
            .in2(_gnd_net_),
            .in3(N__19826),
            .lcout(M_this_external_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_1),
            .carryout(un1_M_this_external_address_q_cry_2),
            .clk(N__21648),
            .ce(),
            .sr(N__21350));
    defparam M_this_external_address_q_3_LC_30_23_3.C_ON=1'b1;
    defparam M_this_external_address_q_3_LC_30_23_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_3_LC_30_23_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_3_LC_30_23_3 (
            .in0(N__21852),
            .in1(N__19813),
            .in2(_gnd_net_),
            .in3(N__19802),
            .lcout(M_this_external_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_2),
            .carryout(un1_M_this_external_address_q_cry_3),
            .clk(N__21648),
            .ce(),
            .sr(N__21350));
    defparam M_this_external_address_q_4_LC_30_23_4.C_ON=1'b1;
    defparam M_this_external_address_q_4_LC_30_23_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_4_LC_30_23_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_4_LC_30_23_4 (
            .in0(N__21845),
            .in1(N__19795),
            .in2(_gnd_net_),
            .in3(N__21176),
            .lcout(M_this_external_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_3),
            .carryout(un1_M_this_external_address_q_cry_4),
            .clk(N__21648),
            .ce(),
            .sr(N__21350));
    defparam M_this_external_address_q_5_LC_30_23_5.C_ON=1'b1;
    defparam M_this_external_address_q_5_LC_30_23_5.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_5_LC_30_23_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_5_LC_30_23_5 (
            .in0(N__21853),
            .in1(N__21166),
            .in2(_gnd_net_),
            .in3(N__21155),
            .lcout(M_this_external_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_4),
            .carryout(un1_M_this_external_address_q_cry_5),
            .clk(N__21648),
            .ce(),
            .sr(N__21350));
    defparam M_this_external_address_q_6_LC_30_23_6.C_ON=1'b1;
    defparam M_this_external_address_q_6_LC_30_23_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_6_LC_30_23_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_6_LC_30_23_6 (
            .in0(N__21846),
            .in1(N__21145),
            .in2(_gnd_net_),
            .in3(N__21134),
            .lcout(M_this_external_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_5),
            .carryout(un1_M_this_external_address_q_cry_6),
            .clk(N__21648),
            .ce(),
            .sr(N__21350));
    defparam M_this_external_address_q_7_LC_30_23_7.C_ON=1'b1;
    defparam M_this_external_address_q_7_LC_30_23_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_7_LC_30_23_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_7_LC_30_23_7 (
            .in0(N__21854),
            .in1(N__21118),
            .in2(_gnd_net_),
            .in3(N__21107),
            .lcout(M_this_external_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_6),
            .carryout(un1_M_this_external_address_q_cry_7),
            .clk(N__21648),
            .ce(),
            .sr(N__21350));
    defparam M_this_external_address_q_8_LC_30_24_0.C_ON=1'b1;
    defparam M_this_external_address_q_8_LC_30_24_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_8_LC_30_24_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_8_LC_30_24_0 (
            .in0(N__21850),
            .in1(N__21085),
            .in2(_gnd_net_),
            .in3(N__21074),
            .lcout(M_this_external_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_30_24_0_),
            .carryout(un1_M_this_external_address_q_cry_8),
            .clk(N__21651),
            .ce(),
            .sr(N__21348));
    defparam M_this_external_address_q_9_LC_30_24_1.C_ON=1'b1;
    defparam M_this_external_address_q_9_LC_30_24_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_9_LC_30_24_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_9_LC_30_24_1 (
            .in0(N__21841),
            .in1(N__21064),
            .in2(_gnd_net_),
            .in3(N__21053),
            .lcout(M_this_external_address_qZ0Z_9),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_8),
            .carryout(un1_M_this_external_address_q_cry_9),
            .clk(N__21651),
            .ce(),
            .sr(N__21348));
    defparam M_this_external_address_q_10_LC_30_24_2.C_ON=1'b1;
    defparam M_this_external_address_q_10_LC_30_24_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_10_LC_30_24_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_10_LC_30_24_2 (
            .in0(N__21847),
            .in1(N__21034),
            .in2(_gnd_net_),
            .in3(N__21023),
            .lcout(M_this_external_address_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_9),
            .carryout(un1_M_this_external_address_q_cry_10),
            .clk(N__21651),
            .ce(),
            .sr(N__21348));
    defparam M_this_external_address_q_11_LC_30_24_3.C_ON=1'b1;
    defparam M_this_external_address_q_11_LC_30_24_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_11_LC_30_24_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_11_LC_30_24_3 (
            .in0(N__21839),
            .in1(N__21016),
            .in2(_gnd_net_),
            .in3(N__21005),
            .lcout(M_this_external_address_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_10),
            .carryout(un1_M_this_external_address_q_cry_11),
            .clk(N__21651),
            .ce(),
            .sr(N__21348));
    defparam M_this_external_address_q_12_LC_30_24_4.C_ON=1'b1;
    defparam M_this_external_address_q_12_LC_30_24_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_12_LC_30_24_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_12_LC_30_24_4 (
            .in0(N__21848),
            .in1(N__20998),
            .in2(_gnd_net_),
            .in3(N__20987),
            .lcout(M_this_external_address_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_11),
            .carryout(un1_M_this_external_address_q_cry_12),
            .clk(N__21651),
            .ce(),
            .sr(N__21348));
    defparam M_this_external_address_q_13_LC_30_24_5.C_ON=1'b1;
    defparam M_this_external_address_q_13_LC_30_24_5.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_13_LC_30_24_5.LUT_INIT=16'b1011101111101110;
    LogicCell40 M_this_external_address_q_13_LC_30_24_5 (
            .in0(N__21840),
            .in1(N__21898),
            .in2(_gnd_net_),
            .in3(N__21887),
            .lcout(M_this_external_address_qZ0Z_13),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_12),
            .carryout(un1_M_this_external_address_q_cry_13),
            .clk(N__21651),
            .ce(),
            .sr(N__21348));
    defparam M_this_external_address_q_14_LC_30_24_6.C_ON=1'b1;
    defparam M_this_external_address_q_14_LC_30_24_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_14_LC_30_24_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_14_LC_30_24_6 (
            .in0(N__21849),
            .in1(N__21874),
            .in2(_gnd_net_),
            .in3(N__21863),
            .lcout(M_this_external_address_qZ0Z_14),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_13),
            .carryout(un1_M_this_external_address_q_cry_14),
            .clk(N__21651),
            .ce(),
            .sr(N__21348));
    defparam M_this_external_address_q_15_LC_30_24_7.C_ON=1'b0;
    defparam M_this_external_address_q_15_LC_30_24_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_15_LC_30_24_7.LUT_INIT=16'b1011101111101110;
    LogicCell40 M_this_external_address_q_15_LC_30_24_7 (
            .in0(N__21842),
            .in1(N__21664),
            .in2(_gnd_net_),
            .in3(N__21680),
            .lcout(M_this_external_address_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21651),
            .ce(),
            .sr(N__21348));
    defparam \this_start_data_delay.M_this_state_d27_6_LC_32_19_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_d27_6_LC_32_19_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_d27_6_LC_32_19_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.M_this_state_d27_6_LC_32_19_5  (
            .in0(N__21266),
            .in1(N__21254),
            .in2(N__21242),
            .in3(N__21218),
            .lcout(\this_start_data_delay.M_this_state_d27Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
