-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     May 8 2022 20:03:30

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : in std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : in std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    debug : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__20240\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7101\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal port_rw_c_i : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \this_vga_signals_M_hstate_q_i_1\ : std_logic;
signal port_nmib_c_i : std_logic;
signal rgb_c_2 : std_logic;
signal rgb_c_5 : std_logic;
signal \this_vga_signals_M_hstate_q_i_4\ : std_logic;
signal rgb_c_4 : std_logic;
signal rgb_c_0 : std_logic;
signal m5 : std_logic;
signal rgb_c_1 : std_logic;
signal \rgb_2_5_0__i2_mux_0\ : std_logic;
signal \rgb_2_5_0__i2_mux\ : std_logic;
signal m19 : std_logic;
signal rgb72 : std_logic;
signal rgb_c_3 : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_0\ : std_logic;
signal port_clk_c : std_logic;
signal \this_start_data_delay_this_edge_detector_M_last_q\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_0\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_1\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_2\ : std_logic;
signal m16 : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_8\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_6\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_7\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_5\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_3\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_4\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_10_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_10_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_10_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_10_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_10_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_10_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_10_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_10_cry_7\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_10_cry_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_10_cry_2_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_10_cry_1_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_10_cry_0_THRU_CO\ : std_logic;
signal \this_vga_signals.N_238_0_cascade_\ : std_logic;
signal \this_vga_signals.N_221_0_cascade_\ : std_logic;
signal \this_vga_signals.N_232_0\ : std_logic;
signal \this_vga_signals.N_237_0_cascade_\ : std_logic;
signal \this_vga_signals.M_vstate_d_0_sqmuxa\ : std_logic;
signal \this_vga_signals.N_221_0\ : std_logic;
signal \this_vga_signals.N_225_0\ : std_logic;
signal \this_vga_signals.N_225_0_cascade_\ : std_logic;
signal \this_vga_signals.N_239_0\ : std_logic;
signal \this_vga_signals.N_239_0_cascade_\ : std_logic;
signal port_nmib_c : std_logic;
signal \this_vga_signals.N_258_cascade_\ : std_logic;
signal \this_vga_signals.N_238_0\ : std_logic;
signal \this_vga_signals.M_vstate_qZ0Z_2\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_1\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_6\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_2\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_3\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_4\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_5\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_13\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_11\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_12\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_9\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_10\ : std_logic;
signal \this_vga_signals.M_vstate_q_RNI3M6M4Z0Z_0\ : std_logic;
signal \this_vga_signals.N_251_cascade_\ : std_logic;
signal \this_vga_signals.N_237_0\ : std_logic;
signal \this_vga_signals.M_vstate_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vstate_q_srsts_0_a4_0_4_cascade_\ : std_logic;
signal \this_vga_signals.M_vstate_q_srsts_0_a4_0_4\ : std_logic;
signal \this_vga_signals.N_230_0_cascade_\ : std_logic;
signal vsync_c : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.N_230_0\ : std_logic;
signal \this_vga_signals.M_vstate_q_srsts_0_o2_2_5_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.N_248_0\ : std_logic;
signal \this_vga_signals.N_248_0_cascade_\ : std_logic;
signal \this_vga_signals.M_vstate_qZ0Z_5\ : std_logic;
signal \this_vga_signals.N_252\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_vstate_q_srsts_0_o2_2_3_cascade_\ : std_logic;
signal \this_vga_signals.N_255\ : std_logic;
signal \this_vga_signals.M_vstate_q_srsts_0_o2_2_3\ : std_logic;
signal \this_vga_signals.M_vstate_qZ0Z_3\ : std_logic;
signal \this_vga_signals.N_226_0\ : std_logic;
signal \this_vga_signals.N_256\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_7\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_10\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_11\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_8\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_9\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_14\ : std_logic;
signal \this_vga_signals.N_417_cascade_\ : std_logic;
signal \this_vga_signals.N_412_cascade_\ : std_logic;
signal \this_vga_signals.N_390_0_cascade_\ : std_logic;
signal \this_vga_signals.N_390_0\ : std_logic;
signal \this_vga_signals.M_hstate_qZ0Z_2\ : std_logic;
signal \this_vga_signals.N_413_cascade_\ : std_logic;
signal \this_vga_signals.N_398_0\ : std_logic;
signal \this_vga_signals.M_hstate_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_hstate_q_srsts_0_a3_0_4\ : std_logic;
signal \this_vga_signals.N_416\ : std_logic;
signal \this_vga_signals.M_hstate_q_srsts_0_a3_0_4_cascade_\ : std_logic;
signal \this_vga_signals.M_hstate_qZ0Z_4\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_12\ : std_logic;
signal \this_vga_signals.M_hstate_d_0_sqmuxa_cascade_\ : std_logic;
signal \this_vga_signals.N_405_0\ : std_logic;
signal \this_vga_signals.M_hstate_qZ0Z_0\ : std_logic;
signal \this_vga_signals.N_405_0_cascade_\ : std_logic;
signal \this_vga_signals.N_409\ : std_logic;
signal \this_vga_signals.N_397_0\ : std_logic;
signal \this_vga_signals.M_hstate_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_hstate_q_srsts_0_o3_2_3_5_cascade_\ : std_logic;
signal \this_vga_signals.N_385_0\ : std_logic;
signal \this_vga_signals.N_385_0_cascade_\ : std_logic;
signal \this_vga_signals.N_391_0\ : std_logic;
signal \this_vga_signals.N_386_0\ : std_logic;
signal \this_vga_signals.N_386_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hstate_q_srsts_0_o3_2_1\ : std_logic;
signal \this_vga_signals.N_388_0\ : std_logic;
signal \this_vga_signals.M_hstate_q_srsts_0_o3_2_3_5\ : std_logic;
signal \this_vga_signals.N_393_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \this_vga_signals.g2_2_cascade_\ : std_logic;
signal \this_vga_signals.g1_cascade_\ : std_logic;
signal \this_vga_signals.g2_5_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_4\ : std_logic;
signal \this_vga_signals.g0_14_N_8L16_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c3_0_0_cascade_\ : std_logic;
signal this_vga_signals_un14_address_if_generate_plus_mult1_un75_sum_i_3 : std_logic;
signal \this_vga_signals.if_N_2_6_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0\ : std_logic;
signal \this_vga_signals.g0_14_N_7L14\ : std_logic;
signal \this_vga_signals.if_N_9_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals.if_m3_1_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_3_out\ : std_logic;
signal \this_vga_signals.if_i2_mux_0\ : std_logic;
signal \this_vga_signals.if_N_6_0_0_cascade_\ : std_logic;
signal this_vga_signals_un6_address_if_generate_plus_mult1_un75_sum_i_3 : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_13\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_ac0_3_2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_ac0_3_0_a1_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_ac0_3_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_ac0_3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_ac0_3_2\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_14\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_15\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_10\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_9\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_10\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_11\ : std_logic;
signal \this_vga_signals.g1_1_1\ : std_logic;
signal \this_vga_signals.g2_1_0_cascade_\ : std_logic;
signal \this_vga_signals.g2_3_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_2_4_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_2_cascade_\ : std_logic;
signal \this_vga_signals.g0_0_6_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3\ : std_logic;
signal \this_vga_signals.g0_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb2_i\ : std_logic;
signal \this_vga_signals.g0_14_N_4L6\ : std_logic;
signal \this_vga_signals.g1_2_1\ : std_logic;
signal \this_vga_signals.g2_5_0\ : std_logic;
signal \this_vga_signals.M_vaddress_q_RNI85LKP4Z0Z_2\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_1_1_0_cascade_\ : std_logic;
signal \this_vga_signals.g3_0_0_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g1_2\ : std_logic;
signal \this_vga_signals.g2\ : std_logic;
signal \this_vga_signals.g1_0_1_0_0\ : std_logic;
signal \this_vga_signals.N_4_i\ : std_logic;
signal \this_vga_signals.g0_14_N_7L14_1\ : std_logic;
signal \this_vga_signals.if_m2_0_1\ : std_logic;
signal \this_vga_signals.if_N_3_0_i\ : std_logic;
signal \this_vga_signals.if_N_3_0_i_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c3_0\ : std_logic;
signal \this_vga_signals.if_i1_mux_0\ : std_logic;
signal \this_vga_signals.if_m2\ : std_logic;
signal \this_vga_signals.M_haddress_q_RNILVKM8Z0Z_6_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.if_N_8_i\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_3_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_1_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_4_i\ : std_logic;
signal \this_vga_signals_un6_address_if_N_5_mux_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.if_m1_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m1_9_1\ : std_logic;
signal \this_vga_signals.M_hstate_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_haddress_qZ0Z_0\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \this_vga_signals.M_haddress_qZ0Z_1\ : std_logic;
signal \this_vga_signals.un1_M_haddress_q_cry_0\ : std_logic;
signal \this_vga_signals.M_haddress_qZ0Z_2\ : std_logic;
signal \this_vga_signals.un1_M_haddress_q_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_haddress_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_haddress_q_cry_3\ : std_logic;
signal \this_vga_signals.M_haddress_qZ0Z_5\ : std_logic;
signal \this_vga_signals.un1_M_haddress_q_cry_4\ : std_logic;
signal \this_vga_signals.M_haddress_qZ0Z_6\ : std_logic;
signal \this_vga_signals.un1_M_haddress_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_haddress_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_haddress_q_cry_7\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \this_vga_signals.un1_M_haddress_q_cry_8\ : std_logic;
signal \this_vga_signals.un1_M_haddress_q_cry_9\ : std_logic;
signal \this_vga_signals.un1_M_haddress_q_cry_10\ : std_logic;
signal \this_vga_signals.M_hstate_q_RNIFIH84Z0Z_5\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_16\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_17\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_0_i\ : std_logic;
signal this_vga_signals_un6_address_if_generate_plus_mult1_un54_sum_i_3 : std_logic;
signal \this_vga_signals.g1_3_1_cascade_\ : std_logic;
signal \this_vga_signals.if_N_7_cascade_\ : std_logic;
signal \this_vga_signals.if_m1_3\ : std_logic;
signal \this_vga_signals.if_m1_3_cascade_\ : std_logic;
signal \this_vga_signals.if_m8_am_cascade_\ : std_logic;
signal \this_vga_signals.if_m8_bm\ : std_logic;
signal \this_vga_signals.g1_0_0\ : std_logic;
signal \this_vga_signals.g0_0_2_cascade_\ : std_logic;
signal \this_vga_signals.g0_0_3_0\ : std_logic;
signal \this_vga_signals.g3_2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_0_0_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_2\ : std_logic;
signal \this_vga_signals.g1_N_2L1\ : std_logic;
signal \this_vga_signals.G_5_0_x2_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals.g2_4_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_1\ : std_logic;
signal \this_vga_signals.g0_0_0_2\ : std_logic;
signal \this_vga_signals.g0_29_1\ : std_logic;
signal \this_vga_signals.N_3_0_0_0\ : std_logic;
signal \this_vga_signals.if_N_7\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_2\ : std_logic;
signal \this_vga_signals_un6_address_if_N_5_mux_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3\ : std_logic;
signal this_vga_signals_un6_address_if_generate_plus_mult1_un47_sum_i_3 : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_1\ : std_logic;
signal \this_vga_signals.CO1_1_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axb1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axbxc2_0\ : std_logic;
signal \this_vga_signals.N_2_1_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axbxc3_a4_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum1_0_3\ : std_logic;
signal \this_vga_signals.M_haddress_qZ0Z_7\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axbxc3_a5\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_ac0_2\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_15\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_18\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_16\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_17\ : std_logic;
signal \M_state_qZ0Z_5\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_252_0\ : std_logic;
signal \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_o3_0_0\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_252_0_cascade_\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_18\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_267_cascade_\ : std_logic;
signal \this_vga_signals.if_m12_bm\ : std_logic;
signal \this_vga_signals.if_m12_am\ : std_logic;
signal \this_vga_signals.if_m13_ns_1\ : std_logic;
signal if_m13_ns : std_logic;
signal \this_vga_signals.N_9_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_4_2\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_0_0_1_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_d_cascade_\ : std_logic;
signal \this_vga_signals.if_N_2_1_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_2_cascade_\ : std_logic;
signal \this_vga_signals.N_3_1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_1_x\ : std_logic;
signal \this_vga_signals.g0_3_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_2_5\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_2\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_0_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_0\ : std_logic;
signal \this_vga_signals.g0_0_5_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_3_1\ : std_logic;
signal \this_vga_signals.if_N_2_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_1_0_0\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_253_0\ : std_logic;
signal \this_vga_signals.M_haddress_qZ0Z_3\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_261_cascade_\ : std_logic;
signal \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_0Z0Z_0\ : std_logic;
signal \M_this_start_address_delay_out_0\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_267\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_275_cascade_\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_263_cascade_\ : std_logic;
signal \M_state_qZ0Z_0\ : std_logic;
signal port_address_c_0 : std_logic;
signal port_address_c_1 : std_logic;
signal \this_start_data_delay.this_edge_detector.N_275\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_259_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_i_1_3\ : std_logic;
signal \this_vga_signals.M_haddress_qZ0Z_4\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0_2\ : std_logic;
signal this_vga_signals_un6_address_if_generate_plus_mult1_un68_sum_i_3 : std_logic;
signal \this_vga_signals.g0_14_N_8L16_sx\ : std_logic;
signal \this_vga_signals.mult1_un40_sum1_3_cascade_\ : std_logic;
signal \this_vga_signals.g0_4_0\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \this_vga_signals.g0_1_1_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_1_1\ : std_logic;
signal \this_vga_signals.N_2_1_0\ : std_logic;
signal \this_vga_signals.g0_3_2_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_am_x_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_ns_2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axbxc3_5_3\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_x1_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_ns_3_cascade_\ : std_logic;
signal \this_vga_signals.N_6_i\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_am_2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum1_3\ : std_logic;
signal \this_vga_signals.N_6_i_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0\ : std_logic;
signal \this_vga_signals.if_m5_0_s\ : std_logic;
signal \this_vga_signals.if_m1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_2_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_1_0\ : std_logic;
signal \M_state_qZ0Z_2\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_d\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_0_0\ : std_logic;
signal this_vga_signals_un14_address_if_generate_plus_mult1_un54_sum_i_3 : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axbxc3_5_4\ : std_logic;
signal \this_vga_signals.M_vaddress_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_axb1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_1_1\ : std_logic;
signal \this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_0_1\ : std_logic;
signal \this_vga_signals.M_vaddress_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axbxc3_5_2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axbxc3_5_2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_1_axbxc3_a4_1_0\ : std_logic;
signal \this_vga_signals.M_vaddress_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.M_vaddress_q_fastZ0Z_9\ : std_logic;
signal \this_vga_signals.M_vaddress_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8\ : std_logic;
signal \this_vga_signals.N_353_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_bm_2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_axbxc3_5_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_axbxc3_5_3\ : std_logic;
signal \this_vga_signals.mult1_un40_sum0_3\ : std_logic;
signal \this_vga_signals.M_vaddress_q_5_repZ0Z1\ : std_logic;
signal \this_vga_signals.N_9_0\ : std_logic;
signal \this_vga_signals.M_vaddress_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vaddress_q_7_repZ0Z1\ : std_logic;
signal \this_vga_signals.N_15_0\ : std_logic;
signal \this_vga_signals.N_15_0_0_cascade_\ : std_logic;
signal \this_vga_signals.M_haddress_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_haddress_qZ0Z_8\ : std_logic;
signal \this_vga_signals.M_haddress_qZ0Z_10\ : std_logic;
signal \this_vga_signals.CO0_0\ : std_logic;
signal \M_haddress_q_RNI8ARU_11\ : std_logic;
signal \M_state_qZ0Z_1\ : std_logic;
signal port_enb_c : std_logic;
signal \M_state_qZ0Z_3\ : std_logic;
signal \M_this_start_data_delay_out_0\ : std_logic;
signal \this_vram.mem_WE_2\ : std_logic;
signal port_address_c_5 : std_logic;
signal port_address_c_2 : std_logic;
signal port_address_c_6 : std_logic;
signal \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_3Z0Z_0\ : std_logic;
signal \M_current_data_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_hstate_d_0_sqmuxa\ : std_logic;
signal \this_vga_signals.M_vaddress_qZ0Z_0\ : std_logic;
signal \bfn_23_9_0_\ : std_logic;
signal \this_vga_signals.M_vaddress_qZ0Z_1\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_0\ : std_logic;
signal \this_vga_signals.M_vaddress_qZ0Z_2\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNEZ0\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_6_c_RNISQOEZ0\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_7\ : std_logic;
signal \bfn_23_10_0_\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_8\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01REZ0\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPEZ0\ : std_logic;
signal \this_vga_signals.M_vaddress_qZ0Z_3\ : std_logic;
signal \this_vga_signals.N_1253_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_cascade_\ : std_logic;
signal \this_vga_signals.N_15_0_0\ : std_logic;
signal \this_vga_signals.N_353_0\ : std_logic;
signal \this_vga_signals.N_3520_0_cascade_\ : std_logic;
signal \this_vga_signals.CO1_2_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_2\ : std_logic;
signal \this_vga_signals.g0_1_N_2L1\ : std_logic;
signal \this_vga_signals.N_1253_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_0_2_cascade_\ : std_logic;
signal \this_vga_signals.N_3_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_0_0\ : std_logic;
signal \this_vga_signals.g0_1_N_5L7_x0_cascade_\ : std_logic;
signal \this_vga_signals.g0_1_N_5L7_x1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_m_ns_3\ : std_logic;
signal \this_vga_signals.M_vaddress_qZ0Z_4\ : std_logic;
signal \this_vga_signals.g0_1_N_5L7_ns_cascade_\ : std_logic;
signal \this_vga_signals.g0_1_1_0\ : std_logic;
signal \this_vga_signals.N_355_0\ : std_logic;
signal \this_vga_signals.g1_4\ : std_logic;
signal \this_vga_signals.M_vaddress_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_vaddress_qZ0Z_8\ : std_logic;
signal \this_vga_signals.M_vaddress_qZ0Z_6\ : std_logic;
signal \this_vga_signals.CO0\ : std_logic;
signal \this_vga_signals.if_i2_mux\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \this_vram.mem_WE_6\ : std_logic;
signal \M_current_address_qZ1Z_0\ : std_logic;
signal \M_current_address_qZ0Z_0\ : std_logic;
signal \this_vram.mem_out_bus5_0\ : std_logic;
signal \this_vram.mem_out_bus1_0\ : std_logic;
signal \this_vram.mem_mem_1_0_RNISSKZ0Z11\ : std_logic;
signal \this_vram.mem_radregZ0Z_11\ : std_logic;
signal \this_vram.mem_N_109_cascade_\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \this_vram.mem_out_bus0_0\ : std_logic;
signal \this_vram.mem_out_bus4_0\ : std_logic;
signal \this_vram.mem_mem_0_0_RNIQOIZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_N_112\ : std_logic;
signal \this_vram.mem_out_bus2_0\ : std_logic;
signal \this_vram.mem_out_bus6_0\ : std_logic;
signal \this_vram.mem_mem_2_0_RNIU0NZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus1_1\ : std_logic;
signal \this_vram.mem_out_bus5_1\ : std_logic;
signal \this_vram.mem_mem_1_0_RNISSK11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_N_88\ : std_logic;
signal \this_vram.mem_out_bus4_2\ : std_logic;
signal \this_vram.mem_out_bus0_2\ : std_logic;
signal \this_vram.mem_out_bus6_2\ : std_logic;
signal \this_vram.mem_out_bus2_2\ : std_logic;
signal \this_vram.mem_mem_0_1_RNISOIZ0Z11\ : std_logic;
signal \this_vram.mem_mem_2_1_RNI01NZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_N_98\ : std_logic;
signal \this_vram.mem_out_bus6_1\ : std_logic;
signal \this_vram.mem_out_bus2_1\ : std_logic;
signal \this_vram.mem_out_bus4_1\ : std_logic;
signal \this_vram.mem_out_bus0_1\ : std_logic;
signal \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0\ : std_logic;
signal \this_vram.mem_N_91\ : std_logic;
signal \this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKMEZ0\ : std_logic;
signal \this_vga_signals.M_vaddress_qZ0Z_5\ : std_logic;
signal \this_vga_signals.N_583_g\ : std_logic;
signal \this_vram.mem_out_bus6_3\ : std_logic;
signal \this_vram.mem_out_bus2_3\ : std_logic;
signal \this_vram.mem_mem_2_1_RNI01N11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_N_105\ : std_logic;
signal \this_vram.mem_out_bus0_3\ : std_logic;
signal \this_vram.mem_out_bus4_3\ : std_logic;
signal \this_vram.mem_mem_0_1_RNISOI11Z0Z_0\ : std_logic;
signal \this_vram.mem_WE_12\ : std_logic;
signal \this_vram.mem_out_bus7_1\ : std_logic;
signal \this_vram.mem_out_bus3_1\ : std_logic;
signal \this_vram.mem_mem_3_0_RNI05P11Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus5_3\ : std_logic;
signal \this_vram.mem_out_bus1_3\ : std_logic;
signal \this_vram.mem_mem_1_1_RNIUSK11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_N_102\ : std_logic;
signal \this_vram.mem_out_bus1_2\ : std_logic;
signal \this_vram.mem_out_bus5_2\ : std_logic;
signal \this_vram.mem_radregZ0Z_12\ : std_logic;
signal \this_vram.mem_mem_1_1_RNIUSKZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_N_95\ : std_logic;
signal \this_vram.mem_out_bus3_0\ : std_logic;
signal \this_vram.mem_out_bus7_0\ : std_logic;
signal \this_vram.mem_mem_3_0_RNI05PZ0Z11\ : std_logic;
signal \this_vram.mem_WE_10\ : std_logic;
signal \this_vram.mem_WE_8\ : std_logic;
signal \this_vram.mem_WE_14\ : std_logic;
signal \this_vram.mem_out_bus7_3\ : std_logic;
signal \this_vram.mem_out_bus3_3\ : std_logic;
signal \this_vram.mem_mem_3_1_RNI25P11Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus3_2\ : std_logic;
signal \this_vram.mem_out_bus7_2\ : std_logic;
signal \this_vram.mem_radregZ0Z_13\ : std_logic;
signal \this_vram.mem_mem_3_1_RNI25PZ0Z11\ : std_logic;
signal port_data_c_6 : std_logic;
signal \M_current_address_qZ0Z_6\ : std_logic;
signal \this_vram.mem_WE_4\ : std_logic;
signal \M_current_address_qZ0Z_12\ : std_logic;
signal \M_current_address_qZ0Z_13\ : std_logic;
signal debug_c : std_logic;
signal \this_vram.mem_WE_0\ : std_logic;
signal port_data_c_5 : std_logic;
signal \M_current_address_qZ0Z_5\ : std_logic;
signal \M_current_address_qZ0Z_11\ : std_logic;
signal port_data_c_4 : std_logic;
signal \M_current_address_qZ0Z_4\ : std_logic;
signal \M_current_address_qZ0Z_2\ : std_logic;
signal \M_current_address_qZ0Z_9\ : std_logic;
signal \M_current_data_qZ0Z_0\ : std_logic;
signal \M_current_address_qZ0Z_1\ : std_logic;
signal \M_current_address_qZ0Z_3\ : std_logic;
signal \M_current_address_q_0_0\ : std_logic;
signal \M_current_address_qZ0Z_10\ : std_logic;
signal port_data_c_0 : std_logic;
signal \M_current_address_qZ0Z_7\ : std_logic;
signal port_data_c_1 : std_logic;
signal \M_current_address_qZ0Z_8\ : std_logic;
signal \M_current_address_q_0_6_0\ : std_logic;
signal \N_631_g\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_0\ : std_logic;
signal this_vga_signals_un14_address_if_generate_plus_mult1_un61_sum_i_3 : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_i\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3\ : std_logic;
signal this_vga_signals_un6_address_if_generate_plus_mult1_un61_sum_i_3 : std_logic;
signal port_data_c_2 : std_logic;
signal \M_current_data_qZ0Z_2\ : std_logic;
signal \M_current_data_d_0_sqmuxa\ : std_logic;
signal port_data_c_3 : std_logic;
signal \M_this_reset_cond_out_0\ : std_logic;
signal \M_current_data_qZ0Z_3\ : std_logic;
signal clk_c_g : std_logic;
signal port_address_c_4 : std_logic;
signal port_address_c_7 : std_logic;
signal port_address_c_3 : std_logic;
signal port_rw_c : std_logic;
signal \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_4Z0Z_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic;
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal port_address_wire : std_logic_vector(15 downto 0);
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal port_rw_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    port_address_wire <= port_address;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    port_rw_wire <= port_rw;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \this_vram.mem_out_bus0_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus0_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= \N__12194\&\N__17591\&\N__11120\&\N__9092\&\N__13331\&\N__10685\&\N__10502\&\N__10151\&\N__19829\&\N__11618\&\N__9221\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= \N__18278\&\N__18722\&\N__17987\&\N__18137\&\N__17474\&\N__17084\&\N__16889\&\N__18431\&\N__18830\&\N__18536\&\N__15770\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14210\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18614\&'0'&'0'&'0';
    \this_vram.mem_out_bus0_3\ <= \this_vram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus0_2\ <= \this_vram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_0_1_physical_RADDR_wire\ <= \N__12188\&\N__17585\&\N__11114\&\N__9086\&\N__13325\&\N__10679\&\N__10496\&\N__10145\&\N__19823\&\N__11612\&\N__9215\;
    \this_vram.mem_mem_0_1_physical_WADDR_wire\ <= \N__18272\&\N__18716\&\N__17981\&\N__18131\&\N__17468\&\N__17078\&\N__16883\&\N__18425\&\N__18824\&\N__18530\&\N__15764\;
    \this_vram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19280\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19697\&'0'&'0'&'0';
    \this_vram.mem_out_bus1_1\ <= \this_vram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus1_0\ <= \this_vram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_1_0_physical_RADDR_wire\ <= \N__12182\&\N__17579\&\N__11108\&\N__9080\&\N__13319\&\N__10673\&\N__10490\&\N__10139\&\N__19817\&\N__11606\&\N__9209\;
    \this_vram.mem_mem_1_0_physical_WADDR_wire\ <= \N__18266\&\N__18710\&\N__17975\&\N__18125\&\N__17462\&\N__17072\&\N__16877\&\N__18419\&\N__18818\&\N__18524\&\N__15758\;
    \this_vram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14206\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18610\&'0'&'0'&'0';
    \this_vram.mem_out_bus1_3\ <= \this_vram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus1_2\ <= \this_vram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_1_1_physical_RADDR_wire\ <= \N__12176\&\N__17573\&\N__11102\&\N__9074\&\N__13313\&\N__10667\&\N__10484\&\N__10133\&\N__19811\&\N__11600\&\N__9203\;
    \this_vram.mem_mem_1_1_physical_WADDR_wire\ <= \N__18260\&\N__18704\&\N__17969\&\N__18119\&\N__17456\&\N__17066\&\N__16871\&\N__18413\&\N__18812\&\N__18518\&\N__15752\;
    \this_vram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19276\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19693\&'0'&'0'&'0';
    \this_vram.mem_out_bus2_1\ <= \this_vram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus2_0\ <= \this_vram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_2_0_physical_RADDR_wire\ <= \N__12170\&\N__17567\&\N__11096\&\N__9068\&\N__13307\&\N__10661\&\N__10478\&\N__10127\&\N__19805\&\N__11594\&\N__9197\;
    \this_vram.mem_mem_2_0_physical_WADDR_wire\ <= \N__18254\&\N__18698\&\N__17963\&\N__18113\&\N__17450\&\N__17060\&\N__16865\&\N__18407\&\N__18806\&\N__18512\&\N__15746\;
    \this_vram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14199\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18603\&'0'&'0'&'0';
    \this_vram.mem_out_bus2_3\ <= \this_vram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus2_2\ <= \this_vram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_2_1_physical_RADDR_wire\ <= \N__12164\&\N__17561\&\N__11090\&\N__9062\&\N__13301\&\N__10655\&\N__10472\&\N__10121\&\N__19799\&\N__11588\&\N__9191\;
    \this_vram.mem_mem_2_1_physical_WADDR_wire\ <= \N__18248\&\N__18692\&\N__17957\&\N__18107\&\N__17444\&\N__17054\&\N__16859\&\N__18401\&\N__18800\&\N__18506\&\N__15740\;
    \this_vram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19269\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19686\&'0'&'0'&'0';
    \this_vram.mem_out_bus3_1\ <= \this_vram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus3_0\ <= \this_vram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_3_0_physical_RADDR_wire\ <= \N__12158\&\N__17555\&\N__11084\&\N__9056\&\N__13295\&\N__10649\&\N__10466\&\N__10115\&\N__19793\&\N__11582\&\N__9185\;
    \this_vram.mem_mem_3_0_physical_WADDR_wire\ <= \N__18242\&\N__18686\&\N__17951\&\N__18101\&\N__17438\&\N__17048\&\N__16853\&\N__18395\&\N__18794\&\N__18500\&\N__15734\;
    \this_vram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14189\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18594\&'0'&'0'&'0';
    \this_vram.mem_out_bus3_3\ <= \this_vram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus3_2\ <= \this_vram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_3_1_physical_RADDR_wire\ <= \N__12152\&\N__17549\&\N__11078\&\N__9050\&\N__13289\&\N__10643\&\N__10460\&\N__10109\&\N__19787\&\N__11576\&\N__9179\;
    \this_vram.mem_mem_3_1_physical_WADDR_wire\ <= \N__18236\&\N__18680\&\N__17945\&\N__18095\&\N__17432\&\N__17042\&\N__16847\&\N__18389\&\N__18788\&\N__18494\&\N__15728\;
    \this_vram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19260\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19676\&'0'&'0'&'0';
    \this_vram.mem_out_bus4_1\ <= \this_vram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus4_0\ <= \this_vram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_4_0_physical_RADDR_wire\ <= \N__12146\&\N__17543\&\N__11072\&\N__9044\&\N__13283\&\N__10637\&\N__10454\&\N__10103\&\N__19781\&\N__11570\&\N__9173\;
    \this_vram.mem_mem_4_0_physical_WADDR_wire\ <= \N__18230\&\N__18674\&\N__17939\&\N__18089\&\N__17426\&\N__17036\&\N__16841\&\N__18383\&\N__18782\&\N__18488\&\N__15722\;
    \this_vram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14177\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18585\&'0'&'0'&'0';
    \this_vram.mem_out_bus4_3\ <= \this_vram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus4_2\ <= \this_vram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_4_1_physical_RADDR_wire\ <= \N__12140\&\N__17537\&\N__11066\&\N__9038\&\N__13277\&\N__10631\&\N__10448\&\N__10097\&\N__19775\&\N__11564\&\N__9167\;
    \this_vram.mem_mem_4_1_physical_WADDR_wire\ <= \N__18224\&\N__18668\&\N__17933\&\N__18083\&\N__17420\&\N__17030\&\N__16835\&\N__18377\&\N__18776\&\N__18482\&\N__15716\;
    \this_vram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19251\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19675\&'0'&'0'&'0';
    \this_vram.mem_out_bus5_1\ <= \this_vram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus5_0\ <= \this_vram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_5_0_physical_RADDR_wire\ <= \N__12134\&\N__17531\&\N__11060\&\N__9032\&\N__13271\&\N__10625\&\N__10442\&\N__10091\&\N__19769\&\N__11558\&\N__9161\;
    \this_vram.mem_mem_5_0_physical_WADDR_wire\ <= \N__18218\&\N__18662\&\N__17927\&\N__18077\&\N__17414\&\N__17024\&\N__16829\&\N__18371\&\N__18770\&\N__18476\&\N__15710\;
    \this_vram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14165\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18576\&'0'&'0'&'0';
    \this_vram.mem_out_bus5_3\ <= \this_vram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus5_2\ <= \this_vram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_5_1_physical_RADDR_wire\ <= \N__12128\&\N__17525\&\N__11054\&\N__9026\&\N__13265\&\N__10619\&\N__10436\&\N__10085\&\N__19763\&\N__11552\&\N__9155\;
    \this_vram.mem_mem_5_1_physical_WADDR_wire\ <= \N__18212\&\N__18656\&\N__17921\&\N__18071\&\N__17408\&\N__17018\&\N__16823\&\N__18365\&\N__18764\&\N__18470\&\N__15704\;
    \this_vram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19241\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19640\&'0'&'0'&'0';
    \this_vram.mem_out_bus6_1\ <= \this_vram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus6_0\ <= \this_vram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_6_0_physical_RADDR_wire\ <= \N__12122\&\N__17519\&\N__11048\&\N__9020\&\N__13259\&\N__10613\&\N__10430\&\N__10079\&\N__19757\&\N__11546\&\N__9149\;
    \this_vram.mem_mem_6_0_physical_WADDR_wire\ <= \N__18206\&\N__18650\&\N__17915\&\N__18065\&\N__17402\&\N__17012\&\N__16817\&\N__18359\&\N__18758\&\N__18464\&\N__15698\;
    \this_vram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14153\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18555\&'0'&'0'&'0';
    \this_vram.mem_out_bus6_3\ <= \this_vram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus6_2\ <= \this_vram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_6_1_physical_RADDR_wire\ <= \N__12116\&\N__17513\&\N__11042\&\N__9014\&\N__13253\&\N__10607\&\N__10424\&\N__10073\&\N__19751\&\N__11540\&\N__9143\;
    \this_vram.mem_mem_6_1_physical_WADDR_wire\ <= \N__18200\&\N__18644\&\N__17909\&\N__18059\&\N__17396\&\N__17006\&\N__16811\&\N__18353\&\N__18752\&\N__18458\&\N__15692\;
    \this_vram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19221\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19671\&'0'&'0'&'0';
    \this_vram.mem_out_bus7_1\ <= \this_vram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus7_0\ <= \this_vram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_7_0_physical_RADDR_wire\ <= \N__12110\&\N__17507\&\N__11036\&\N__9008\&\N__13247\&\N__10601\&\N__10418\&\N__10067\&\N__19745\&\N__11534\&\N__9137\;
    \this_vram.mem_mem_7_0_physical_WADDR_wire\ <= \N__18194\&\N__18638\&\N__17903\&\N__18053\&\N__17390\&\N__17000\&\N__16805\&\N__18347\&\N__18746\&\N__18452\&\N__15686\;
    \this_vram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__14152\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18575\&'0'&'0'&'0';
    \this_vram.mem_out_bus7_3\ <= \this_vram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus7_2\ <= \this_vram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_7_1_physical_RADDR_wire\ <= \N__12104\&\N__17501\&\N__11030\&\N__9002\&\N__13241\&\N__10595\&\N__10412\&\N__10061\&\N__19739\&\N__11528\&\N__9131\;
    \this_vram.mem_mem_7_1_physical_WADDR_wire\ <= \N__18188\&\N__18632\&\N__17897\&\N__18047\&\N__17384\&\N__16994\&\N__16799\&\N__18341\&\N__18740\&\N__18446\&\N__15680\;
    \this_vram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__19250\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19685\&'0'&'0'&'0';

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19111\,
            RE => \N__7404\,
            WCLKE => \N__16601\,
            WCLK => \N__19112\,
            WE => \N__7314\
        );

    \this_vram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19114\,
            RE => \N__7385\,
            WCLKE => \N__16597\,
            WCLK => \N__19115\,
            WE => \N__7389\
        );

    \this_vram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19119\,
            RE => \N__7384\,
            WCLKE => \N__16142\,
            WCLK => \N__19120\,
            WE => \N__7255\
        );

    \this_vram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19130\,
            RE => \N__7360\,
            WCLKE => \N__16138\,
            WCLK => \N__19131\,
            WE => \N__7421\
        );

    \this_vram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19145\,
            RE => \N__7359\,
            WCLKE => \N__16640\,
            WCLK => \N__19144\,
            WE => \N__7417\
        );

    \this_vram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19158\,
            RE => \N__7332\,
            WCLKE => \N__16636\,
            WCLK => \N__19159\,
            WE => \N__7416\
        );

    \this_vram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19166\,
            RE => \N__7331\,
            WCLKE => \N__16612\,
            WCLK => \N__19167\,
            WE => \N__7406\
        );

    \this_vram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19170\,
            RE => \N__7298\,
            WCLKE => \N__16619\,
            WCLK => \N__19171\,
            WE => \N__7405\
        );

    \this_vram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19173\,
            RE => \N__7390\,
            WCLKE => \N__15799\,
            WCLK => \N__19174\,
            WE => \N__7209\
        );

    \this_vram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19176\,
            RE => \N__7349\,
            WCLKE => \N__15800\,
            WCLK => \N__19177\,
            WE => \N__7373\
        );

    \this_vram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19180\,
            RE => \N__7350\,
            WCLKE => \N__17362\,
            WCLK => \N__19181\,
            WE => \N__7329\
        );

    \this_vram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19184\,
            RE => \N__7316\,
            WCLKE => \N__17366\,
            WCLK => \N__19185\,
            WE => \N__7320\
        );

    \this_vram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19190\,
            RE => \N__7283\,
            WCLKE => \N__14281\,
            WCLK => \N__19191\,
            WE => \N__7274\
        );

    \this_vram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19195\,
            RE => \N__7315\,
            WCLKE => \N__14285\,
            WCLK => \N__19196\,
            WE => \N__7273\
        );

    \this_vram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19199\,
            RE => \N__7218\,
            WCLKE => \N__17128\,
            WCLK => \N__19200\,
            WE => \N__7269\
        );

    \this_vram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__19201\,
            RE => \N__7282\,
            WCLKE => \N__17132\,
            WCLK => \N__19202\,
            WE => \N__7281\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__20238\,
            GLOBALBUFFEROUTPUT => clk_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20240\,
            DIN => \N__20239\,
            DOUT => \N__20238\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20240\,
            PADOUT => \N__20239\,
            PADIN => \N__20238\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20229\,
            DIN => \N__20228\,
            DOUT => \N__20227\,
            PACKAGEPIN => debug_wire
        );

    \debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20229\,
            PADOUT => \N__20228\,
            PADIN => \N__20227\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__17225\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20220\,
            DIN => \N__20219\,
            DOUT => \N__20218\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20220\,
            PADOUT => \N__20219\,
            PADIN => \N__20218\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7556\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20211\,
            DIN => \N__20210\,
            DOUT => \N__20209\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20211\,
            PADOUT => \N__20210\,
            PADIN => \N__20209\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7499\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20202\,
            DIN => \N__20201\,
            DOUT => \N__20200\,
            PACKAGEPIN => port_address_wire(0)
        );

    \port_address_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20202\,
            PADOUT => \N__20201\,
            PADIN => \N__20200\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20193\,
            DIN => \N__20192\,
            DOUT => \N__20191\,
            PACKAGEPIN => port_address_wire(1)
        );

    \port_address_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20193\,
            PADOUT => \N__20192\,
            PADIN => \N__20191\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20184\,
            DIN => \N__20183\,
            DOUT => \N__20182\,
            PACKAGEPIN => port_address_wire(2)
        );

    \port_address_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20184\,
            PADOUT => \N__20183\,
            PADIN => \N__20182\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20175\,
            DIN => \N__20174\,
            DOUT => \N__20173\,
            PACKAGEPIN => port_address_wire(3)
        );

    \port_address_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20175\,
            PADOUT => \N__20174\,
            PADIN => \N__20173\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20166\,
            DIN => \N__20165\,
            DOUT => \N__20164\,
            PACKAGEPIN => port_address_wire(4)
        );

    \port_address_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20166\,
            PADOUT => \N__20165\,
            PADIN => \N__20164\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20157\,
            DIN => \N__20156\,
            DOUT => \N__20155\,
            PACKAGEPIN => port_address_wire(5)
        );

    \port_address_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20157\,
            PADOUT => \N__20156\,
            PADIN => \N__20155\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20148\,
            DIN => \N__20147\,
            DOUT => \N__20146\,
            PACKAGEPIN => port_address_wire(6)
        );

    \port_address_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20148\,
            PADOUT => \N__20147\,
            PADIN => \N__20146\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20139\,
            DIN => \N__20138\,
            DOUT => \N__20137\,
            PACKAGEPIN => port_address_wire(7)
        );

    \port_address_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20139\,
            PADOUT => \N__20138\,
            PADIN => \N__20137\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20130\,
            DIN => \N__20129\,
            DOUT => \N__20128\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20130\,
            PADOUT => \N__20129\,
            PADIN => \N__20128\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20121\,
            DIN => \N__20120\,
            DOUT => \N__20119\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20121\,
            PADOUT => \N__20120\,
            PADIN => \N__20119\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20112\,
            DIN => \N__20111\,
            DOUT => \N__20110\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20112\,
            PADOUT => \N__20111\,
            PADIN => \N__20110\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20103\,
            DIN => \N__20102\,
            DOUT => \N__20101\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20103\,
            PADOUT => \N__20102\,
            PADIN => \N__20101\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20094\,
            DIN => \N__20093\,
            DOUT => \N__20092\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20094\,
            PADOUT => \N__20093\,
            PADIN => \N__20092\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20085\,
            DIN => \N__20084\,
            DOUT => \N__20083\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20085\,
            PADOUT => \N__20084\,
            PADIN => \N__20083\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20076\,
            DIN => \N__20075\,
            DOUT => \N__20074\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20076\,
            PADOUT => \N__20075\,
            PADIN => \N__20074\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20067\,
            DIN => \N__20066\,
            DOUT => \N__20065\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20067\,
            PADOUT => \N__20066\,
            PADIN => \N__20065\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20058\,
            DIN => \N__20057\,
            DOUT => \N__20056\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20058\,
            PADOUT => \N__20057\,
            PADIN => \N__20056\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7427\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20049\,
            DIN => \N__20048\,
            DOUT => \N__20047\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20049\,
            PADOUT => \N__20048\,
            PADIN => \N__20047\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7330\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20040\,
            DIN => \N__20039\,
            DOUT => \N__20038\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20040\,
            PADOUT => \N__20039\,
            PADIN => \N__20038\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20031\,
            DIN => \N__20030\,
            DOUT => \N__20029\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20031\,
            PADOUT => \N__20030\,
            PADIN => \N__20029\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7910\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20022\,
            DIN => \N__20021\,
            DOUT => \N__20020\,
            PACKAGEPIN => port_rw_wire
        );

    \port_rw_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20022\,
            PADOUT => \N__20021\,
            PADIN => \N__20020\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20013\,
            DIN => \N__20012\,
            DOUT => \N__20011\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20013\,
            PADOUT => \N__20012\,
            PADIN => \N__20011\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7469\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20004\,
            DIN => \N__20003\,
            DOUT => \N__20002\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20004\,
            PADOUT => \N__20003\,
            PADIN => \N__20002\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7439\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19995\,
            DIN => \N__19994\,
            DOUT => \N__19993\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__19995\,
            PADOUT => \N__19994\,
            PADIN => \N__19993\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7526\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19986\,
            DIN => \N__19985\,
            DOUT => \N__19984\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__19986\,
            PADOUT => \N__19985\,
            PADIN => \N__19984\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7580\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19977\,
            DIN => \N__19976\,
            DOUT => \N__19975\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__19977\,
            PADOUT => \N__19976\,
            PADIN => \N__19975\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7481\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19968\,
            DIN => \N__19967\,
            DOUT => \N__19966\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__19968\,
            PADOUT => \N__19967\,
            PADIN => \N__19966\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7517\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19959\,
            DIN => \N__19958\,
            DOUT => \N__19957\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__19959\,
            PADOUT => \N__19958\,
            PADIN => \N__19957\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19950\,
            DIN => \N__19949\,
            DOUT => \N__19948\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__19950\,
            PADOUT => \N__19949\,
            PADIN => \N__19948\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7538\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19941\,
            DIN => \N__19940\,
            DOUT => \N__19939\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__19941\,
            PADOUT => \N__19940\,
            PADIN => \N__19939\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8126\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__4782\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__19919\,
            I => \N__19916\
        );

    \I__4780\ : Span4Mux_v
    port map (
            O => \N__19916\,
            I => \N__19912\
        );

    \I__4779\ : InMux
    port map (
            O => \N__19915\,
            I => \N__19909\
        );

    \I__4778\ : Sp12to4
    port map (
            O => \N__19912\,
            I => \N__19905\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__19909\,
            I => \N__19901\
        );

    \I__4776\ : InMux
    port map (
            O => \N__19908\,
            I => \N__19898\
        );

    \I__4775\ : Span12Mux_v
    port map (
            O => \N__19905\,
            I => \N__19895\
        );

    \I__4774\ : InMux
    port map (
            O => \N__19904\,
            I => \N__19892\
        );

    \I__4773\ : Span4Mux_v
    port map (
            O => \N__19901\,
            I => \N__19887\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__19898\,
            I => \N__19887\
        );

    \I__4771\ : Odrv12
    port map (
            O => \N__19895\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__19892\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__4769\ : Odrv4
    port map (
            O => \N__19887\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\
        );

    \I__4768\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__4766\ : Span4Mux_s3_v
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__4765\ : Span4Mux_h
    port map (
            O => \N__19871\,
            I => \N__19868\
        );

    \I__4764\ : Span4Mux_v
    port map (
            O => \N__19868\,
            I => \N__19865\
        );

    \I__4763\ : Span4Mux_v
    port map (
            O => \N__19865\,
            I => \N__19861\
        );

    \I__4762\ : InMux
    port map (
            O => \N__19864\,
            I => \N__19858\
        );

    \I__4761\ : Span4Mux_v
    port map (
            O => \N__19861\,
            I => \N__19853\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__19858\,
            I => \N__19853\
        );

    \I__4759\ : Span4Mux_v
    port map (
            O => \N__19853\,
            I => \N__19846\
        );

    \I__4758\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19839\
        );

    \I__4757\ : InMux
    port map (
            O => \N__19851\,
            I => \N__19839\
        );

    \I__4756\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19839\
        );

    \I__4755\ : InMux
    port map (
            O => \N__19849\,
            I => \N__19836\
        );

    \I__4754\ : Odrv4
    port map (
            O => \N__19846\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__19839\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__19836\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3\
        );

    \I__4751\ : CascadeMux
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__4750\ : CascadeBuf
    port map (
            O => \N__19826\,
            I => \N__19823\
        );

    \I__4749\ : CascadeMux
    port map (
            O => \N__19823\,
            I => \N__19820\
        );

    \I__4748\ : CascadeBuf
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__19817\,
            I => \N__19814\
        );

    \I__4746\ : CascadeBuf
    port map (
            O => \N__19814\,
            I => \N__19811\
        );

    \I__4745\ : CascadeMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__4744\ : CascadeBuf
    port map (
            O => \N__19808\,
            I => \N__19805\
        );

    \I__4743\ : CascadeMux
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__4742\ : CascadeBuf
    port map (
            O => \N__19802\,
            I => \N__19799\
        );

    \I__4741\ : CascadeMux
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__4740\ : CascadeBuf
    port map (
            O => \N__19796\,
            I => \N__19793\
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__19793\,
            I => \N__19790\
        );

    \I__4738\ : CascadeBuf
    port map (
            O => \N__19790\,
            I => \N__19787\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__4736\ : CascadeBuf
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__4734\ : CascadeBuf
    port map (
            O => \N__19778\,
            I => \N__19775\
        );

    \I__4733\ : CascadeMux
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__4732\ : CascadeBuf
    port map (
            O => \N__19772\,
            I => \N__19769\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__4730\ : CascadeBuf
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__4728\ : CascadeBuf
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__4727\ : CascadeMux
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__4726\ : CascadeBuf
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__4724\ : CascadeBuf
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__4722\ : CascadeBuf
    port map (
            O => \N__19742\,
            I => \N__19739\
        );

    \I__4721\ : CascadeMux
    port map (
            O => \N__19739\,
            I => \N__19736\
        );

    \I__4720\ : InMux
    port map (
            O => \N__19736\,
            I => \N__19733\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__19733\,
            I => this_vga_signals_un6_address_if_generate_plus_mult1_un61_sum_i_3
        );

    \I__4718\ : InMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__4716\ : Span4Mux_v
    port map (
            O => \N__19724\,
            I => \N__19719\
        );

    \I__4715\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19716\
        );

    \I__4714\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19713\
        );

    \I__4713\ : Sp12to4
    port map (
            O => \N__19719\,
            I => \N__19708\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__19716\,
            I => \N__19708\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__19713\,
            I => \N__19705\
        );

    \I__4710\ : Span12Mux_h
    port map (
            O => \N__19708\,
            I => \N__19700\
        );

    \I__4709\ : Sp12to4
    port map (
            O => \N__19705\,
            I => \N__19700\
        );

    \I__4708\ : Odrv12
    port map (
            O => \N__19700\,
            I => port_data_c_2
        );

    \I__4707\ : InMux
    port map (
            O => \N__19697\,
            I => \N__19694\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__19694\,
            I => \N__19690\
        );

    \I__4705\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19687\
        );

    \I__4704\ : Span4Mux_v
    port map (
            O => \N__19690\,
            I => \N__19680\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__19687\,
            I => \N__19680\
        );

    \I__4702\ : InMux
    port map (
            O => \N__19686\,
            I => \N__19677\
        );

    \I__4701\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19672\
        );

    \I__4700\ : Span4Mux_v
    port map (
            O => \N__19680\,
            I => \N__19666\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__19677\,
            I => \N__19666\
        );

    \I__4698\ : InMux
    port map (
            O => \N__19676\,
            I => \N__19663\
        );

    \I__4697\ : InMux
    port map (
            O => \N__19675\,
            I => \N__19660\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__19672\,
            I => \N__19657\
        );

    \I__4695\ : InMux
    port map (
            O => \N__19671\,
            I => \N__19654\
        );

    \I__4694\ : Span4Mux_v
    port map (
            O => \N__19666\,
            I => \N__19649\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__19663\,
            I => \N__19649\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__19660\,
            I => \N__19646\
        );

    \I__4691\ : Span4Mux_v
    port map (
            O => \N__19657\,
            I => \N__19641\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__19654\,
            I => \N__19641\
        );

    \I__4689\ : Sp12to4
    port map (
            O => \N__19649\,
            I => \N__19636\
        );

    \I__4688\ : Span4Mux_h
    port map (
            O => \N__19646\,
            I => \N__19633\
        );

    \I__4687\ : Span4Mux_v
    port map (
            O => \N__19641\,
            I => \N__19630\
        );

    \I__4686\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19627\
        );

    \I__4685\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19624\
        );

    \I__4684\ : Odrv12
    port map (
            O => \N__19636\,
            I => \M_current_data_qZ0Z_2\
        );

    \I__4683\ : Odrv4
    port map (
            O => \N__19633\,
            I => \M_current_data_qZ0Z_2\
        );

    \I__4682\ : Odrv4
    port map (
            O => \N__19630\,
            I => \M_current_data_qZ0Z_2\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__19627\,
            I => \M_current_data_qZ0Z_2\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__19624\,
            I => \M_current_data_qZ0Z_2\
        );

    \I__4679\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19605\
        );

    \I__4677\ : InMux
    port map (
            O => \N__19609\,
            I => \N__19602\
        );

    \I__4676\ : InMux
    port map (
            O => \N__19608\,
            I => \N__19598\
        );

    \I__4675\ : Span4Mux_v
    port map (
            O => \N__19605\,
            I => \N__19593\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__19602\,
            I => \N__19593\
        );

    \I__4673\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19590\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__19598\,
            I => \N__19587\
        );

    \I__4671\ : Span4Mux_h
    port map (
            O => \N__19593\,
            I => \N__19584\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__19590\,
            I => \N__19581\
        );

    \I__4669\ : Span12Mux_s10_h
    port map (
            O => \N__19587\,
            I => \N__19574\
        );

    \I__4668\ : Sp12to4
    port map (
            O => \N__19584\,
            I => \N__19574\
        );

    \I__4667\ : Span12Mux_s5_v
    port map (
            O => \N__19581\,
            I => \N__19574\
        );

    \I__4666\ : Odrv12
    port map (
            O => \N__19574\,
            I => \M_current_data_d_0_sqmuxa\
        );

    \I__4665\ : InMux
    port map (
            O => \N__19571\,
            I => \N__19567\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__19570\,
            I => \N__19563\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__19567\,
            I => \N__19560\
        );

    \I__4662\ : InMux
    port map (
            O => \N__19566\,
            I => \N__19557\
        );

    \I__4661\ : InMux
    port map (
            O => \N__19563\,
            I => \N__19554\
        );

    \I__4660\ : Span4Mux_v
    port map (
            O => \N__19560\,
            I => \N__19551\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__19557\,
            I => \N__19546\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__19554\,
            I => \N__19546\
        );

    \I__4657\ : Span4Mux_h
    port map (
            O => \N__19551\,
            I => \N__19543\
        );

    \I__4656\ : Span12Mux_h
    port map (
            O => \N__19546\,
            I => \N__19540\
        );

    \I__4655\ : Odrv4
    port map (
            O => \N__19543\,
            I => port_data_c_3
        );

    \I__4654\ : Odrv12
    port map (
            O => \N__19540\,
            I => port_data_c_3
        );

    \I__4653\ : InMux
    port map (
            O => \N__19535\,
            I => \N__19524\
        );

    \I__4652\ : InMux
    port map (
            O => \N__19534\,
            I => \N__19524\
        );

    \I__4651\ : InMux
    port map (
            O => \N__19533\,
            I => \N__19524\
        );

    \I__4650\ : InMux
    port map (
            O => \N__19532\,
            I => \N__19520\
        );

    \I__4649\ : InMux
    port map (
            O => \N__19531\,
            I => \N__19515\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__19524\,
            I => \N__19512\
        );

    \I__4647\ : CascadeMux
    port map (
            O => \N__19523\,
            I => \N__19506\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__19520\,
            I => \N__19501\
        );

    \I__4645\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19496\
        );

    \I__4644\ : InMux
    port map (
            O => \N__19518\,
            I => \N__19496\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__19515\,
            I => \N__19491\
        );

    \I__4642\ : Span4Mux_v
    port map (
            O => \N__19512\,
            I => \N__19491\
        );

    \I__4641\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19488\
        );

    \I__4640\ : IoInMux
    port map (
            O => \N__19510\,
            I => \N__19485\
        );

    \I__4639\ : CascadeMux
    port map (
            O => \N__19509\,
            I => \N__19482\
        );

    \I__4638\ : InMux
    port map (
            O => \N__19506\,
            I => \N__19465\
        );

    \I__4637\ : InMux
    port map (
            O => \N__19505\,
            I => \N__19462\
        );

    \I__4636\ : InMux
    port map (
            O => \N__19504\,
            I => \N__19459\
        );

    \I__4635\ : Span4Mux_v
    port map (
            O => \N__19501\,
            I => \N__19456\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__19496\,
            I => \N__19449\
        );

    \I__4633\ : Span4Mux_h
    port map (
            O => \N__19491\,
            I => \N__19449\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__19488\,
            I => \N__19449\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__19485\,
            I => \N__19446\
        );

    \I__4630\ : InMux
    port map (
            O => \N__19482\,
            I => \N__19442\
        );

    \I__4629\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19439\
        );

    \I__4628\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19434\
        );

    \I__4627\ : InMux
    port map (
            O => \N__19479\,
            I => \N__19434\
        );

    \I__4626\ : InMux
    port map (
            O => \N__19478\,
            I => \N__19429\
        );

    \I__4625\ : InMux
    port map (
            O => \N__19477\,
            I => \N__19429\
        );

    \I__4624\ : InMux
    port map (
            O => \N__19476\,
            I => \N__19426\
        );

    \I__4623\ : InMux
    port map (
            O => \N__19475\,
            I => \N__19421\
        );

    \I__4622\ : InMux
    port map (
            O => \N__19474\,
            I => \N__19421\
        );

    \I__4621\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19418\
        );

    \I__4620\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19415\
        );

    \I__4619\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19412\
        );

    \I__4618\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19407\
        );

    \I__4617\ : InMux
    port map (
            O => \N__19469\,
            I => \N__19407\
        );

    \I__4616\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19404\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__19465\,
            I => \N__19401\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__19462\,
            I => \N__19398\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__19459\,
            I => \N__19395\
        );

    \I__4612\ : Span4Mux_h
    port map (
            O => \N__19456\,
            I => \N__19390\
        );

    \I__4611\ : Span4Mux_v
    port map (
            O => \N__19449\,
            I => \N__19390\
        );

    \I__4610\ : Span4Mux_s3_v
    port map (
            O => \N__19446\,
            I => \N__19387\
        );

    \I__4609\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19384\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__19442\,
            I => \N__19379\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__19439\,
            I => \N__19379\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__19434\,
            I => \N__19370\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__19429\,
            I => \N__19370\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__19426\,
            I => \N__19363\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__19421\,
            I => \N__19363\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__19418\,
            I => \N__19363\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__19415\,
            I => \N__19358\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__19412\,
            I => \N__19358\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__19407\,
            I => \N__19353\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__19404\,
            I => \N__19353\
        );

    \I__4597\ : Span4Mux_v
    port map (
            O => \N__19401\,
            I => \N__19346\
        );

    \I__4596\ : Span4Mux_v
    port map (
            O => \N__19398\,
            I => \N__19346\
        );

    \I__4595\ : Span4Mux_v
    port map (
            O => \N__19395\,
            I => \N__19346\
        );

    \I__4594\ : Span4Mux_v
    port map (
            O => \N__19390\,
            I => \N__19341\
        );

    \I__4593\ : Span4Mux_v
    port map (
            O => \N__19387\,
            I => \N__19341\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__19384\,
            I => \N__19336\
        );

    \I__4591\ : Span4Mux_v
    port map (
            O => \N__19379\,
            I => \N__19336\
        );

    \I__4590\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19327\
        );

    \I__4589\ : InMux
    port map (
            O => \N__19377\,
            I => \N__19327\
        );

    \I__4588\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19327\
        );

    \I__4587\ : InMux
    port map (
            O => \N__19375\,
            I => \N__19327\
        );

    \I__4586\ : Span4Mux_h
    port map (
            O => \N__19370\,
            I => \N__19324\
        );

    \I__4585\ : Span4Mux_h
    port map (
            O => \N__19363\,
            I => \N__19321\
        );

    \I__4584\ : Span4Mux_h
    port map (
            O => \N__19358\,
            I => \N__19316\
        );

    \I__4583\ : Span4Mux_h
    port map (
            O => \N__19353\,
            I => \N__19316\
        );

    \I__4582\ : Sp12to4
    port map (
            O => \N__19346\,
            I => \N__19311\
        );

    \I__4581\ : Sp12to4
    port map (
            O => \N__19341\,
            I => \N__19311\
        );

    \I__4580\ : Span4Mux_h
    port map (
            O => \N__19336\,
            I => \N__19308\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__19327\,
            I => \N__19303\
        );

    \I__4578\ : Span4Mux_v
    port map (
            O => \N__19324\,
            I => \N__19303\
        );

    \I__4577\ : Sp12to4
    port map (
            O => \N__19321\,
            I => \N__19296\
        );

    \I__4576\ : Sp12to4
    port map (
            O => \N__19316\,
            I => \N__19296\
        );

    \I__4575\ : Span12Mux_h
    port map (
            O => \N__19311\,
            I => \N__19296\
        );

    \I__4574\ : Span4Mux_v
    port map (
            O => \N__19308\,
            I => \N__19293\
        );

    \I__4573\ : Span4Mux_v
    port map (
            O => \N__19303\,
            I => \N__19290\
        );

    \I__4572\ : Span12Mux_v
    port map (
            O => \N__19296\,
            I => \N__19287\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__19293\,
            I => \M_this_reset_cond_out_0\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__19290\,
            I => \M_this_reset_cond_out_0\
        );

    \I__4569\ : Odrv12
    port map (
            O => \N__19287\,
            I => \M_this_reset_cond_out_0\
        );

    \I__4568\ : InMux
    port map (
            O => \N__19280\,
            I => \N__19277\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__19277\,
            I => \N__19273\
        );

    \I__4566\ : InMux
    port map (
            O => \N__19276\,
            I => \N__19270\
        );

    \I__4565\ : Span4Mux_v
    port map (
            O => \N__19273\,
            I => \N__19264\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__19270\,
            I => \N__19264\
        );

    \I__4563\ : InMux
    port map (
            O => \N__19269\,
            I => \N__19261\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__19264\,
            I => \N__19255\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__19261\,
            I => \N__19255\
        );

    \I__4560\ : InMux
    port map (
            O => \N__19260\,
            I => \N__19252\
        );

    \I__4559\ : Span4Mux_v
    port map (
            O => \N__19255\,
            I => \N__19245\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__19252\,
            I => \N__19245\
        );

    \I__4557\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19242\
        );

    \I__4556\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19238\
        );

    \I__4555\ : Span4Mux_v
    port map (
            O => \N__19245\,
            I => \N__19233\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__19242\,
            I => \N__19233\
        );

    \I__4553\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19230\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__19238\,
            I => \N__19227\
        );

    \I__4551\ : Span4Mux_v
    port map (
            O => \N__19233\,
            I => \N__19222\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__19230\,
            I => \N__19222\
        );

    \I__4549\ : Span4Mux_s2_v
    port map (
            O => \N__19227\,
            I => \N__19215\
        );

    \I__4548\ : Span4Mux_v
    port map (
            O => \N__19222\,
            I => \N__19215\
        );

    \I__4547\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19212\
        );

    \I__4546\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19209\
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__19215\,
            I => \M_current_data_qZ0Z_3\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__19212\,
            I => \M_current_data_qZ0Z_3\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__19209\,
            I => \M_current_data_qZ0Z_3\
        );

    \I__4542\ : ClkMux
    port map (
            O => \N__19202\,
            I => \N__18923\
        );

    \I__4541\ : ClkMux
    port map (
            O => \N__19201\,
            I => \N__18923\
        );

    \I__4540\ : ClkMux
    port map (
            O => \N__19200\,
            I => \N__18923\
        );

    \I__4539\ : ClkMux
    port map (
            O => \N__19199\,
            I => \N__18923\
        );

    \I__4538\ : ClkMux
    port map (
            O => \N__19198\,
            I => \N__18923\
        );

    \I__4537\ : ClkMux
    port map (
            O => \N__19197\,
            I => \N__18923\
        );

    \I__4536\ : ClkMux
    port map (
            O => \N__19196\,
            I => \N__18923\
        );

    \I__4535\ : ClkMux
    port map (
            O => \N__19195\,
            I => \N__18923\
        );

    \I__4534\ : ClkMux
    port map (
            O => \N__19194\,
            I => \N__18923\
        );

    \I__4533\ : ClkMux
    port map (
            O => \N__19193\,
            I => \N__18923\
        );

    \I__4532\ : ClkMux
    port map (
            O => \N__19192\,
            I => \N__18923\
        );

    \I__4531\ : ClkMux
    port map (
            O => \N__19191\,
            I => \N__18923\
        );

    \I__4530\ : ClkMux
    port map (
            O => \N__19190\,
            I => \N__18923\
        );

    \I__4529\ : ClkMux
    port map (
            O => \N__19189\,
            I => \N__18923\
        );

    \I__4528\ : ClkMux
    port map (
            O => \N__19188\,
            I => \N__18923\
        );

    \I__4527\ : ClkMux
    port map (
            O => \N__19187\,
            I => \N__18923\
        );

    \I__4526\ : ClkMux
    port map (
            O => \N__19186\,
            I => \N__18923\
        );

    \I__4525\ : ClkMux
    port map (
            O => \N__19185\,
            I => \N__18923\
        );

    \I__4524\ : ClkMux
    port map (
            O => \N__19184\,
            I => \N__18923\
        );

    \I__4523\ : ClkMux
    port map (
            O => \N__19183\,
            I => \N__18923\
        );

    \I__4522\ : ClkMux
    port map (
            O => \N__19182\,
            I => \N__18923\
        );

    \I__4521\ : ClkMux
    port map (
            O => \N__19181\,
            I => \N__18923\
        );

    \I__4520\ : ClkMux
    port map (
            O => \N__19180\,
            I => \N__18923\
        );

    \I__4519\ : ClkMux
    port map (
            O => \N__19179\,
            I => \N__18923\
        );

    \I__4518\ : ClkMux
    port map (
            O => \N__19178\,
            I => \N__18923\
        );

    \I__4517\ : ClkMux
    port map (
            O => \N__19177\,
            I => \N__18923\
        );

    \I__4516\ : ClkMux
    port map (
            O => \N__19176\,
            I => \N__18923\
        );

    \I__4515\ : ClkMux
    port map (
            O => \N__19175\,
            I => \N__18923\
        );

    \I__4514\ : ClkMux
    port map (
            O => \N__19174\,
            I => \N__18923\
        );

    \I__4513\ : ClkMux
    port map (
            O => \N__19173\,
            I => \N__18923\
        );

    \I__4512\ : ClkMux
    port map (
            O => \N__19172\,
            I => \N__18923\
        );

    \I__4511\ : ClkMux
    port map (
            O => \N__19171\,
            I => \N__18923\
        );

    \I__4510\ : ClkMux
    port map (
            O => \N__19170\,
            I => \N__18923\
        );

    \I__4509\ : ClkMux
    port map (
            O => \N__19169\,
            I => \N__18923\
        );

    \I__4508\ : ClkMux
    port map (
            O => \N__19168\,
            I => \N__18923\
        );

    \I__4507\ : ClkMux
    port map (
            O => \N__19167\,
            I => \N__18923\
        );

    \I__4506\ : ClkMux
    port map (
            O => \N__19166\,
            I => \N__18923\
        );

    \I__4505\ : ClkMux
    port map (
            O => \N__19165\,
            I => \N__18923\
        );

    \I__4504\ : ClkMux
    port map (
            O => \N__19164\,
            I => \N__18923\
        );

    \I__4503\ : ClkMux
    port map (
            O => \N__19163\,
            I => \N__18923\
        );

    \I__4502\ : ClkMux
    port map (
            O => \N__19162\,
            I => \N__18923\
        );

    \I__4501\ : ClkMux
    port map (
            O => \N__19161\,
            I => \N__18923\
        );

    \I__4500\ : ClkMux
    port map (
            O => \N__19160\,
            I => \N__18923\
        );

    \I__4499\ : ClkMux
    port map (
            O => \N__19159\,
            I => \N__18923\
        );

    \I__4498\ : ClkMux
    port map (
            O => \N__19158\,
            I => \N__18923\
        );

    \I__4497\ : ClkMux
    port map (
            O => \N__19157\,
            I => \N__18923\
        );

    \I__4496\ : ClkMux
    port map (
            O => \N__19156\,
            I => \N__18923\
        );

    \I__4495\ : ClkMux
    port map (
            O => \N__19155\,
            I => \N__18923\
        );

    \I__4494\ : ClkMux
    port map (
            O => \N__19154\,
            I => \N__18923\
        );

    \I__4493\ : ClkMux
    port map (
            O => \N__19153\,
            I => \N__18923\
        );

    \I__4492\ : ClkMux
    port map (
            O => \N__19152\,
            I => \N__18923\
        );

    \I__4491\ : ClkMux
    port map (
            O => \N__19151\,
            I => \N__18923\
        );

    \I__4490\ : ClkMux
    port map (
            O => \N__19150\,
            I => \N__18923\
        );

    \I__4489\ : ClkMux
    port map (
            O => \N__19149\,
            I => \N__18923\
        );

    \I__4488\ : ClkMux
    port map (
            O => \N__19148\,
            I => \N__18923\
        );

    \I__4487\ : ClkMux
    port map (
            O => \N__19147\,
            I => \N__18923\
        );

    \I__4486\ : ClkMux
    port map (
            O => \N__19146\,
            I => \N__18923\
        );

    \I__4485\ : ClkMux
    port map (
            O => \N__19145\,
            I => \N__18923\
        );

    \I__4484\ : ClkMux
    port map (
            O => \N__19144\,
            I => \N__18923\
        );

    \I__4483\ : ClkMux
    port map (
            O => \N__19143\,
            I => \N__18923\
        );

    \I__4482\ : ClkMux
    port map (
            O => \N__19142\,
            I => \N__18923\
        );

    \I__4481\ : ClkMux
    port map (
            O => \N__19141\,
            I => \N__18923\
        );

    \I__4480\ : ClkMux
    port map (
            O => \N__19140\,
            I => \N__18923\
        );

    \I__4479\ : ClkMux
    port map (
            O => \N__19139\,
            I => \N__18923\
        );

    \I__4478\ : ClkMux
    port map (
            O => \N__19138\,
            I => \N__18923\
        );

    \I__4477\ : ClkMux
    port map (
            O => \N__19137\,
            I => \N__18923\
        );

    \I__4476\ : ClkMux
    port map (
            O => \N__19136\,
            I => \N__18923\
        );

    \I__4475\ : ClkMux
    port map (
            O => \N__19135\,
            I => \N__18923\
        );

    \I__4474\ : ClkMux
    port map (
            O => \N__19134\,
            I => \N__18923\
        );

    \I__4473\ : ClkMux
    port map (
            O => \N__19133\,
            I => \N__18923\
        );

    \I__4472\ : ClkMux
    port map (
            O => \N__19132\,
            I => \N__18923\
        );

    \I__4471\ : ClkMux
    port map (
            O => \N__19131\,
            I => \N__18923\
        );

    \I__4470\ : ClkMux
    port map (
            O => \N__19130\,
            I => \N__18923\
        );

    \I__4469\ : ClkMux
    port map (
            O => \N__19129\,
            I => \N__18923\
        );

    \I__4468\ : ClkMux
    port map (
            O => \N__19128\,
            I => \N__18923\
        );

    \I__4467\ : ClkMux
    port map (
            O => \N__19127\,
            I => \N__18923\
        );

    \I__4466\ : ClkMux
    port map (
            O => \N__19126\,
            I => \N__18923\
        );

    \I__4465\ : ClkMux
    port map (
            O => \N__19125\,
            I => \N__18923\
        );

    \I__4464\ : ClkMux
    port map (
            O => \N__19124\,
            I => \N__18923\
        );

    \I__4463\ : ClkMux
    port map (
            O => \N__19123\,
            I => \N__18923\
        );

    \I__4462\ : ClkMux
    port map (
            O => \N__19122\,
            I => \N__18923\
        );

    \I__4461\ : ClkMux
    port map (
            O => \N__19121\,
            I => \N__18923\
        );

    \I__4460\ : ClkMux
    port map (
            O => \N__19120\,
            I => \N__18923\
        );

    \I__4459\ : ClkMux
    port map (
            O => \N__19119\,
            I => \N__18923\
        );

    \I__4458\ : ClkMux
    port map (
            O => \N__19118\,
            I => \N__18923\
        );

    \I__4457\ : ClkMux
    port map (
            O => \N__19117\,
            I => \N__18923\
        );

    \I__4456\ : ClkMux
    port map (
            O => \N__19116\,
            I => \N__18923\
        );

    \I__4455\ : ClkMux
    port map (
            O => \N__19115\,
            I => \N__18923\
        );

    \I__4454\ : ClkMux
    port map (
            O => \N__19114\,
            I => \N__18923\
        );

    \I__4453\ : ClkMux
    port map (
            O => \N__19113\,
            I => \N__18923\
        );

    \I__4452\ : ClkMux
    port map (
            O => \N__19112\,
            I => \N__18923\
        );

    \I__4451\ : ClkMux
    port map (
            O => \N__19111\,
            I => \N__18923\
        );

    \I__4450\ : ClkMux
    port map (
            O => \N__19110\,
            I => \N__18923\
        );

    \I__4449\ : GlobalMux
    port map (
            O => \N__18923\,
            I => \N__18920\
        );

    \I__4448\ : gio2CtrlBuf
    port map (
            O => \N__18920\,
            I => clk_c_g
        );

    \I__4447\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__4445\ : Span4Mux_v
    port map (
            O => \N__18911\,
            I => \N__18908\
        );

    \I__4444\ : Odrv4
    port map (
            O => \N__18908\,
            I => port_address_c_4
        );

    \I__4443\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__18902\,
            I => \N__18899\
        );

    \I__4441\ : Span4Mux_v
    port map (
            O => \N__18899\,
            I => \N__18896\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__4439\ : Span4Mux_v
    port map (
            O => \N__18893\,
            I => \N__18890\
        );

    \I__4438\ : Span4Mux_v
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__4437\ : Odrv4
    port map (
            O => \N__18887\,
            I => port_address_c_7
        );

    \I__4436\ : CascadeMux
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__4435\ : InMux
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__18878\,
            I => \N__18875\
        );

    \I__4433\ : Span12Mux_v
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__4432\ : Odrv12
    port map (
            O => \N__18872\,
            I => port_address_c_3
        );

    \I__4431\ : InMux
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__18866\,
            I => \N__18863\
        );

    \I__4429\ : Span12Mux_s10_h
    port map (
            O => \N__18863\,
            I => \N__18860\
        );

    \I__4428\ : Span12Mux_h
    port map (
            O => \N__18860\,
            I => \N__18856\
        );

    \I__4427\ : InMux
    port map (
            O => \N__18859\,
            I => \N__18853\
        );

    \I__4426\ : Odrv12
    port map (
            O => \N__18856\,
            I => port_rw_c
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__18853\,
            I => port_rw_c
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__18848\,
            I => \N__18845\
        );

    \I__4423\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__18842\,
            I => \N__18839\
        );

    \I__4421\ : Span12Mux_v
    port map (
            O => \N__18839\,
            I => \N__18836\
        );

    \I__4420\ : Span12Mux_h
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__4419\ : Odrv12
    port map (
            O => \N__18833\,
            I => \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_4Z0Z_0\
        );

    \I__4418\ : CascadeMux
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__4417\ : CascadeBuf
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__4416\ : CascadeMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__4415\ : CascadeBuf
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__4414\ : CascadeMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__4413\ : CascadeBuf
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__4411\ : CascadeBuf
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__4410\ : CascadeMux
    port map (
            O => \N__18806\,
            I => \N__18803\
        );

    \I__4409\ : CascadeBuf
    port map (
            O => \N__18803\,
            I => \N__18800\
        );

    \I__4408\ : CascadeMux
    port map (
            O => \N__18800\,
            I => \N__18797\
        );

    \I__4407\ : CascadeBuf
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__4406\ : CascadeMux
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__4405\ : CascadeBuf
    port map (
            O => \N__18791\,
            I => \N__18788\
        );

    \I__4404\ : CascadeMux
    port map (
            O => \N__18788\,
            I => \N__18785\
        );

    \I__4403\ : CascadeBuf
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__4402\ : CascadeMux
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__4401\ : CascadeBuf
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__4400\ : CascadeMux
    port map (
            O => \N__18776\,
            I => \N__18773\
        );

    \I__4399\ : CascadeBuf
    port map (
            O => \N__18773\,
            I => \N__18770\
        );

    \I__4398\ : CascadeMux
    port map (
            O => \N__18770\,
            I => \N__18767\
        );

    \I__4397\ : CascadeBuf
    port map (
            O => \N__18767\,
            I => \N__18764\
        );

    \I__4396\ : CascadeMux
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__4395\ : CascadeBuf
    port map (
            O => \N__18761\,
            I => \N__18758\
        );

    \I__4394\ : CascadeMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__4393\ : CascadeBuf
    port map (
            O => \N__18755\,
            I => \N__18752\
        );

    \I__4392\ : CascadeMux
    port map (
            O => \N__18752\,
            I => \N__18749\
        );

    \I__4391\ : CascadeBuf
    port map (
            O => \N__18749\,
            I => \N__18746\
        );

    \I__4390\ : CascadeMux
    port map (
            O => \N__18746\,
            I => \N__18743\
        );

    \I__4389\ : CascadeBuf
    port map (
            O => \N__18743\,
            I => \N__18740\
        );

    \I__4388\ : CascadeMux
    port map (
            O => \N__18740\,
            I => \N__18737\
        );

    \I__4387\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18734\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__18734\,
            I => \N__18731\
        );

    \I__4385\ : Span4Mux_s1_v
    port map (
            O => \N__18731\,
            I => \N__18728\
        );

    \I__4384\ : Span4Mux_v
    port map (
            O => \N__18728\,
            I => \N__18725\
        );

    \I__4383\ : Odrv4
    port map (
            O => \N__18725\,
            I => \M_current_address_qZ0Z_2\
        );

    \I__4382\ : CascadeMux
    port map (
            O => \N__18722\,
            I => \N__18719\
        );

    \I__4381\ : CascadeBuf
    port map (
            O => \N__18719\,
            I => \N__18716\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__18716\,
            I => \N__18713\
        );

    \I__4379\ : CascadeBuf
    port map (
            O => \N__18713\,
            I => \N__18710\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__18710\,
            I => \N__18707\
        );

    \I__4377\ : CascadeBuf
    port map (
            O => \N__18707\,
            I => \N__18704\
        );

    \I__4376\ : CascadeMux
    port map (
            O => \N__18704\,
            I => \N__18701\
        );

    \I__4375\ : CascadeBuf
    port map (
            O => \N__18701\,
            I => \N__18698\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__18698\,
            I => \N__18695\
        );

    \I__4373\ : CascadeBuf
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__4372\ : CascadeMux
    port map (
            O => \N__18692\,
            I => \N__18689\
        );

    \I__4371\ : CascadeBuf
    port map (
            O => \N__18689\,
            I => \N__18686\
        );

    \I__4370\ : CascadeMux
    port map (
            O => \N__18686\,
            I => \N__18683\
        );

    \I__4369\ : CascadeBuf
    port map (
            O => \N__18683\,
            I => \N__18680\
        );

    \I__4368\ : CascadeMux
    port map (
            O => \N__18680\,
            I => \N__18677\
        );

    \I__4367\ : CascadeBuf
    port map (
            O => \N__18677\,
            I => \N__18674\
        );

    \I__4366\ : CascadeMux
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__4365\ : CascadeBuf
    port map (
            O => \N__18671\,
            I => \N__18668\
        );

    \I__4364\ : CascadeMux
    port map (
            O => \N__18668\,
            I => \N__18665\
        );

    \I__4363\ : CascadeBuf
    port map (
            O => \N__18665\,
            I => \N__18662\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__18662\,
            I => \N__18659\
        );

    \I__4361\ : CascadeBuf
    port map (
            O => \N__18659\,
            I => \N__18656\
        );

    \I__4360\ : CascadeMux
    port map (
            O => \N__18656\,
            I => \N__18653\
        );

    \I__4359\ : CascadeBuf
    port map (
            O => \N__18653\,
            I => \N__18650\
        );

    \I__4358\ : CascadeMux
    port map (
            O => \N__18650\,
            I => \N__18647\
        );

    \I__4357\ : CascadeBuf
    port map (
            O => \N__18647\,
            I => \N__18644\
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__18644\,
            I => \N__18641\
        );

    \I__4355\ : CascadeBuf
    port map (
            O => \N__18641\,
            I => \N__18638\
        );

    \I__4354\ : CascadeMux
    port map (
            O => \N__18638\,
            I => \N__18635\
        );

    \I__4353\ : CascadeBuf
    port map (
            O => \N__18635\,
            I => \N__18632\
        );

    \I__4352\ : CascadeMux
    port map (
            O => \N__18632\,
            I => \N__18629\
        );

    \I__4351\ : InMux
    port map (
            O => \N__18629\,
            I => \N__18626\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__18626\,
            I => \N__18623\
        );

    \I__4349\ : Span4Mux_s1_v
    port map (
            O => \N__18623\,
            I => \N__18620\
        );

    \I__4348\ : Span4Mux_v
    port map (
            O => \N__18620\,
            I => \N__18617\
        );

    \I__4347\ : Odrv4
    port map (
            O => \N__18617\,
            I => \M_current_address_qZ0Z_9\
        );

    \I__4346\ : InMux
    port map (
            O => \N__18614\,
            I => \N__18611\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__18611\,
            I => \N__18607\
        );

    \I__4344\ : InMux
    port map (
            O => \N__18610\,
            I => \N__18604\
        );

    \I__4343\ : Span4Mux_v
    port map (
            O => \N__18607\,
            I => \N__18598\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__18604\,
            I => \N__18598\
        );

    \I__4341\ : InMux
    port map (
            O => \N__18603\,
            I => \N__18595\
        );

    \I__4340\ : Span4Mux_v
    port map (
            O => \N__18598\,
            I => \N__18589\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__18595\,
            I => \N__18589\
        );

    \I__4338\ : InMux
    port map (
            O => \N__18594\,
            I => \N__18586\
        );

    \I__4337\ : Span4Mux_v
    port map (
            O => \N__18589\,
            I => \N__18580\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__18586\,
            I => \N__18580\
        );

    \I__4335\ : InMux
    port map (
            O => \N__18585\,
            I => \N__18577\
        );

    \I__4334\ : Span4Mux_v
    port map (
            O => \N__18580\,
            I => \N__18570\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__18577\,
            I => \N__18570\
        );

    \I__4332\ : InMux
    port map (
            O => \N__18576\,
            I => \N__18567\
        );

    \I__4331\ : InMux
    port map (
            O => \N__18575\,
            I => \N__18564\
        );

    \I__4330\ : Span4Mux_v
    port map (
            O => \N__18570\,
            I => \N__18559\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__18567\,
            I => \N__18559\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__18564\,
            I => \N__18556\
        );

    \I__4327\ : Span4Mux_v
    port map (
            O => \N__18559\,
            I => \N__18549\
        );

    \I__4326\ : Span4Mux_s3_v
    port map (
            O => \N__18556\,
            I => \N__18549\
        );

    \I__4325\ : InMux
    port map (
            O => \N__18555\,
            I => \N__18546\
        );

    \I__4324\ : InMux
    port map (
            O => \N__18554\,
            I => \N__18543\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__18549\,
            I => \M_current_data_qZ0Z_0\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__18546\,
            I => \M_current_data_qZ0Z_0\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__18543\,
            I => \M_current_data_qZ0Z_0\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__18536\,
            I => \N__18533\
        );

    \I__4319\ : CascadeBuf
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__4317\ : CascadeBuf
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__4316\ : CascadeMux
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__4315\ : CascadeBuf
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__4314\ : CascadeMux
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__4313\ : CascadeBuf
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__4311\ : CascadeBuf
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__4309\ : CascadeBuf
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__4307\ : CascadeBuf
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__4306\ : CascadeMux
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__4305\ : CascadeBuf
    port map (
            O => \N__18491\,
            I => \N__18488\
        );

    \I__4304\ : CascadeMux
    port map (
            O => \N__18488\,
            I => \N__18485\
        );

    \I__4303\ : CascadeBuf
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__4301\ : CascadeBuf
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__18476\,
            I => \N__18473\
        );

    \I__4299\ : CascadeBuf
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__4298\ : CascadeMux
    port map (
            O => \N__18470\,
            I => \N__18467\
        );

    \I__4297\ : CascadeBuf
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__4296\ : CascadeMux
    port map (
            O => \N__18464\,
            I => \N__18461\
        );

    \I__4295\ : CascadeBuf
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__4294\ : CascadeMux
    port map (
            O => \N__18458\,
            I => \N__18455\
        );

    \I__4293\ : CascadeBuf
    port map (
            O => \N__18455\,
            I => \N__18452\
        );

    \I__4292\ : CascadeMux
    port map (
            O => \N__18452\,
            I => \N__18449\
        );

    \I__4291\ : CascadeBuf
    port map (
            O => \N__18449\,
            I => \N__18446\
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__18446\,
            I => \N__18443\
        );

    \I__4289\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__18440\,
            I => \N__18437\
        );

    \I__4287\ : Span4Mux_s2_v
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__4286\ : Odrv4
    port map (
            O => \N__18434\,
            I => \M_current_address_qZ0Z_1\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__18431\,
            I => \N__18428\
        );

    \I__4284\ : CascadeBuf
    port map (
            O => \N__18428\,
            I => \N__18425\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__18425\,
            I => \N__18422\
        );

    \I__4282\ : CascadeBuf
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__4281\ : CascadeMux
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__4280\ : CascadeBuf
    port map (
            O => \N__18416\,
            I => \N__18413\
        );

    \I__4279\ : CascadeMux
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__4278\ : CascadeBuf
    port map (
            O => \N__18410\,
            I => \N__18407\
        );

    \I__4277\ : CascadeMux
    port map (
            O => \N__18407\,
            I => \N__18404\
        );

    \I__4276\ : CascadeBuf
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__4275\ : CascadeMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__4274\ : CascadeBuf
    port map (
            O => \N__18398\,
            I => \N__18395\
        );

    \I__4273\ : CascadeMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__4272\ : CascadeBuf
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__4271\ : CascadeMux
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__4270\ : CascadeBuf
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__4269\ : CascadeMux
    port map (
            O => \N__18383\,
            I => \N__18380\
        );

    \I__4268\ : CascadeBuf
    port map (
            O => \N__18380\,
            I => \N__18377\
        );

    \I__4267\ : CascadeMux
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__4266\ : CascadeBuf
    port map (
            O => \N__18374\,
            I => \N__18371\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__18371\,
            I => \N__18368\
        );

    \I__4264\ : CascadeBuf
    port map (
            O => \N__18368\,
            I => \N__18365\
        );

    \I__4263\ : CascadeMux
    port map (
            O => \N__18365\,
            I => \N__18362\
        );

    \I__4262\ : CascadeBuf
    port map (
            O => \N__18362\,
            I => \N__18359\
        );

    \I__4261\ : CascadeMux
    port map (
            O => \N__18359\,
            I => \N__18356\
        );

    \I__4260\ : CascadeBuf
    port map (
            O => \N__18356\,
            I => \N__18353\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__18353\,
            I => \N__18350\
        );

    \I__4258\ : CascadeBuf
    port map (
            O => \N__18350\,
            I => \N__18347\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__18347\,
            I => \N__18344\
        );

    \I__4256\ : CascadeBuf
    port map (
            O => \N__18344\,
            I => \N__18341\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__18341\,
            I => \N__18338\
        );

    \I__4254\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18335\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__4252\ : Span4Mux_s3_v
    port map (
            O => \N__18332\,
            I => \N__18329\
        );

    \I__4251\ : Odrv4
    port map (
            O => \N__18329\,
            I => \M_current_address_qZ0Z_3\
        );

    \I__4250\ : CEMux
    port map (
            O => \N__18326\,
            I => \N__18322\
        );

    \I__4249\ : CEMux
    port map (
            O => \N__18325\,
            I => \N__18319\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__18322\,
            I => \N__18311\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__18319\,
            I => \N__18311\
        );

    \I__4246\ : CEMux
    port map (
            O => \N__18318\,
            I => \N__18308\
        );

    \I__4245\ : CEMux
    port map (
            O => \N__18317\,
            I => \N__18305\
        );

    \I__4244\ : CEMux
    port map (
            O => \N__18316\,
            I => \N__18302\
        );

    \I__4243\ : Span4Mux_v
    port map (
            O => \N__18311\,
            I => \N__18296\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__18308\,
            I => \N__18296\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__18305\,
            I => \N__18291\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__18302\,
            I => \N__18291\
        );

    \I__4239\ : CEMux
    port map (
            O => \N__18301\,
            I => \N__18288\
        );

    \I__4238\ : Span4Mux_v
    port map (
            O => \N__18296\,
            I => \N__18281\
        );

    \I__4237\ : Span4Mux_v
    port map (
            O => \N__18291\,
            I => \N__18281\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__18288\,
            I => \N__18281\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__18281\,
            I => \M_current_address_q_0_0\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__18278\,
            I => \N__18275\
        );

    \I__4233\ : CascadeBuf
    port map (
            O => \N__18275\,
            I => \N__18272\
        );

    \I__4232\ : CascadeMux
    port map (
            O => \N__18272\,
            I => \N__18269\
        );

    \I__4231\ : CascadeBuf
    port map (
            O => \N__18269\,
            I => \N__18266\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__18266\,
            I => \N__18263\
        );

    \I__4229\ : CascadeBuf
    port map (
            O => \N__18263\,
            I => \N__18260\
        );

    \I__4228\ : CascadeMux
    port map (
            O => \N__18260\,
            I => \N__18257\
        );

    \I__4227\ : CascadeBuf
    port map (
            O => \N__18257\,
            I => \N__18254\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__18254\,
            I => \N__18251\
        );

    \I__4225\ : CascadeBuf
    port map (
            O => \N__18251\,
            I => \N__18248\
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__18248\,
            I => \N__18245\
        );

    \I__4223\ : CascadeBuf
    port map (
            O => \N__18245\,
            I => \N__18242\
        );

    \I__4222\ : CascadeMux
    port map (
            O => \N__18242\,
            I => \N__18239\
        );

    \I__4221\ : CascadeBuf
    port map (
            O => \N__18239\,
            I => \N__18236\
        );

    \I__4220\ : CascadeMux
    port map (
            O => \N__18236\,
            I => \N__18233\
        );

    \I__4219\ : CascadeBuf
    port map (
            O => \N__18233\,
            I => \N__18230\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__18230\,
            I => \N__18227\
        );

    \I__4217\ : CascadeBuf
    port map (
            O => \N__18227\,
            I => \N__18224\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__18224\,
            I => \N__18221\
        );

    \I__4215\ : CascadeBuf
    port map (
            O => \N__18221\,
            I => \N__18218\
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__18218\,
            I => \N__18215\
        );

    \I__4213\ : CascadeBuf
    port map (
            O => \N__18215\,
            I => \N__18212\
        );

    \I__4212\ : CascadeMux
    port map (
            O => \N__18212\,
            I => \N__18209\
        );

    \I__4211\ : CascadeBuf
    port map (
            O => \N__18209\,
            I => \N__18206\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__18206\,
            I => \N__18203\
        );

    \I__4209\ : CascadeBuf
    port map (
            O => \N__18203\,
            I => \N__18200\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__18200\,
            I => \N__18197\
        );

    \I__4207\ : CascadeBuf
    port map (
            O => \N__18197\,
            I => \N__18194\
        );

    \I__4206\ : CascadeMux
    port map (
            O => \N__18194\,
            I => \N__18191\
        );

    \I__4205\ : CascadeBuf
    port map (
            O => \N__18191\,
            I => \N__18188\
        );

    \I__4204\ : CascadeMux
    port map (
            O => \N__18188\,
            I => \N__18185\
        );

    \I__4203\ : InMux
    port map (
            O => \N__18185\,
            I => \N__18182\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__4201\ : Span4Mux_s1_v
    port map (
            O => \N__18179\,
            I => \N__18176\
        );

    \I__4200\ : Odrv4
    port map (
            O => \N__18176\,
            I => \M_current_address_qZ0Z_10\
        );

    \I__4199\ : CascadeMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__4198\ : InMux
    port map (
            O => \N__18170\,
            I => \N__18166\
        );

    \I__4197\ : InMux
    port map (
            O => \N__18169\,
            I => \N__18163\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__18166\,
            I => \N__18160\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__18163\,
            I => \N__18157\
        );

    \I__4194\ : Span4Mux_v
    port map (
            O => \N__18160\,
            I => \N__18151\
        );

    \I__4193\ : Span4Mux_v
    port map (
            O => \N__18157\,
            I => \N__18151\
        );

    \I__4192\ : InMux
    port map (
            O => \N__18156\,
            I => \N__18148\
        );

    \I__4191\ : Sp12to4
    port map (
            O => \N__18151\,
            I => \N__18143\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__18148\,
            I => \N__18143\
        );

    \I__4189\ : Span12Mux_h
    port map (
            O => \N__18143\,
            I => \N__18140\
        );

    \I__4188\ : Odrv12
    port map (
            O => \N__18140\,
            I => port_data_c_0
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__18137\,
            I => \N__18134\
        );

    \I__4186\ : CascadeBuf
    port map (
            O => \N__18134\,
            I => \N__18131\
        );

    \I__4185\ : CascadeMux
    port map (
            O => \N__18131\,
            I => \N__18128\
        );

    \I__4184\ : CascadeBuf
    port map (
            O => \N__18128\,
            I => \N__18125\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__18125\,
            I => \N__18122\
        );

    \I__4182\ : CascadeBuf
    port map (
            O => \N__18122\,
            I => \N__18119\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__18119\,
            I => \N__18116\
        );

    \I__4180\ : CascadeBuf
    port map (
            O => \N__18116\,
            I => \N__18113\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__18113\,
            I => \N__18110\
        );

    \I__4178\ : CascadeBuf
    port map (
            O => \N__18110\,
            I => \N__18107\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__18107\,
            I => \N__18104\
        );

    \I__4176\ : CascadeBuf
    port map (
            O => \N__18104\,
            I => \N__18101\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__18101\,
            I => \N__18098\
        );

    \I__4174\ : CascadeBuf
    port map (
            O => \N__18098\,
            I => \N__18095\
        );

    \I__4173\ : CascadeMux
    port map (
            O => \N__18095\,
            I => \N__18092\
        );

    \I__4172\ : CascadeBuf
    port map (
            O => \N__18092\,
            I => \N__18089\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__4170\ : CascadeBuf
    port map (
            O => \N__18086\,
            I => \N__18083\
        );

    \I__4169\ : CascadeMux
    port map (
            O => \N__18083\,
            I => \N__18080\
        );

    \I__4168\ : CascadeBuf
    port map (
            O => \N__18080\,
            I => \N__18077\
        );

    \I__4167\ : CascadeMux
    port map (
            O => \N__18077\,
            I => \N__18074\
        );

    \I__4166\ : CascadeBuf
    port map (
            O => \N__18074\,
            I => \N__18071\
        );

    \I__4165\ : CascadeMux
    port map (
            O => \N__18071\,
            I => \N__18068\
        );

    \I__4164\ : CascadeBuf
    port map (
            O => \N__18068\,
            I => \N__18065\
        );

    \I__4163\ : CascadeMux
    port map (
            O => \N__18065\,
            I => \N__18062\
        );

    \I__4162\ : CascadeBuf
    port map (
            O => \N__18062\,
            I => \N__18059\
        );

    \I__4161\ : CascadeMux
    port map (
            O => \N__18059\,
            I => \N__18056\
        );

    \I__4160\ : CascadeBuf
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__18053\,
            I => \N__18050\
        );

    \I__4158\ : CascadeBuf
    port map (
            O => \N__18050\,
            I => \N__18047\
        );

    \I__4157\ : CascadeMux
    port map (
            O => \N__18047\,
            I => \N__18044\
        );

    \I__4156\ : InMux
    port map (
            O => \N__18044\,
            I => \N__18041\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__18041\,
            I => \N__18038\
        );

    \I__4154\ : Span4Mux_s1_v
    port map (
            O => \N__18038\,
            I => \N__18035\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__18035\,
            I => \M_current_address_qZ0Z_7\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__18032\,
            I => \N__18028\
        );

    \I__4151\ : InMux
    port map (
            O => \N__18031\,
            I => \N__18025\
        );

    \I__4150\ : InMux
    port map (
            O => \N__18028\,
            I => \N__18022\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__18025\,
            I => \N__18018\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__18022\,
            I => \N__18015\
        );

    \I__4147\ : InMux
    port map (
            O => \N__18021\,
            I => \N__18012\
        );

    \I__4146\ : Span4Mux_v
    port map (
            O => \N__18018\,
            I => \N__18009\
        );

    \I__4145\ : Span4Mux_v
    port map (
            O => \N__18015\,
            I => \N__18006\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__18012\,
            I => \N__18003\
        );

    \I__4143\ : Sp12to4
    port map (
            O => \N__18009\,
            I => \N__17998\
        );

    \I__4142\ : Sp12to4
    port map (
            O => \N__18006\,
            I => \N__17998\
        );

    \I__4141\ : Span12Mux_h
    port map (
            O => \N__18003\,
            I => \N__17995\
        );

    \I__4140\ : Span12Mux_h
    port map (
            O => \N__17998\,
            I => \N__17992\
        );

    \I__4139\ : Odrv12
    port map (
            O => \N__17995\,
            I => port_data_c_1
        );

    \I__4138\ : Odrv12
    port map (
            O => \N__17992\,
            I => port_data_c_1
        );

    \I__4137\ : CascadeMux
    port map (
            O => \N__17987\,
            I => \N__17984\
        );

    \I__4136\ : CascadeBuf
    port map (
            O => \N__17984\,
            I => \N__17981\
        );

    \I__4135\ : CascadeMux
    port map (
            O => \N__17981\,
            I => \N__17978\
        );

    \I__4134\ : CascadeBuf
    port map (
            O => \N__17978\,
            I => \N__17975\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__17975\,
            I => \N__17972\
        );

    \I__4132\ : CascadeBuf
    port map (
            O => \N__17972\,
            I => \N__17969\
        );

    \I__4131\ : CascadeMux
    port map (
            O => \N__17969\,
            I => \N__17966\
        );

    \I__4130\ : CascadeBuf
    port map (
            O => \N__17966\,
            I => \N__17963\
        );

    \I__4129\ : CascadeMux
    port map (
            O => \N__17963\,
            I => \N__17960\
        );

    \I__4128\ : CascadeBuf
    port map (
            O => \N__17960\,
            I => \N__17957\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__17957\,
            I => \N__17954\
        );

    \I__4126\ : CascadeBuf
    port map (
            O => \N__17954\,
            I => \N__17951\
        );

    \I__4125\ : CascadeMux
    port map (
            O => \N__17951\,
            I => \N__17948\
        );

    \I__4124\ : CascadeBuf
    port map (
            O => \N__17948\,
            I => \N__17945\
        );

    \I__4123\ : CascadeMux
    port map (
            O => \N__17945\,
            I => \N__17942\
        );

    \I__4122\ : CascadeBuf
    port map (
            O => \N__17942\,
            I => \N__17939\
        );

    \I__4121\ : CascadeMux
    port map (
            O => \N__17939\,
            I => \N__17936\
        );

    \I__4120\ : CascadeBuf
    port map (
            O => \N__17936\,
            I => \N__17933\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__17933\,
            I => \N__17930\
        );

    \I__4118\ : CascadeBuf
    port map (
            O => \N__17930\,
            I => \N__17927\
        );

    \I__4117\ : CascadeMux
    port map (
            O => \N__17927\,
            I => \N__17924\
        );

    \I__4116\ : CascadeBuf
    port map (
            O => \N__17924\,
            I => \N__17921\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__17921\,
            I => \N__17918\
        );

    \I__4114\ : CascadeBuf
    port map (
            O => \N__17918\,
            I => \N__17915\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__17915\,
            I => \N__17912\
        );

    \I__4112\ : CascadeBuf
    port map (
            O => \N__17912\,
            I => \N__17909\
        );

    \I__4111\ : CascadeMux
    port map (
            O => \N__17909\,
            I => \N__17906\
        );

    \I__4110\ : CascadeBuf
    port map (
            O => \N__17906\,
            I => \N__17903\
        );

    \I__4109\ : CascadeMux
    port map (
            O => \N__17903\,
            I => \N__17900\
        );

    \I__4108\ : CascadeBuf
    port map (
            O => \N__17900\,
            I => \N__17897\
        );

    \I__4107\ : CascadeMux
    port map (
            O => \N__17897\,
            I => \N__17894\
        );

    \I__4106\ : InMux
    port map (
            O => \N__17894\,
            I => \N__17891\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__17891\,
            I => \N__17888\
        );

    \I__4104\ : Odrv4
    port map (
            O => \N__17888\,
            I => \M_current_address_qZ0Z_8\
        );

    \I__4103\ : CEMux
    port map (
            O => \N__17885\,
            I => \N__17882\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__17882\,
            I => \N__17876\
        );

    \I__4101\ : CEMux
    port map (
            O => \N__17881\,
            I => \N__17873\
        );

    \I__4100\ : CEMux
    port map (
            O => \N__17880\,
            I => \N__17870\
        );

    \I__4099\ : CEMux
    port map (
            O => \N__17879\,
            I => \N__17865\
        );

    \I__4098\ : Span4Mux_v
    port map (
            O => \N__17876\,
            I => \N__17860\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__17873\,
            I => \N__17860\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__17870\,
            I => \N__17857\
        );

    \I__4095\ : CEMux
    port map (
            O => \N__17869\,
            I => \N__17854\
        );

    \I__4094\ : CEMux
    port map (
            O => \N__17868\,
            I => \N__17851\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__17865\,
            I => \N__17846\
        );

    \I__4092\ : Sp12to4
    port map (
            O => \N__17860\,
            I => \N__17846\
        );

    \I__4091\ : Span4Mux_h
    port map (
            O => \N__17857\,
            I => \N__17843\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__17854\,
            I => \N__17840\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__17851\,
            I => \N__17837\
        );

    \I__4088\ : Span12Mux_v
    port map (
            O => \N__17846\,
            I => \N__17834\
        );

    \I__4087\ : Span4Mux_v
    port map (
            O => \N__17843\,
            I => \N__17831\
        );

    \I__4086\ : Span4Mux_h
    port map (
            O => \N__17840\,
            I => \N__17828\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__17837\,
            I => \N__17825\
        );

    \I__4084\ : Odrv12
    port map (
            O => \N__17834\,
            I => \M_current_address_q_0_6_0\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__17831\,
            I => \M_current_address_q_0_6_0\
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__17828\,
            I => \M_current_address_q_0_6_0\
        );

    \I__4081\ : Odrv4
    port map (
            O => \N__17825\,
            I => \M_current_address_q_0_6_0\
        );

    \I__4080\ : InMux
    port map (
            O => \N__17816\,
            I => \N__17812\
        );

    \I__4079\ : InMux
    port map (
            O => \N__17815\,
            I => \N__17809\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__17812\,
            I => \N__17788\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__17809\,
            I => \N__17785\
        );

    \I__4076\ : SRMux
    port map (
            O => \N__17808\,
            I => \N__17744\
        );

    \I__4075\ : SRMux
    port map (
            O => \N__17807\,
            I => \N__17744\
        );

    \I__4074\ : SRMux
    port map (
            O => \N__17806\,
            I => \N__17744\
        );

    \I__4073\ : SRMux
    port map (
            O => \N__17805\,
            I => \N__17744\
        );

    \I__4072\ : SRMux
    port map (
            O => \N__17804\,
            I => \N__17744\
        );

    \I__4071\ : SRMux
    port map (
            O => \N__17803\,
            I => \N__17744\
        );

    \I__4070\ : SRMux
    port map (
            O => \N__17802\,
            I => \N__17744\
        );

    \I__4069\ : SRMux
    port map (
            O => \N__17801\,
            I => \N__17744\
        );

    \I__4068\ : SRMux
    port map (
            O => \N__17800\,
            I => \N__17744\
        );

    \I__4067\ : SRMux
    port map (
            O => \N__17799\,
            I => \N__17744\
        );

    \I__4066\ : SRMux
    port map (
            O => \N__17798\,
            I => \N__17744\
        );

    \I__4065\ : SRMux
    port map (
            O => \N__17797\,
            I => \N__17744\
        );

    \I__4064\ : SRMux
    port map (
            O => \N__17796\,
            I => \N__17744\
        );

    \I__4063\ : SRMux
    port map (
            O => \N__17795\,
            I => \N__17744\
        );

    \I__4062\ : SRMux
    port map (
            O => \N__17794\,
            I => \N__17744\
        );

    \I__4061\ : SRMux
    port map (
            O => \N__17793\,
            I => \N__17744\
        );

    \I__4060\ : SRMux
    port map (
            O => \N__17792\,
            I => \N__17744\
        );

    \I__4059\ : SRMux
    port map (
            O => \N__17791\,
            I => \N__17744\
        );

    \I__4058\ : Glb2LocalMux
    port map (
            O => \N__17788\,
            I => \N__17744\
        );

    \I__4057\ : Glb2LocalMux
    port map (
            O => \N__17785\,
            I => \N__17744\
        );

    \I__4056\ : GlobalMux
    port map (
            O => \N__17744\,
            I => \N__17741\
        );

    \I__4055\ : gio2CtrlBuf
    port map (
            O => \N__17741\,
            I => \N_631_g\
        );

    \I__4054\ : InMux
    port map (
            O => \N__17738\,
            I => \N__17735\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__17735\,
            I => \N__17732\
        );

    \I__4052\ : Span4Mux_h
    port map (
            O => \N__17732\,
            I => \N__17729\
        );

    \I__4051\ : Sp12to4
    port map (
            O => \N__17729\,
            I => \N__17726\
        );

    \I__4050\ : Span12Mux_s10_v
    port map (
            O => \N__17726\,
            I => \N__17721\
        );

    \I__4049\ : InMux
    port map (
            O => \N__17725\,
            I => \N__17715\
        );

    \I__4048\ : InMux
    port map (
            O => \N__17724\,
            I => \N__17715\
        );

    \I__4047\ : Span12Mux_v
    port map (
            O => \N__17721\,
            I => \N__17712\
        );

    \I__4046\ : InMux
    port map (
            O => \N__17720\,
            I => \N__17709\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__17715\,
            I => \N__17706\
        );

    \I__4044\ : Odrv12
    port map (
            O => \N__17712\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_2\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__17709\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_2\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__17706\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_2\
        );

    \I__4041\ : InMux
    port map (
            O => \N__17699\,
            I => \N__17696\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__17696\,
            I => \N__17693\
        );

    \I__4039\ : Span4Mux_v
    port map (
            O => \N__17693\,
            I => \N__17690\
        );

    \I__4038\ : Sp12to4
    port map (
            O => \N__17690\,
            I => \N__17687\
        );

    \I__4037\ : Span12Mux_h
    port map (
            O => \N__17687\,
            I => \N__17684\
        );

    \I__4036\ : Span12Mux_v
    port map (
            O => \N__17684\,
            I => \N__17680\
        );

    \I__4035\ : InMux
    port map (
            O => \N__17683\,
            I => \N__17677\
        );

    \I__4034\ : Odrv12
    port map (
            O => \N__17680\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__17677\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__4032\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17669\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__17669\,
            I => \N__17666\
        );

    \I__4030\ : Span4Mux_h
    port map (
            O => \N__17666\,
            I => \N__17663\
        );

    \I__4029\ : Span4Mux_h
    port map (
            O => \N__17663\,
            I => \N__17659\
        );

    \I__4028\ : InMux
    port map (
            O => \N__17662\,
            I => \N__17655\
        );

    \I__4027\ : Sp12to4
    port map (
            O => \N__17659\,
            I => \N__17651\
        );

    \I__4026\ : InMux
    port map (
            O => \N__17658\,
            I => \N__17648\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__17655\,
            I => \N__17645\
        );

    \I__4024\ : InMux
    port map (
            O => \N__17654\,
            I => \N__17640\
        );

    \I__4023\ : Span12Mux_v
    port map (
            O => \N__17651\,
            I => \N__17633\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__17648\,
            I => \N__17630\
        );

    \I__4021\ : Span4Mux_h
    port map (
            O => \N__17645\,
            I => \N__17627\
        );

    \I__4020\ : InMux
    port map (
            O => \N__17644\,
            I => \N__17622\
        );

    \I__4019\ : InMux
    port map (
            O => \N__17643\,
            I => \N__17622\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__17640\,
            I => \N__17619\
        );

    \I__4017\ : InMux
    port map (
            O => \N__17639\,
            I => \N__17614\
        );

    \I__4016\ : InMux
    port map (
            O => \N__17638\,
            I => \N__17614\
        );

    \I__4015\ : InMux
    port map (
            O => \N__17637\,
            I => \N__17611\
        );

    \I__4014\ : InMux
    port map (
            O => \N__17636\,
            I => \N__17608\
        );

    \I__4013\ : Odrv12
    port map (
            O => \N__17633\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0\
        );

    \I__4012\ : Odrv4
    port map (
            O => \N__17630\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0\
        );

    \I__4011\ : Odrv4
    port map (
            O => \N__17627\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__17622\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0\
        );

    \I__4009\ : Odrv4
    port map (
            O => \N__17619\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__17614\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__17611\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__17608\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0\
        );

    \I__4005\ : CascadeMux
    port map (
            O => \N__17591\,
            I => \N__17588\
        );

    \I__4004\ : CascadeBuf
    port map (
            O => \N__17588\,
            I => \N__17585\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__17585\,
            I => \N__17582\
        );

    \I__4002\ : CascadeBuf
    port map (
            O => \N__17582\,
            I => \N__17579\
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__17579\,
            I => \N__17576\
        );

    \I__4000\ : CascadeBuf
    port map (
            O => \N__17576\,
            I => \N__17573\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__3998\ : CascadeBuf
    port map (
            O => \N__17570\,
            I => \N__17567\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__17567\,
            I => \N__17564\
        );

    \I__3996\ : CascadeBuf
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__3995\ : CascadeMux
    port map (
            O => \N__17561\,
            I => \N__17558\
        );

    \I__3994\ : CascadeBuf
    port map (
            O => \N__17558\,
            I => \N__17555\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__17555\,
            I => \N__17552\
        );

    \I__3992\ : CascadeBuf
    port map (
            O => \N__17552\,
            I => \N__17549\
        );

    \I__3991\ : CascadeMux
    port map (
            O => \N__17549\,
            I => \N__17546\
        );

    \I__3990\ : CascadeBuf
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__17543\,
            I => \N__17540\
        );

    \I__3988\ : CascadeBuf
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__3987\ : CascadeMux
    port map (
            O => \N__17537\,
            I => \N__17534\
        );

    \I__3986\ : CascadeBuf
    port map (
            O => \N__17534\,
            I => \N__17531\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__17531\,
            I => \N__17528\
        );

    \I__3984\ : CascadeBuf
    port map (
            O => \N__17528\,
            I => \N__17525\
        );

    \I__3983\ : CascadeMux
    port map (
            O => \N__17525\,
            I => \N__17522\
        );

    \I__3982\ : CascadeBuf
    port map (
            O => \N__17522\,
            I => \N__17519\
        );

    \I__3981\ : CascadeMux
    port map (
            O => \N__17519\,
            I => \N__17516\
        );

    \I__3980\ : CascadeBuf
    port map (
            O => \N__17516\,
            I => \N__17513\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__17513\,
            I => \N__17510\
        );

    \I__3978\ : CascadeBuf
    port map (
            O => \N__17510\,
            I => \N__17507\
        );

    \I__3977\ : CascadeMux
    port map (
            O => \N__17507\,
            I => \N__17504\
        );

    \I__3976\ : CascadeBuf
    port map (
            O => \N__17504\,
            I => \N__17501\
        );

    \I__3975\ : CascadeMux
    port map (
            O => \N__17501\,
            I => \N__17498\
        );

    \I__3974\ : InMux
    port map (
            O => \N__17498\,
            I => \N__17495\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__17495\,
            I => this_vga_signals_un14_address_if_generate_plus_mult1_un61_sum_i_3
        );

    \I__3972\ : InMux
    port map (
            O => \N__17492\,
            I => \N__17488\
        );

    \I__3971\ : InMux
    port map (
            O => \N__17491\,
            I => \N__17485\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__17488\,
            I => \N__17480\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__17485\,
            I => \N__17480\
        );

    \I__3968\ : Span12Mux_v
    port map (
            O => \N__17480\,
            I => \N__17477\
        );

    \I__3967\ : Odrv12
    port map (
            O => \N__17477\,
            I => port_data_c_6
        );

    \I__3966\ : CascadeMux
    port map (
            O => \N__17474\,
            I => \N__17471\
        );

    \I__3965\ : CascadeBuf
    port map (
            O => \N__17471\,
            I => \N__17468\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__17468\,
            I => \N__17465\
        );

    \I__3963\ : CascadeBuf
    port map (
            O => \N__17465\,
            I => \N__17462\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__17462\,
            I => \N__17459\
        );

    \I__3961\ : CascadeBuf
    port map (
            O => \N__17459\,
            I => \N__17456\
        );

    \I__3960\ : CascadeMux
    port map (
            O => \N__17456\,
            I => \N__17453\
        );

    \I__3959\ : CascadeBuf
    port map (
            O => \N__17453\,
            I => \N__17450\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__17450\,
            I => \N__17447\
        );

    \I__3957\ : CascadeBuf
    port map (
            O => \N__17447\,
            I => \N__17444\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__17444\,
            I => \N__17441\
        );

    \I__3955\ : CascadeBuf
    port map (
            O => \N__17441\,
            I => \N__17438\
        );

    \I__3954\ : CascadeMux
    port map (
            O => \N__17438\,
            I => \N__17435\
        );

    \I__3953\ : CascadeBuf
    port map (
            O => \N__17435\,
            I => \N__17432\
        );

    \I__3952\ : CascadeMux
    port map (
            O => \N__17432\,
            I => \N__17429\
        );

    \I__3951\ : CascadeBuf
    port map (
            O => \N__17429\,
            I => \N__17426\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__17426\,
            I => \N__17423\
        );

    \I__3949\ : CascadeBuf
    port map (
            O => \N__17423\,
            I => \N__17420\
        );

    \I__3948\ : CascadeMux
    port map (
            O => \N__17420\,
            I => \N__17417\
        );

    \I__3947\ : CascadeBuf
    port map (
            O => \N__17417\,
            I => \N__17414\
        );

    \I__3946\ : CascadeMux
    port map (
            O => \N__17414\,
            I => \N__17411\
        );

    \I__3945\ : CascadeBuf
    port map (
            O => \N__17411\,
            I => \N__17408\
        );

    \I__3944\ : CascadeMux
    port map (
            O => \N__17408\,
            I => \N__17405\
        );

    \I__3943\ : CascadeBuf
    port map (
            O => \N__17405\,
            I => \N__17402\
        );

    \I__3942\ : CascadeMux
    port map (
            O => \N__17402\,
            I => \N__17399\
        );

    \I__3941\ : CascadeBuf
    port map (
            O => \N__17399\,
            I => \N__17396\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__17396\,
            I => \N__17393\
        );

    \I__3939\ : CascadeBuf
    port map (
            O => \N__17393\,
            I => \N__17390\
        );

    \I__3938\ : CascadeMux
    port map (
            O => \N__17390\,
            I => \N__17387\
        );

    \I__3937\ : CascadeBuf
    port map (
            O => \N__17387\,
            I => \N__17384\
        );

    \I__3936\ : CascadeMux
    port map (
            O => \N__17384\,
            I => \N__17381\
        );

    \I__3935\ : InMux
    port map (
            O => \N__17381\,
            I => \N__17378\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__17378\,
            I => \N__17375\
        );

    \I__3933\ : Span12Mux_s2_v
    port map (
            O => \N__17375\,
            I => \N__17372\
        );

    \I__3932\ : Span12Mux_v
    port map (
            O => \N__17372\,
            I => \N__17369\
        );

    \I__3931\ : Odrv12
    port map (
            O => \N__17369\,
            I => \M_current_address_qZ0Z_6\
        );

    \I__3930\ : CEMux
    port map (
            O => \N__17366\,
            I => \N__17363\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__17363\,
            I => \N__17359\
        );

    \I__3928\ : CEMux
    port map (
            O => \N__17362\,
            I => \N__17356\
        );

    \I__3927\ : Span4Mux_v
    port map (
            O => \N__17359\,
            I => \N__17351\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__17356\,
            I => \N__17351\
        );

    \I__3925\ : Odrv4
    port map (
            O => \N__17351\,
            I => \this_vram.mem_WE_4\
        );

    \I__3924\ : InMux
    port map (
            O => \N__17348\,
            I => \N__17341\
        );

    \I__3923\ : InMux
    port map (
            O => \N__17347\,
            I => \N__17338\
        );

    \I__3922\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17331\
        );

    \I__3921\ : InMux
    port map (
            O => \N__17345\,
            I => \N__17331\
        );

    \I__3920\ : InMux
    port map (
            O => \N__17344\,
            I => \N__17331\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__17341\,
            I => \N__17327\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__17338\,
            I => \N__17322\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__17331\,
            I => \N__17322\
        );

    \I__3916\ : InMux
    port map (
            O => \N__17330\,
            I => \N__17319\
        );

    \I__3915\ : Span4Mux_h
    port map (
            O => \N__17327\,
            I => \N__17314\
        );

    \I__3914\ : Span4Mux_v
    port map (
            O => \N__17322\,
            I => \N__17309\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__17319\,
            I => \N__17309\
        );

    \I__3912\ : InMux
    port map (
            O => \N__17318\,
            I => \N__17304\
        );

    \I__3911\ : InMux
    port map (
            O => \N__17317\,
            I => \N__17304\
        );

    \I__3910\ : Odrv4
    port map (
            O => \N__17314\,
            I => \M_current_address_qZ0Z_12\
        );

    \I__3909\ : Odrv4
    port map (
            O => \N__17309\,
            I => \M_current_address_qZ0Z_12\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__17304\,
            I => \M_current_address_qZ0Z_12\
        );

    \I__3907\ : CascadeMux
    port map (
            O => \N__17297\,
            I => \N__17294\
        );

    \I__3906\ : InMux
    port map (
            O => \N__17294\,
            I => \N__17285\
        );

    \I__3905\ : CascadeMux
    port map (
            O => \N__17293\,
            I => \N__17281\
        );

    \I__3904\ : CascadeMux
    port map (
            O => \N__17292\,
            I => \N__17278\
        );

    \I__3903\ : CascadeMux
    port map (
            O => \N__17291\,
            I => \N__17275\
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__17290\,
            I => \N__17272\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__17289\,
            I => \N__17269\
        );

    \I__3900\ : CascadeMux
    port map (
            O => \N__17288\,
            I => \N__17266\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__17285\,
            I => \N__17263\
        );

    \I__3898\ : CascadeMux
    port map (
            O => \N__17284\,
            I => \N__17260\
        );

    \I__3897\ : InMux
    port map (
            O => \N__17281\,
            I => \N__17255\
        );

    \I__3896\ : InMux
    port map (
            O => \N__17278\,
            I => \N__17255\
        );

    \I__3895\ : InMux
    port map (
            O => \N__17275\,
            I => \N__17252\
        );

    \I__3894\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17245\
        );

    \I__3893\ : InMux
    port map (
            O => \N__17269\,
            I => \N__17245\
        );

    \I__3892\ : InMux
    port map (
            O => \N__17266\,
            I => \N__17245\
        );

    \I__3891\ : Span4Mux_h
    port map (
            O => \N__17263\,
            I => \N__17242\
        );

    \I__3890\ : InMux
    port map (
            O => \N__17260\,
            I => \N__17239\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__17255\,
            I => \N__17232\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__17252\,
            I => \N__17232\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__17245\,
            I => \N__17232\
        );

    \I__3886\ : Odrv4
    port map (
            O => \N__17242\,
            I => \M_current_address_qZ0Z_13\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__17239\,
            I => \M_current_address_qZ0Z_13\
        );

    \I__3884\ : Odrv12
    port map (
            O => \N__17232\,
            I => \M_current_address_qZ0Z_13\
        );

    \I__3883\ : IoInMux
    port map (
            O => \N__17225\,
            I => \N__17222\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__17222\,
            I => \N__17219\
        );

    \I__3881\ : IoSpan4Mux
    port map (
            O => \N__17219\,
            I => \N__17210\
        );

    \I__3880\ : InMux
    port map (
            O => \N__17218\,
            I => \N__17207\
        );

    \I__3879\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17202\
        );

    \I__3878\ : InMux
    port map (
            O => \N__17216\,
            I => \N__17202\
        );

    \I__3877\ : InMux
    port map (
            O => \N__17215\,
            I => \N__17195\
        );

    \I__3876\ : InMux
    port map (
            O => \N__17214\,
            I => \N__17195\
        );

    \I__3875\ : InMux
    port map (
            O => \N__17213\,
            I => \N__17195\
        );

    \I__3874\ : IoSpan4Mux
    port map (
            O => \N__17210\,
            I => \N__17191\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__17207\,
            I => \N__17188\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__17202\,
            I => \N__17185\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__17195\,
            I => \N__17182\
        );

    \I__3870\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17179\
        );

    \I__3869\ : Sp12to4
    port map (
            O => \N__17191\,
            I => \N__17175\
        );

    \I__3868\ : Span4Mux_v
    port map (
            O => \N__17188\,
            I => \N__17172\
        );

    \I__3867\ : Span4Mux_h
    port map (
            O => \N__17185\,
            I => \N__17169\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__17182\,
            I => \N__17164\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__17179\,
            I => \N__17164\
        );

    \I__3864\ : InMux
    port map (
            O => \N__17178\,
            I => \N__17161\
        );

    \I__3863\ : Span12Mux_s9_v
    port map (
            O => \N__17175\,
            I => \N__17157\
        );

    \I__3862\ : Span4Mux_h
    port map (
            O => \N__17172\,
            I => \N__17154\
        );

    \I__3861\ : Span4Mux_h
    port map (
            O => \N__17169\,
            I => \N__17151\
        );

    \I__3860\ : Span4Mux_v
    port map (
            O => \N__17164\,
            I => \N__17146\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__17161\,
            I => \N__17146\
        );

    \I__3858\ : InMux
    port map (
            O => \N__17160\,
            I => \N__17143\
        );

    \I__3857\ : Odrv12
    port map (
            O => \N__17157\,
            I => debug_c
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__17154\,
            I => debug_c
        );

    \I__3855\ : Odrv4
    port map (
            O => \N__17151\,
            I => debug_c
        );

    \I__3854\ : Odrv4
    port map (
            O => \N__17146\,
            I => debug_c
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__17143\,
            I => debug_c
        );

    \I__3852\ : CEMux
    port map (
            O => \N__17132\,
            I => \N__17129\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__17129\,
            I => \N__17125\
        );

    \I__3850\ : CEMux
    port map (
            O => \N__17128\,
            I => \N__17122\
        );

    \I__3849\ : Span4Mux_s2_v
    port map (
            O => \N__17125\,
            I => \N__17117\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__17122\,
            I => \N__17117\
        );

    \I__3847\ : Span4Mux_v
    port map (
            O => \N__17117\,
            I => \N__17114\
        );

    \I__3846\ : Span4Mux_v
    port map (
            O => \N__17114\,
            I => \N__17111\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__17111\,
            I => \this_vram.mem_WE_0\
        );

    \I__3844\ : InMux
    port map (
            O => \N__17108\,
            I => \N__17105\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__17105\,
            I => \N__17102\
        );

    \I__3842\ : Span4Mux_v
    port map (
            O => \N__17102\,
            I => \N__17098\
        );

    \I__3841\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17095\
        );

    \I__3840\ : Span4Mux_h
    port map (
            O => \N__17098\,
            I => \N__17092\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__17095\,
            I => \N__17089\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__17092\,
            I => port_data_c_5
        );

    \I__3837\ : Odrv12
    port map (
            O => \N__17089\,
            I => port_data_c_5
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__17084\,
            I => \N__17081\
        );

    \I__3835\ : CascadeBuf
    port map (
            O => \N__17081\,
            I => \N__17078\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__17078\,
            I => \N__17075\
        );

    \I__3833\ : CascadeBuf
    port map (
            O => \N__17075\,
            I => \N__17072\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__17072\,
            I => \N__17069\
        );

    \I__3831\ : CascadeBuf
    port map (
            O => \N__17069\,
            I => \N__17066\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__17066\,
            I => \N__17063\
        );

    \I__3829\ : CascadeBuf
    port map (
            O => \N__17063\,
            I => \N__17060\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__17060\,
            I => \N__17057\
        );

    \I__3827\ : CascadeBuf
    port map (
            O => \N__17057\,
            I => \N__17054\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__17054\,
            I => \N__17051\
        );

    \I__3825\ : CascadeBuf
    port map (
            O => \N__17051\,
            I => \N__17048\
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__17048\,
            I => \N__17045\
        );

    \I__3823\ : CascadeBuf
    port map (
            O => \N__17045\,
            I => \N__17042\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__17042\,
            I => \N__17039\
        );

    \I__3821\ : CascadeBuf
    port map (
            O => \N__17039\,
            I => \N__17036\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__17036\,
            I => \N__17033\
        );

    \I__3819\ : CascadeBuf
    port map (
            O => \N__17033\,
            I => \N__17030\
        );

    \I__3818\ : CascadeMux
    port map (
            O => \N__17030\,
            I => \N__17027\
        );

    \I__3817\ : CascadeBuf
    port map (
            O => \N__17027\,
            I => \N__17024\
        );

    \I__3816\ : CascadeMux
    port map (
            O => \N__17024\,
            I => \N__17021\
        );

    \I__3815\ : CascadeBuf
    port map (
            O => \N__17021\,
            I => \N__17018\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__17018\,
            I => \N__17015\
        );

    \I__3813\ : CascadeBuf
    port map (
            O => \N__17015\,
            I => \N__17012\
        );

    \I__3812\ : CascadeMux
    port map (
            O => \N__17012\,
            I => \N__17009\
        );

    \I__3811\ : CascadeBuf
    port map (
            O => \N__17009\,
            I => \N__17006\
        );

    \I__3810\ : CascadeMux
    port map (
            O => \N__17006\,
            I => \N__17003\
        );

    \I__3809\ : CascadeBuf
    port map (
            O => \N__17003\,
            I => \N__17000\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__17000\,
            I => \N__16997\
        );

    \I__3807\ : CascadeBuf
    port map (
            O => \N__16997\,
            I => \N__16994\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__16994\,
            I => \N__16991\
        );

    \I__3805\ : InMux
    port map (
            O => \N__16991\,
            I => \N__16988\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__16988\,
            I => \N__16985\
        );

    \I__3803\ : Span4Mux_s1_v
    port map (
            O => \N__16985\,
            I => \N__16982\
        );

    \I__3802\ : Span4Mux_v
    port map (
            O => \N__16982\,
            I => \N__16979\
        );

    \I__3801\ : Span4Mux_v
    port map (
            O => \N__16979\,
            I => \N__16976\
        );

    \I__3800\ : Odrv4
    port map (
            O => \N__16976\,
            I => \M_current_address_qZ0Z_5\
        );

    \I__3799\ : InMux
    port map (
            O => \N__16973\,
            I => \N__16969\
        );

    \I__3798\ : InMux
    port map (
            O => \N__16972\,
            I => \N__16962\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__16969\,
            I => \N__16959\
        );

    \I__3796\ : InMux
    port map (
            O => \N__16968\,
            I => \N__16956\
        );

    \I__3795\ : InMux
    port map (
            O => \N__16967\,
            I => \N__16947\
        );

    \I__3794\ : InMux
    port map (
            O => \N__16966\,
            I => \N__16947\
        );

    \I__3793\ : InMux
    port map (
            O => \N__16965\,
            I => \N__16947\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__16962\,
            I => \N__16944\
        );

    \I__3791\ : Span4Mux_v
    port map (
            O => \N__16959\,
            I => \N__16939\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__16956\,
            I => \N__16939\
        );

    \I__3789\ : InMux
    port map (
            O => \N__16955\,
            I => \N__16934\
        );

    \I__3788\ : InMux
    port map (
            O => \N__16954\,
            I => \N__16934\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__16947\,
            I => \N__16931\
        );

    \I__3786\ : Span4Mux_h
    port map (
            O => \N__16944\,
            I => \N__16928\
        );

    \I__3785\ : Span4Mux_v
    port map (
            O => \N__16939\,
            I => \N__16923\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__16934\,
            I => \N__16923\
        );

    \I__3783\ : Odrv12
    port map (
            O => \N__16931\,
            I => \M_current_address_qZ0Z_11\
        );

    \I__3782\ : Odrv4
    port map (
            O => \N__16928\,
            I => \M_current_address_qZ0Z_11\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__16923\,
            I => \M_current_address_qZ0Z_11\
        );

    \I__3780\ : InMux
    port map (
            O => \N__16916\,
            I => \N__16913\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__16913\,
            I => \N__16909\
        );

    \I__3778\ : InMux
    port map (
            O => \N__16912\,
            I => \N__16906\
        );

    \I__3777\ : Span4Mux_v
    port map (
            O => \N__16909\,
            I => \N__16901\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__16906\,
            I => \N__16901\
        );

    \I__3775\ : Span4Mux_h
    port map (
            O => \N__16901\,
            I => \N__16898\
        );

    \I__3774\ : Span4Mux_v
    port map (
            O => \N__16898\,
            I => \N__16895\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__16895\,
            I => \N__16892\
        );

    \I__3772\ : Odrv4
    port map (
            O => \N__16892\,
            I => port_data_c_4
        );

    \I__3771\ : CascadeMux
    port map (
            O => \N__16889\,
            I => \N__16886\
        );

    \I__3770\ : CascadeBuf
    port map (
            O => \N__16886\,
            I => \N__16883\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__16883\,
            I => \N__16880\
        );

    \I__3768\ : CascadeBuf
    port map (
            O => \N__16880\,
            I => \N__16877\
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__16877\,
            I => \N__16874\
        );

    \I__3766\ : CascadeBuf
    port map (
            O => \N__16874\,
            I => \N__16871\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__16871\,
            I => \N__16868\
        );

    \I__3764\ : CascadeBuf
    port map (
            O => \N__16868\,
            I => \N__16865\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__16865\,
            I => \N__16862\
        );

    \I__3762\ : CascadeBuf
    port map (
            O => \N__16862\,
            I => \N__16859\
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__16859\,
            I => \N__16856\
        );

    \I__3760\ : CascadeBuf
    port map (
            O => \N__16856\,
            I => \N__16853\
        );

    \I__3759\ : CascadeMux
    port map (
            O => \N__16853\,
            I => \N__16850\
        );

    \I__3758\ : CascadeBuf
    port map (
            O => \N__16850\,
            I => \N__16847\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__16847\,
            I => \N__16844\
        );

    \I__3756\ : CascadeBuf
    port map (
            O => \N__16844\,
            I => \N__16841\
        );

    \I__3755\ : CascadeMux
    port map (
            O => \N__16841\,
            I => \N__16838\
        );

    \I__3754\ : CascadeBuf
    port map (
            O => \N__16838\,
            I => \N__16835\
        );

    \I__3753\ : CascadeMux
    port map (
            O => \N__16835\,
            I => \N__16832\
        );

    \I__3752\ : CascadeBuf
    port map (
            O => \N__16832\,
            I => \N__16829\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__16829\,
            I => \N__16826\
        );

    \I__3750\ : CascadeBuf
    port map (
            O => \N__16826\,
            I => \N__16823\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__16823\,
            I => \N__16820\
        );

    \I__3748\ : CascadeBuf
    port map (
            O => \N__16820\,
            I => \N__16817\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__16817\,
            I => \N__16814\
        );

    \I__3746\ : CascadeBuf
    port map (
            O => \N__16814\,
            I => \N__16811\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__16811\,
            I => \N__16808\
        );

    \I__3744\ : CascadeBuf
    port map (
            O => \N__16808\,
            I => \N__16805\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__16805\,
            I => \N__16802\
        );

    \I__3742\ : CascadeBuf
    port map (
            O => \N__16802\,
            I => \N__16799\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__16799\,
            I => \N__16796\
        );

    \I__3740\ : InMux
    port map (
            O => \N__16796\,
            I => \N__16793\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__16793\,
            I => \N__16790\
        );

    \I__3738\ : Span4Mux_s2_v
    port map (
            O => \N__16790\,
            I => \N__16787\
        );

    \I__3737\ : Span4Mux_v
    port map (
            O => \N__16787\,
            I => \N__16784\
        );

    \I__3736\ : Odrv4
    port map (
            O => \N__16784\,
            I => \M_current_address_qZ0Z_4\
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__16781\,
            I => \this_vram.mem_mem_1_1_RNIUSK11Z0Z_0_cascade_\
        );

    \I__3734\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16775\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__16775\,
            I => \N__16772\
        );

    \I__3732\ : Span4Mux_h
    port map (
            O => \N__16772\,
            I => \N__16769\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__16769\,
            I => \this_vram.mem_N_102\
        );

    \I__3730\ : InMux
    port map (
            O => \N__16766\,
            I => \N__16763\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__16763\,
            I => \N__16760\
        );

    \I__3728\ : Span4Mux_v
    port map (
            O => \N__16760\,
            I => \N__16757\
        );

    \I__3727\ : Span4Mux_v
    port map (
            O => \N__16757\,
            I => \N__16754\
        );

    \I__3726\ : Odrv4
    port map (
            O => \N__16754\,
            I => \this_vram.mem_out_bus1_2\
        );

    \I__3725\ : InMux
    port map (
            O => \N__16751\,
            I => \N__16748\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__16748\,
            I => \N__16745\
        );

    \I__3723\ : Sp12to4
    port map (
            O => \N__16745\,
            I => \N__16742\
        );

    \I__3722\ : Span12Mux_v
    port map (
            O => \N__16742\,
            I => \N__16739\
        );

    \I__3721\ : Odrv12
    port map (
            O => \N__16739\,
            I => \this_vram.mem_out_bus5_2\
        );

    \I__3720\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16725\
        );

    \I__3719\ : InMux
    port map (
            O => \N__16735\,
            I => \N__16725\
        );

    \I__3718\ : InMux
    port map (
            O => \N__16734\,
            I => \N__16722\
        );

    \I__3717\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16717\
        );

    \I__3716\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16717\
        );

    \I__3715\ : InMux
    port map (
            O => \N__16731\,
            I => \N__16712\
        );

    \I__3714\ : InMux
    port map (
            O => \N__16730\,
            I => \N__16712\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__16725\,
            I => \N__16704\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__16722\,
            I => \N__16704\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__16717\,
            I => \N__16704\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__16712\,
            I => \N__16701\
        );

    \I__3709\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16698\
        );

    \I__3708\ : Span4Mux_v
    port map (
            O => \N__16704\,
            I => \N__16691\
        );

    \I__3707\ : Span4Mux_v
    port map (
            O => \N__16701\,
            I => \N__16691\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__16698\,
            I => \N__16691\
        );

    \I__3705\ : Odrv4
    port map (
            O => \N__16691\,
            I => \this_vram.mem_radregZ0Z_12\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__16688\,
            I => \this_vram.mem_mem_1_1_RNIUSKZ0Z11_cascade_\
        );

    \I__3703\ : InMux
    port map (
            O => \N__16685\,
            I => \N__16682\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__16682\,
            I => \this_vram.mem_N_95\
        );

    \I__3701\ : InMux
    port map (
            O => \N__16679\,
            I => \N__16676\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__16676\,
            I => \N__16673\
        );

    \I__3699\ : Span4Mux_h
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__3698\ : Odrv4
    port map (
            O => \N__16670\,
            I => \this_vram.mem_out_bus3_0\
        );

    \I__3697\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16664\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__16664\,
            I => \N__16661\
        );

    \I__3695\ : Sp12to4
    port map (
            O => \N__16661\,
            I => \N__16658\
        );

    \I__3694\ : Span12Mux_v
    port map (
            O => \N__16658\,
            I => \N__16655\
        );

    \I__3693\ : Odrv12
    port map (
            O => \N__16655\,
            I => \this_vram.mem_out_bus7_0\
        );

    \I__3692\ : InMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__3690\ : Span4Mux_v
    port map (
            O => \N__16646\,
            I => \N__16643\
        );

    \I__3689\ : Odrv4
    port map (
            O => \N__16643\,
            I => \this_vram.mem_mem_3_0_RNI05PZ0Z11\
        );

    \I__3688\ : CEMux
    port map (
            O => \N__16640\,
            I => \N__16637\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__16637\,
            I => \N__16633\
        );

    \I__3686\ : CEMux
    port map (
            O => \N__16636\,
            I => \N__16630\
        );

    \I__3685\ : Span4Mux_v
    port map (
            O => \N__16633\,
            I => \N__16625\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__16630\,
            I => \N__16625\
        );

    \I__3683\ : Span4Mux_h
    port map (
            O => \N__16625\,
            I => \N__16622\
        );

    \I__3682\ : Odrv4
    port map (
            O => \N__16622\,
            I => \this_vram.mem_WE_10\
        );

    \I__3681\ : CEMux
    port map (
            O => \N__16619\,
            I => \N__16616\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__16616\,
            I => \N__16613\
        );

    \I__3679\ : Span12Mux_s8_h
    port map (
            O => \N__16613\,
            I => \N__16609\
        );

    \I__3678\ : CEMux
    port map (
            O => \N__16612\,
            I => \N__16606\
        );

    \I__3677\ : Odrv12
    port map (
            O => \N__16609\,
            I => \this_vram.mem_WE_8\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__16606\,
            I => \this_vram.mem_WE_8\
        );

    \I__3675\ : CEMux
    port map (
            O => \N__16601\,
            I => \N__16598\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__16598\,
            I => \N__16594\
        );

    \I__3673\ : CEMux
    port map (
            O => \N__16597\,
            I => \N__16591\
        );

    \I__3672\ : Span4Mux_s1_v
    port map (
            O => \N__16594\,
            I => \N__16586\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__16591\,
            I => \N__16586\
        );

    \I__3670\ : Span4Mux_v
    port map (
            O => \N__16586\,
            I => \N__16583\
        );

    \I__3669\ : Span4Mux_v
    port map (
            O => \N__16583\,
            I => \N__16580\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__16580\,
            I => \this_vram.mem_WE_14\
        );

    \I__3667\ : InMux
    port map (
            O => \N__16577\,
            I => \N__16574\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__16574\,
            I => \N__16571\
        );

    \I__3665\ : Span4Mux_v
    port map (
            O => \N__16571\,
            I => \N__16568\
        );

    \I__3664\ : Span4Mux_v
    port map (
            O => \N__16568\,
            I => \N__16565\
        );

    \I__3663\ : Sp12to4
    port map (
            O => \N__16565\,
            I => \N__16562\
        );

    \I__3662\ : Odrv12
    port map (
            O => \N__16562\,
            I => \this_vram.mem_out_bus7_3\
        );

    \I__3661\ : InMux
    port map (
            O => \N__16559\,
            I => \N__16556\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__16556\,
            I => \this_vram.mem_out_bus3_3\
        );

    \I__3659\ : InMux
    port map (
            O => \N__16553\,
            I => \N__16550\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__16550\,
            I => \N__16547\
        );

    \I__3657\ : Odrv4
    port map (
            O => \N__16547\,
            I => \this_vram.mem_mem_3_1_RNI25P11Z0Z_0\
        );

    \I__3656\ : InMux
    port map (
            O => \N__16544\,
            I => \N__16541\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__16541\,
            I => \this_vram.mem_out_bus3_2\
        );

    \I__3654\ : InMux
    port map (
            O => \N__16538\,
            I => \N__16535\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__16535\,
            I => \N__16532\
        );

    \I__3652\ : Span4Mux_v
    port map (
            O => \N__16532\,
            I => \N__16529\
        );

    \I__3651\ : Span4Mux_v
    port map (
            O => \N__16529\,
            I => \N__16526\
        );

    \I__3650\ : Sp12to4
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__3649\ : Odrv12
    port map (
            O => \N__16523\,
            I => \this_vram.mem_out_bus7_2\
        );

    \I__3648\ : InMux
    port map (
            O => \N__16520\,
            I => \N__16516\
        );

    \I__3647\ : InMux
    port map (
            O => \N__16519\,
            I => \N__16509\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__16516\,
            I => \N__16502\
        );

    \I__3645\ : InMux
    port map (
            O => \N__16515\,
            I => \N__16497\
        );

    \I__3644\ : InMux
    port map (
            O => \N__16514\,
            I => \N__16497\
        );

    \I__3643\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16492\
        );

    \I__3642\ : InMux
    port map (
            O => \N__16512\,
            I => \N__16492\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__16509\,
            I => \N__16489\
        );

    \I__3640\ : InMux
    port map (
            O => \N__16508\,
            I => \N__16480\
        );

    \I__3639\ : InMux
    port map (
            O => \N__16507\,
            I => \N__16480\
        );

    \I__3638\ : InMux
    port map (
            O => \N__16506\,
            I => \N__16480\
        );

    \I__3637\ : InMux
    port map (
            O => \N__16505\,
            I => \N__16480\
        );

    \I__3636\ : Span4Mux_v
    port map (
            O => \N__16502\,
            I => \N__16469\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__16497\,
            I => \N__16469\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__16492\,
            I => \N__16466\
        );

    \I__3633\ : Span4Mux_v
    port map (
            O => \N__16489\,
            I => \N__16461\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__16480\,
            I => \N__16461\
        );

    \I__3631\ : InMux
    port map (
            O => \N__16479\,
            I => \N__16452\
        );

    \I__3630\ : InMux
    port map (
            O => \N__16478\,
            I => \N__16452\
        );

    \I__3629\ : InMux
    port map (
            O => \N__16477\,
            I => \N__16452\
        );

    \I__3628\ : InMux
    port map (
            O => \N__16476\,
            I => \N__16452\
        );

    \I__3627\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16447\
        );

    \I__3626\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16447\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__16469\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__16466\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__16461\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__16452\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__16447\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__3620\ : InMux
    port map (
            O => \N__16436\,
            I => \N__16433\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__16433\,
            I => \N__16430\
        );

    \I__3618\ : Odrv12
    port map (
            O => \N__16430\,
            I => \this_vram.mem_mem_3_1_RNI25PZ0Z11\
        );

    \I__3617\ : CascadeMux
    port map (
            O => \N__16427\,
            I => \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0_cascade_\
        );

    \I__3616\ : InMux
    port map (
            O => \N__16424\,
            I => \N__16421\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__16421\,
            I => \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0\
        );

    \I__3614\ : InMux
    port map (
            O => \N__16418\,
            I => \N__16415\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__16415\,
            I => \N__16412\
        );

    \I__3612\ : Span4Mux_v
    port map (
            O => \N__16412\,
            I => \N__16409\
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__16409\,
            I => \this_vram.mem_N_91\
        );

    \I__3610\ : InMux
    port map (
            O => \N__16406\,
            I => \N__16402\
        );

    \I__3609\ : InMux
    port map (
            O => \N__16405\,
            I => \N__16398\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__16402\,
            I => \N__16395\
        );

    \I__3607\ : InMux
    port map (
            O => \N__16401\,
            I => \N__16392\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__16398\,
            I => \N__16387\
        );

    \I__3605\ : Span4Mux_h
    port map (
            O => \N__16395\,
            I => \N__16387\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__16392\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKMEZ0\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__16387\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKMEZ0\
        );

    \I__3602\ : CascadeMux
    port map (
            O => \N__16382\,
            I => \N__16379\
        );

    \I__3601\ : InMux
    port map (
            O => \N__16379\,
            I => \N__16372\
        );

    \I__3600\ : InMux
    port map (
            O => \N__16378\,
            I => \N__16372\
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__16377\,
            I => \N__16366\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__16372\,
            I => \N__16360\
        );

    \I__3597\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16357\
        );

    \I__3596\ : InMux
    port map (
            O => \N__16370\,
            I => \N__16353\
        );

    \I__3595\ : InMux
    port map (
            O => \N__16369\,
            I => \N__16350\
        );

    \I__3594\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16342\
        );

    \I__3593\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16339\
        );

    \I__3592\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16334\
        );

    \I__3591\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16334\
        );

    \I__3590\ : Span4Mux_v
    port map (
            O => \N__16360\,
            I => \N__16329\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__16357\,
            I => \N__16329\
        );

    \I__3588\ : InMux
    port map (
            O => \N__16356\,
            I => \N__16326\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__16353\,
            I => \N__16321\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__16350\,
            I => \N__16321\
        );

    \I__3585\ : InMux
    port map (
            O => \N__16349\,
            I => \N__16314\
        );

    \I__3584\ : InMux
    port map (
            O => \N__16348\,
            I => \N__16314\
        );

    \I__3583\ : InMux
    port map (
            O => \N__16347\,
            I => \N__16314\
        );

    \I__3582\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16311\
        );

    \I__3581\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16305\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__16342\,
            I => \N__16300\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__16339\,
            I => \N__16300\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__16334\,
            I => \N__16297\
        );

    \I__3577\ : Span4Mux_h
    port map (
            O => \N__16329\,
            I => \N__16294\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__16326\,
            I => \N__16290\
        );

    \I__3575\ : Span4Mux_v
    port map (
            O => \N__16321\,
            I => \N__16285\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__16314\,
            I => \N__16285\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__16311\,
            I => \N__16282\
        );

    \I__3572\ : InMux
    port map (
            O => \N__16310\,
            I => \N__16275\
        );

    \I__3571\ : InMux
    port map (
            O => \N__16309\,
            I => \N__16275\
        );

    \I__3570\ : InMux
    port map (
            O => \N__16308\,
            I => \N__16275\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__16305\,
            I => \N__16272\
        );

    \I__3568\ : Span4Mux_v
    port map (
            O => \N__16300\,
            I => \N__16267\
        );

    \I__3567\ : Span4Mux_v
    port map (
            O => \N__16297\,
            I => \N__16267\
        );

    \I__3566\ : Span4Mux_h
    port map (
            O => \N__16294\,
            I => \N__16264\
        );

    \I__3565\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16261\
        );

    \I__3564\ : Span4Mux_v
    port map (
            O => \N__16290\,
            I => \N__16252\
        );

    \I__3563\ : Span4Mux_h
    port map (
            O => \N__16285\,
            I => \N__16252\
        );

    \I__3562\ : Span4Mux_v
    port map (
            O => \N__16282\,
            I => \N__16252\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__16275\,
            I => \N__16252\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__16272\,
            I => \this_vga_signals.M_vaddress_qZ0Z_5\
        );

    \I__3559\ : Odrv4
    port map (
            O => \N__16267\,
            I => \this_vga_signals.M_vaddress_qZ0Z_5\
        );

    \I__3558\ : Odrv4
    port map (
            O => \N__16264\,
            I => \this_vga_signals.M_vaddress_qZ0Z_5\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__16261\,
            I => \this_vga_signals.M_vaddress_qZ0Z_5\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__16252\,
            I => \this_vga_signals.M_vaddress_qZ0Z_5\
        );

    \I__3555\ : SRMux
    port map (
            O => \N__16241\,
            I => \N__16220\
        );

    \I__3554\ : SRMux
    port map (
            O => \N__16240\,
            I => \N__16220\
        );

    \I__3553\ : SRMux
    port map (
            O => \N__16239\,
            I => \N__16220\
        );

    \I__3552\ : SRMux
    port map (
            O => \N__16238\,
            I => \N__16220\
        );

    \I__3551\ : SRMux
    port map (
            O => \N__16237\,
            I => \N__16220\
        );

    \I__3550\ : SRMux
    port map (
            O => \N__16236\,
            I => \N__16220\
        );

    \I__3549\ : SRMux
    port map (
            O => \N__16235\,
            I => \N__16220\
        );

    \I__3548\ : GlobalMux
    port map (
            O => \N__16220\,
            I => \N__16217\
        );

    \I__3547\ : gio2CtrlBuf
    port map (
            O => \N__16217\,
            I => \this_vga_signals.N_583_g\
        );

    \I__3546\ : InMux
    port map (
            O => \N__16214\,
            I => \N__16211\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__16211\,
            I => \N__16208\
        );

    \I__3544\ : Sp12to4
    port map (
            O => \N__16208\,
            I => \N__16205\
        );

    \I__3543\ : Span12Mux_v
    port map (
            O => \N__16205\,
            I => \N__16202\
        );

    \I__3542\ : Span12Mux_v
    port map (
            O => \N__16202\,
            I => \N__16199\
        );

    \I__3541\ : Odrv12
    port map (
            O => \N__16199\,
            I => \this_vram.mem_out_bus6_3\
        );

    \I__3540\ : InMux
    port map (
            O => \N__16196\,
            I => \N__16193\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__16193\,
            I => \this_vram.mem_out_bus2_3\
        );

    \I__3538\ : CascadeMux
    port map (
            O => \N__16190\,
            I => \this_vram.mem_mem_2_1_RNI01N11Z0Z_0_cascade_\
        );

    \I__3537\ : InMux
    port map (
            O => \N__16187\,
            I => \N__16184\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__16184\,
            I => \N__16181\
        );

    \I__3535\ : Span4Mux_h
    port map (
            O => \N__16181\,
            I => \N__16178\
        );

    \I__3534\ : Odrv4
    port map (
            O => \N__16178\,
            I => \this_vram.mem_N_105\
        );

    \I__3533\ : InMux
    port map (
            O => \N__16175\,
            I => \N__16172\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__16172\,
            I => \N__16169\
        );

    \I__3531\ : Span4Mux_v
    port map (
            O => \N__16169\,
            I => \N__16166\
        );

    \I__3530\ : Span4Mux_v
    port map (
            O => \N__16166\,
            I => \N__16163\
        );

    \I__3529\ : Odrv4
    port map (
            O => \N__16163\,
            I => \this_vram.mem_out_bus0_3\
        );

    \I__3528\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16157\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__16157\,
            I => \N__16154\
        );

    \I__3526\ : Span4Mux_v
    port map (
            O => \N__16154\,
            I => \N__16151\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__16151\,
            I => \this_vram.mem_out_bus4_3\
        );

    \I__3524\ : InMux
    port map (
            O => \N__16148\,
            I => \N__16145\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__16145\,
            I => \this_vram.mem_mem_0_1_RNISOI11Z0Z_0\
        );

    \I__3522\ : CEMux
    port map (
            O => \N__16142\,
            I => \N__16139\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__16139\,
            I => \N__16135\
        );

    \I__3520\ : CEMux
    port map (
            O => \N__16138\,
            I => \N__16132\
        );

    \I__3519\ : Span4Mux_v
    port map (
            O => \N__16135\,
            I => \N__16127\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__16132\,
            I => \N__16127\
        );

    \I__3517\ : Span4Mux_v
    port map (
            O => \N__16127\,
            I => \N__16124\
        );

    \I__3516\ : Odrv4
    port map (
            O => \N__16124\,
            I => \this_vram.mem_WE_12\
        );

    \I__3515\ : InMux
    port map (
            O => \N__16121\,
            I => \N__16118\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__16118\,
            I => \N__16115\
        );

    \I__3513\ : Span4Mux_v
    port map (
            O => \N__16115\,
            I => \N__16112\
        );

    \I__3512\ : Span4Mux_v
    port map (
            O => \N__16112\,
            I => \N__16109\
        );

    \I__3511\ : Sp12to4
    port map (
            O => \N__16109\,
            I => \N__16106\
        );

    \I__3510\ : Odrv12
    port map (
            O => \N__16106\,
            I => \this_vram.mem_out_bus7_1\
        );

    \I__3509\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16100\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__16100\,
            I => \this_vram.mem_out_bus3_1\
        );

    \I__3507\ : InMux
    port map (
            O => \N__16097\,
            I => \N__16094\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__16094\,
            I => \N__16091\
        );

    \I__3505\ : Odrv12
    port map (
            O => \N__16091\,
            I => \this_vram.mem_mem_3_0_RNI05P11Z0Z_0\
        );

    \I__3504\ : InMux
    port map (
            O => \N__16088\,
            I => \N__16085\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__16085\,
            I => \N__16082\
        );

    \I__3502\ : Sp12to4
    port map (
            O => \N__16082\,
            I => \N__16079\
        );

    \I__3501\ : Span12Mux_v
    port map (
            O => \N__16079\,
            I => \N__16076\
        );

    \I__3500\ : Odrv12
    port map (
            O => \N__16076\,
            I => \this_vram.mem_out_bus5_3\
        );

    \I__3499\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16070\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__16070\,
            I => \N__16067\
        );

    \I__3497\ : Span4Mux_v
    port map (
            O => \N__16067\,
            I => \N__16064\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__16064\,
            I => \this_vram.mem_out_bus1_3\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__16061\,
            I => \N__16058\
        );

    \I__3494\ : InMux
    port map (
            O => \N__16058\,
            I => \N__16055\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__16055\,
            I => \this_vram.mem_out_bus2_0\
        );

    \I__3492\ : InMux
    port map (
            O => \N__16052\,
            I => \N__16049\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__16049\,
            I => \N__16046\
        );

    \I__3490\ : Span4Mux_v
    port map (
            O => \N__16046\,
            I => \N__16043\
        );

    \I__3489\ : Span4Mux_v
    port map (
            O => \N__16043\,
            I => \N__16040\
        );

    \I__3488\ : Sp12to4
    port map (
            O => \N__16040\,
            I => \N__16037\
        );

    \I__3487\ : Odrv12
    port map (
            O => \N__16037\,
            I => \this_vram.mem_out_bus6_0\
        );

    \I__3486\ : InMux
    port map (
            O => \N__16034\,
            I => \N__16031\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__16031\,
            I => \this_vram.mem_mem_2_0_RNIU0NZ0Z11\
        );

    \I__3484\ : InMux
    port map (
            O => \N__16028\,
            I => \N__16025\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__16025\,
            I => \N__16022\
        );

    \I__3482\ : Span4Mux_v
    port map (
            O => \N__16022\,
            I => \N__16019\
        );

    \I__3481\ : Odrv4
    port map (
            O => \N__16019\,
            I => \this_vram.mem_out_bus1_1\
        );

    \I__3480\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16013\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__16013\,
            I => \N__16010\
        );

    \I__3478\ : Sp12to4
    port map (
            O => \N__16010\,
            I => \N__16007\
        );

    \I__3477\ : Span12Mux_v
    port map (
            O => \N__16007\,
            I => \N__16004\
        );

    \I__3476\ : Odrv12
    port map (
            O => \N__16004\,
            I => \this_vram.mem_out_bus5_1\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__16001\,
            I => \this_vram.mem_mem_1_0_RNISSK11Z0Z_0_cascade_\
        );

    \I__3474\ : InMux
    port map (
            O => \N__15998\,
            I => \N__15995\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__15995\,
            I => \N__15992\
        );

    \I__3472\ : Odrv4
    port map (
            O => \N__15992\,
            I => \this_vram.mem_N_88\
        );

    \I__3471\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15986\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__15986\,
            I => \N__15983\
        );

    \I__3469\ : Sp12to4
    port map (
            O => \N__15983\,
            I => \N__15980\
        );

    \I__3468\ : Span12Mux_v
    port map (
            O => \N__15980\,
            I => \N__15977\
        );

    \I__3467\ : Odrv12
    port map (
            O => \N__15977\,
            I => \this_vram.mem_out_bus4_2\
        );

    \I__3466\ : InMux
    port map (
            O => \N__15974\,
            I => \N__15971\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__15971\,
            I => \N__15968\
        );

    \I__3464\ : Span4Mux_v
    port map (
            O => \N__15968\,
            I => \N__15965\
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__15965\,
            I => \this_vram.mem_out_bus0_2\
        );

    \I__3462\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15959\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__15959\,
            I => \N__15956\
        );

    \I__3460\ : Sp12to4
    port map (
            O => \N__15956\,
            I => \N__15953\
        );

    \I__3459\ : Span12Mux_v
    port map (
            O => \N__15953\,
            I => \N__15950\
        );

    \I__3458\ : Span12Mux_v
    port map (
            O => \N__15950\,
            I => \N__15947\
        );

    \I__3457\ : Odrv12
    port map (
            O => \N__15947\,
            I => \this_vram.mem_out_bus6_2\
        );

    \I__3456\ : InMux
    port map (
            O => \N__15944\,
            I => \N__15941\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__15941\,
            I => \N__15938\
        );

    \I__3454\ : Odrv4
    port map (
            O => \N__15938\,
            I => \this_vram.mem_out_bus2_2\
        );

    \I__3453\ : InMux
    port map (
            O => \N__15935\,
            I => \N__15932\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__15932\,
            I => \this_vram.mem_mem_0_1_RNISOIZ0Z11\
        );

    \I__3451\ : CascadeMux
    port map (
            O => \N__15929\,
            I => \this_vram.mem_mem_2_1_RNI01NZ0Z11_cascade_\
        );

    \I__3450\ : InMux
    port map (
            O => \N__15926\,
            I => \N__15923\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__15923\,
            I => \N__15920\
        );

    \I__3448\ : Odrv4
    port map (
            O => \N__15920\,
            I => \this_vram.mem_N_98\
        );

    \I__3447\ : InMux
    port map (
            O => \N__15917\,
            I => \N__15914\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__15914\,
            I => \N__15911\
        );

    \I__3445\ : Sp12to4
    port map (
            O => \N__15911\,
            I => \N__15908\
        );

    \I__3444\ : Span12Mux_v
    port map (
            O => \N__15908\,
            I => \N__15905\
        );

    \I__3443\ : Odrv12
    port map (
            O => \N__15905\,
            I => \this_vram.mem_out_bus6_1\
        );

    \I__3442\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15899\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__15899\,
            I => \this_vram.mem_out_bus2_1\
        );

    \I__3440\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15893\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__15893\,
            I => \N__15890\
        );

    \I__3438\ : Span4Mux_v
    port map (
            O => \N__15890\,
            I => \N__15887\
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__15887\,
            I => \this_vram.mem_out_bus4_1\
        );

    \I__3436\ : InMux
    port map (
            O => \N__15884\,
            I => \N__15881\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__15881\,
            I => \N__15878\
        );

    \I__3434\ : Span4Mux_v
    port map (
            O => \N__15878\,
            I => \N__15875\
        );

    \I__3433\ : Span4Mux_v
    port map (
            O => \N__15875\,
            I => \N__15872\
        );

    \I__3432\ : Odrv4
    port map (
            O => \N__15872\,
            I => \this_vram.mem_out_bus0_1\
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__15869\,
            I => \N__15866\
        );

    \I__3430\ : InMux
    port map (
            O => \N__15866\,
            I => \N__15860\
        );

    \I__3429\ : InMux
    port map (
            O => \N__15865\,
            I => \N__15857\
        );

    \I__3428\ : InMux
    port map (
            O => \N__15864\,
            I => \N__15852\
        );

    \I__3427\ : CascadeMux
    port map (
            O => \N__15863\,
            I => \N__15849\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__15860\,
            I => \N__15844\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__15857\,
            I => \N__15844\
        );

    \I__3424\ : InMux
    port map (
            O => \N__15856\,
            I => \N__15841\
        );

    \I__3423\ : CascadeMux
    port map (
            O => \N__15855\,
            I => \N__15838\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__15852\,
            I => \N__15835\
        );

    \I__3421\ : InMux
    port map (
            O => \N__15849\,
            I => \N__15832\
        );

    \I__3420\ : Span4Mux_v
    port map (
            O => \N__15844\,
            I => \N__15827\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__15841\,
            I => \N__15827\
        );

    \I__3418\ : InMux
    port map (
            O => \N__15838\,
            I => \N__15824\
        );

    \I__3417\ : Span4Mux_v
    port map (
            O => \N__15835\,
            I => \N__15821\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__15832\,
            I => \N__15814\
        );

    \I__3415\ : Sp12to4
    port map (
            O => \N__15827\,
            I => \N__15814\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__15824\,
            I => \N__15814\
        );

    \I__3413\ : Sp12to4
    port map (
            O => \N__15821\,
            I => \N__15811\
        );

    \I__3412\ : Span12Mux_v
    port map (
            O => \N__15814\,
            I => \N__15808\
        );

    \I__3411\ : Span12Mux_h
    port map (
            O => \N__15811\,
            I => \N__15803\
        );

    \I__3410\ : Span12Mux_h
    port map (
            O => \N__15808\,
            I => \N__15803\
        );

    \I__3409\ : Odrv12
    port map (
            O => \N__15803\,
            I => \M_this_vram_read_data_2\
        );

    \I__3408\ : CEMux
    port map (
            O => \N__15800\,
            I => \N__15796\
        );

    \I__3407\ : CEMux
    port map (
            O => \N__15799\,
            I => \N__15793\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__15796\,
            I => \N__15788\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__15793\,
            I => \N__15788\
        );

    \I__3404\ : Span4Mux_v
    port map (
            O => \N__15788\,
            I => \N__15785\
        );

    \I__3403\ : Span4Mux_h
    port map (
            O => \N__15785\,
            I => \N__15782\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__15782\,
            I => \this_vram.mem_WE_6\
        );

    \I__3401\ : InMux
    port map (
            O => \N__15779\,
            I => \N__15776\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__15776\,
            I => \N__15773\
        );

    \I__3399\ : Odrv4
    port map (
            O => \N__15773\,
            I => \M_current_address_qZ1Z_0\
        );

    \I__3398\ : CascadeMux
    port map (
            O => \N__15770\,
            I => \N__15767\
        );

    \I__3397\ : CascadeBuf
    port map (
            O => \N__15767\,
            I => \N__15764\
        );

    \I__3396\ : CascadeMux
    port map (
            O => \N__15764\,
            I => \N__15761\
        );

    \I__3395\ : CascadeBuf
    port map (
            O => \N__15761\,
            I => \N__15758\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__15758\,
            I => \N__15755\
        );

    \I__3393\ : CascadeBuf
    port map (
            O => \N__15755\,
            I => \N__15752\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__15752\,
            I => \N__15749\
        );

    \I__3391\ : CascadeBuf
    port map (
            O => \N__15749\,
            I => \N__15746\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__15746\,
            I => \N__15743\
        );

    \I__3389\ : CascadeBuf
    port map (
            O => \N__15743\,
            I => \N__15740\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__15740\,
            I => \N__15737\
        );

    \I__3387\ : CascadeBuf
    port map (
            O => \N__15737\,
            I => \N__15734\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__15734\,
            I => \N__15731\
        );

    \I__3385\ : CascadeBuf
    port map (
            O => \N__15731\,
            I => \N__15728\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__15728\,
            I => \N__15725\
        );

    \I__3383\ : CascadeBuf
    port map (
            O => \N__15725\,
            I => \N__15722\
        );

    \I__3382\ : CascadeMux
    port map (
            O => \N__15722\,
            I => \N__15719\
        );

    \I__3381\ : CascadeBuf
    port map (
            O => \N__15719\,
            I => \N__15716\
        );

    \I__3380\ : CascadeMux
    port map (
            O => \N__15716\,
            I => \N__15713\
        );

    \I__3379\ : CascadeBuf
    port map (
            O => \N__15713\,
            I => \N__15710\
        );

    \I__3378\ : CascadeMux
    port map (
            O => \N__15710\,
            I => \N__15707\
        );

    \I__3377\ : CascadeBuf
    port map (
            O => \N__15707\,
            I => \N__15704\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__15704\,
            I => \N__15701\
        );

    \I__3375\ : CascadeBuf
    port map (
            O => \N__15701\,
            I => \N__15698\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__15698\,
            I => \N__15695\
        );

    \I__3373\ : CascadeBuf
    port map (
            O => \N__15695\,
            I => \N__15692\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__15692\,
            I => \N__15689\
        );

    \I__3371\ : CascadeBuf
    port map (
            O => \N__15689\,
            I => \N__15686\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__15686\,
            I => \N__15683\
        );

    \I__3369\ : CascadeBuf
    port map (
            O => \N__15683\,
            I => \N__15680\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__15680\,
            I => \N__15677\
        );

    \I__3367\ : InMux
    port map (
            O => \N__15677\,
            I => \N__15674\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__15674\,
            I => \N__15671\
        );

    \I__3365\ : Span4Mux_s1_v
    port map (
            O => \N__15671\,
            I => \N__15668\
        );

    \I__3364\ : Span4Mux_v
    port map (
            O => \N__15668\,
            I => \N__15665\
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__15665\,
            I => \M_current_address_qZ0Z_0\
        );

    \I__3362\ : InMux
    port map (
            O => \N__15662\,
            I => \N__15659\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__15659\,
            I => \N__15656\
        );

    \I__3360\ : Span4Mux_v
    port map (
            O => \N__15656\,
            I => \N__15653\
        );

    \I__3359\ : Span4Mux_v
    port map (
            O => \N__15653\,
            I => \N__15650\
        );

    \I__3358\ : Span4Mux_v
    port map (
            O => \N__15650\,
            I => \N__15647\
        );

    \I__3357\ : Odrv4
    port map (
            O => \N__15647\,
            I => \this_vram.mem_out_bus5_0\
        );

    \I__3356\ : InMux
    port map (
            O => \N__15644\,
            I => \N__15641\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__15641\,
            I => \this_vram.mem_out_bus1_0\
        );

    \I__3354\ : InMux
    port map (
            O => \N__15638\,
            I => \N__15635\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__15635\,
            I => \this_vram.mem_mem_1_0_RNISSKZ0Z11\
        );

    \I__3352\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15629\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__15629\,
            I => \N__15625\
        );

    \I__3350\ : InMux
    port map (
            O => \N__15628\,
            I => \N__15622\
        );

    \I__3349\ : Span4Mux_v
    port map (
            O => \N__15625\,
            I => \N__15618\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__15622\,
            I => \N__15615\
        );

    \I__3347\ : InMux
    port map (
            O => \N__15621\,
            I => \N__15612\
        );

    \I__3346\ : Span4Mux_h
    port map (
            O => \N__15618\,
            I => \N__15606\
        );

    \I__3345\ : Span4Mux_v
    port map (
            O => \N__15615\,
            I => \N__15606\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__15612\,
            I => \N__15603\
        );

    \I__3343\ : InMux
    port map (
            O => \N__15611\,
            I => \N__15600\
        );

    \I__3342\ : Odrv4
    port map (
            O => \N__15606\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__3341\ : Odrv12
    port map (
            O => \N__15603\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__15600\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__3339\ : CascadeMux
    port map (
            O => \N__15593\,
            I => \this_vram.mem_N_109_cascade_\
        );

    \I__3338\ : InMux
    port map (
            O => \N__15590\,
            I => \N__15585\
        );

    \I__3337\ : InMux
    port map (
            O => \N__15589\,
            I => \N__15581\
        );

    \I__3336\ : InMux
    port map (
            O => \N__15588\,
            I => \N__15578\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__15585\,
            I => \N__15575\
        );

    \I__3334\ : InMux
    port map (
            O => \N__15584\,
            I => \N__15572\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__15581\,
            I => \N__15567\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__15578\,
            I => \N__15567\
        );

    \I__3331\ : Span4Mux_v
    port map (
            O => \N__15575\,
            I => \N__15558\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__15572\,
            I => \N__15558\
        );

    \I__3329\ : Span4Mux_v
    port map (
            O => \N__15567\,
            I => \N__15558\
        );

    \I__3328\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15555\
        );

    \I__3327\ : InMux
    port map (
            O => \N__15565\,
            I => \N__15552\
        );

    \I__3326\ : Span4Mux_v
    port map (
            O => \N__15558\,
            I => \N__15547\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__15555\,
            I => \N__15547\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__15552\,
            I => \N__15544\
        );

    \I__3323\ : Span4Mux_v
    port map (
            O => \N__15547\,
            I => \N__15541\
        );

    \I__3322\ : Span12Mux_v
    port map (
            O => \N__15544\,
            I => \N__15538\
        );

    \I__3321\ : Sp12to4
    port map (
            O => \N__15541\,
            I => \N__15535\
        );

    \I__3320\ : Span12Mux_h
    port map (
            O => \N__15538\,
            I => \N__15532\
        );

    \I__3319\ : Span12Mux_h
    port map (
            O => \N__15535\,
            I => \N__15529\
        );

    \I__3318\ : Odrv12
    port map (
            O => \N__15532\,
            I => \M_this_vram_read_data_0\
        );

    \I__3317\ : Odrv12
    port map (
            O => \N__15529\,
            I => \M_this_vram_read_data_0\
        );

    \I__3316\ : InMux
    port map (
            O => \N__15524\,
            I => \N__15521\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__15521\,
            I => \N__15518\
        );

    \I__3314\ : Span4Mux_v
    port map (
            O => \N__15518\,
            I => \N__15515\
        );

    \I__3313\ : Odrv4
    port map (
            O => \N__15515\,
            I => \this_vram.mem_out_bus0_0\
        );

    \I__3312\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15509\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__15509\,
            I => \N__15506\
        );

    \I__3310\ : Sp12to4
    port map (
            O => \N__15506\,
            I => \N__15503\
        );

    \I__3309\ : Span12Mux_v
    port map (
            O => \N__15503\,
            I => \N__15500\
        );

    \I__3308\ : Odrv12
    port map (
            O => \N__15500\,
            I => \this_vram.mem_out_bus4_0\
        );

    \I__3307\ : CascadeMux
    port map (
            O => \N__15497\,
            I => \this_vram.mem_mem_0_0_RNIQOIZ0Z11_cascade_\
        );

    \I__3306\ : InMux
    port map (
            O => \N__15494\,
            I => \N__15491\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__15491\,
            I => \this_vram.mem_N_112\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__15488\,
            I => \this_vga_signals.g1_1_cascade_\
        );

    \I__3303\ : InMux
    port map (
            O => \N__15485\,
            I => \N__15482\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__15482\,
            I => \this_vga_signals.N_15_0_0\
        );

    \I__3301\ : InMux
    port map (
            O => \N__15479\,
            I => \N__15476\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__15476\,
            I => \this_vga_signals.N_353_0\
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__15473\,
            I => \this_vga_signals.N_3520_0_cascade_\
        );

    \I__3298\ : InMux
    port map (
            O => \N__15470\,
            I => \N__15463\
        );

    \I__3297\ : InMux
    port map (
            O => \N__15469\,
            I => \N__15460\
        );

    \I__3296\ : InMux
    port map (
            O => \N__15468\,
            I => \N__15447\
        );

    \I__3295\ : InMux
    port map (
            O => \N__15467\,
            I => \N__15447\
        );

    \I__3294\ : InMux
    port map (
            O => \N__15466\,
            I => \N__15444\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__15463\,
            I => \N__15439\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__15460\,
            I => \N__15439\
        );

    \I__3291\ : InMux
    port map (
            O => \N__15459\,
            I => \N__15434\
        );

    \I__3290\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15434\
        );

    \I__3289\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15429\
        );

    \I__3288\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15429\
        );

    \I__3287\ : InMux
    port map (
            O => \N__15455\,
            I => \N__15424\
        );

    \I__3286\ : InMux
    port map (
            O => \N__15454\,
            I => \N__15424\
        );

    \I__3285\ : InMux
    port map (
            O => \N__15453\,
            I => \N__15419\
        );

    \I__3284\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15419\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__15447\,
            I => \this_vga_signals.CO1_2_1\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__15444\,
            I => \this_vga_signals.CO1_2_1\
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__15439\,
            I => \this_vga_signals.CO1_2_1\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__15434\,
            I => \this_vga_signals.CO1_2_1\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__15429\,
            I => \this_vga_signals.CO1_2_1\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__15424\,
            I => \this_vga_signals.CO1_2_1\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__15419\,
            I => \this_vga_signals.CO1_2_1\
        );

    \I__3276\ : InMux
    port map (
            O => \N__15404\,
            I => \N__15401\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__15401\,
            I => \this_vga_signals.mult1_un40_sum_0_2\
        );

    \I__3274\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15392\
        );

    \I__3273\ : InMux
    port map (
            O => \N__15397\,
            I => \N__15392\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__15392\,
            I => \this_vga_signals.g0_1_N_2L1\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__15389\,
            I => \N__15386\
        );

    \I__3270\ : InMux
    port map (
            O => \N__15386\,
            I => \N__15383\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__15383\,
            I => \N__15380\
        );

    \I__3268\ : Span4Mux_h
    port map (
            O => \N__15380\,
            I => \N__15377\
        );

    \I__3267\ : Span4Mux_h
    port map (
            O => \N__15377\,
            I => \N__15373\
        );

    \I__3266\ : InMux
    port map (
            O => \N__15376\,
            I => \N__15370\
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__15373\,
            I => \this_vga_signals.N_1253_0\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__15370\,
            I => \this_vga_signals.N_1253_0\
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__15365\,
            I => \this_vga_signals.mult1_un40_sum_0_2_cascade_\
        );

    \I__3262\ : InMux
    port map (
            O => \N__15362\,
            I => \N__15356\
        );

    \I__3261\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15356\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__15356\,
            I => \this_vga_signals.N_3_0\
        );

    \I__3259\ : InMux
    port map (
            O => \N__15353\,
            I => \N__15340\
        );

    \I__3258\ : InMux
    port map (
            O => \N__15352\,
            I => \N__15340\
        );

    \I__3257\ : InMux
    port map (
            O => \N__15351\,
            I => \N__15335\
        );

    \I__3256\ : InMux
    port map (
            O => \N__15350\,
            I => \N__15335\
        );

    \I__3255\ : InMux
    port map (
            O => \N__15349\,
            I => \N__15330\
        );

    \I__3254\ : InMux
    port map (
            O => \N__15348\,
            I => \N__15323\
        );

    \I__3253\ : InMux
    port map (
            O => \N__15347\,
            I => \N__15323\
        );

    \I__3252\ : InMux
    port map (
            O => \N__15346\,
            I => \N__15318\
        );

    \I__3251\ : InMux
    port map (
            O => \N__15345\,
            I => \N__15315\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__15340\,
            I => \N__15311\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__15335\,
            I => \N__15308\
        );

    \I__3248\ : InMux
    port map (
            O => \N__15334\,
            I => \N__15305\
        );

    \I__3247\ : CascadeMux
    port map (
            O => \N__15333\,
            I => \N__15302\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__15330\,
            I => \N__15294\
        );

    \I__3245\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15289\
        );

    \I__3244\ : InMux
    port map (
            O => \N__15328\,
            I => \N__15289\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__15323\,
            I => \N__15286\
        );

    \I__3242\ : InMux
    port map (
            O => \N__15322\,
            I => \N__15283\
        );

    \I__3241\ : InMux
    port map (
            O => \N__15321\,
            I => \N__15280\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__15318\,
            I => \N__15275\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__15315\,
            I => \N__15275\
        );

    \I__3238\ : InMux
    port map (
            O => \N__15314\,
            I => \N__15272\
        );

    \I__3237\ : Span4Mux_h
    port map (
            O => \N__15311\,
            I => \N__15269\
        );

    \I__3236\ : Span4Mux_h
    port map (
            O => \N__15308\,
            I => \N__15264\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__15305\,
            I => \N__15264\
        );

    \I__3234\ : InMux
    port map (
            O => \N__15302\,
            I => \N__15255\
        );

    \I__3233\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15255\
        );

    \I__3232\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15255\
        );

    \I__3231\ : InMux
    port map (
            O => \N__15299\,
            I => \N__15255\
        );

    \I__3230\ : InMux
    port map (
            O => \N__15298\,
            I => \N__15250\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15297\,
            I => \N__15250\
        );

    \I__3228\ : Span4Mux_v
    port map (
            O => \N__15294\,
            I => \N__15241\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__15289\,
            I => \N__15241\
        );

    \I__3226\ : Span4Mux_v
    port map (
            O => \N__15286\,
            I => \N__15241\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__15283\,
            I => \N__15241\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__15280\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_0\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__15275\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_0\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__15272\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_0\
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__15269\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_0\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__15264\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_0\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__15255\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_0\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__15250\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_0\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__15241\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_0\
        );

    \I__3216\ : CascadeMux
    port map (
            O => \N__15224\,
            I => \this_vga_signals.g0_1_N_5L7_x0_cascade_\
        );

    \I__3215\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15218\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__15218\,
            I => \this_vga_signals.g0_1_N_5L7_x1\
        );

    \I__3213\ : InMux
    port map (
            O => \N__15215\,
            I => \N__15211\
        );

    \I__3212\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15208\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__15211\,
            I => \N__15201\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__15208\,
            I => \N__15197\
        );

    \I__3209\ : InMux
    port map (
            O => \N__15207\,
            I => \N__15192\
        );

    \I__3208\ : InMux
    port map (
            O => \N__15206\,
            I => \N__15192\
        );

    \I__3207\ : InMux
    port map (
            O => \N__15205\,
            I => \N__15180\
        );

    \I__3206\ : InMux
    port map (
            O => \N__15204\,
            I => \N__15180\
        );

    \I__3205\ : Span4Mux_h
    port map (
            O => \N__15201\,
            I => \N__15176\
        );

    \I__3204\ : InMux
    port map (
            O => \N__15200\,
            I => \N__15173\
        );

    \I__3203\ : Span4Mux_h
    port map (
            O => \N__15197\,
            I => \N__15170\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__15192\,
            I => \N__15167\
        );

    \I__3201\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15164\
        );

    \I__3200\ : InMux
    port map (
            O => \N__15190\,
            I => \N__15159\
        );

    \I__3199\ : InMux
    port map (
            O => \N__15189\,
            I => \N__15159\
        );

    \I__3198\ : InMux
    port map (
            O => \N__15188\,
            I => \N__15150\
        );

    \I__3197\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15150\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15186\,
            I => \N__15150\
        );

    \I__3195\ : InMux
    port map (
            O => \N__15185\,
            I => \N__15150\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__15180\,
            I => \N__15147\
        );

    \I__3193\ : InMux
    port map (
            O => \N__15179\,
            I => \N__15144\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__15176\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__15173\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3\
        );

    \I__3190\ : Odrv4
    port map (
            O => \N__15170\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__15167\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__15164\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__15159\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__15150\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3\
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__15147\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__15144\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3\
        );

    \I__3183\ : CascadeMux
    port map (
            O => \N__15125\,
            I => \N__15114\
        );

    \I__3182\ : InMux
    port map (
            O => \N__15124\,
            I => \N__15106\
        );

    \I__3181\ : InMux
    port map (
            O => \N__15123\,
            I => \N__15106\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__15122\,
            I => \N__15102\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__15121\,
            I => \N__15097\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__15120\,
            I => \N__15094\
        );

    \I__3177\ : CascadeMux
    port map (
            O => \N__15119\,
            I => \N__15086\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__15118\,
            I => \N__15079\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15117\,
            I => \N__15074\
        );

    \I__3174\ : InMux
    port map (
            O => \N__15114\,
            I => \N__15074\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__15113\,
            I => \N__15071\
        );

    \I__3172\ : InMux
    port map (
            O => \N__15112\,
            I => \N__15068\
        );

    \I__3171\ : InMux
    port map (
            O => \N__15111\,
            I => \N__15065\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__15106\,
            I => \N__15061\
        );

    \I__3169\ : InMux
    port map (
            O => \N__15105\,
            I => \N__15058\
        );

    \I__3168\ : InMux
    port map (
            O => \N__15102\,
            I => \N__15055\
        );

    \I__3167\ : InMux
    port map (
            O => \N__15101\,
            I => \N__15050\
        );

    \I__3166\ : InMux
    port map (
            O => \N__15100\,
            I => \N__15050\
        );

    \I__3165\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15047\
        );

    \I__3164\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15041\
        );

    \I__3163\ : InMux
    port map (
            O => \N__15093\,
            I => \N__15038\
        );

    \I__3162\ : InMux
    port map (
            O => \N__15092\,
            I => \N__15033\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15091\,
            I => \N__15033\
        );

    \I__3160\ : InMux
    port map (
            O => \N__15090\,
            I => \N__15026\
        );

    \I__3159\ : InMux
    port map (
            O => \N__15089\,
            I => \N__15026\
        );

    \I__3158\ : InMux
    port map (
            O => \N__15086\,
            I => \N__15026\
        );

    \I__3157\ : InMux
    port map (
            O => \N__15085\,
            I => \N__15019\
        );

    \I__3156\ : InMux
    port map (
            O => \N__15084\,
            I => \N__15019\
        );

    \I__3155\ : InMux
    port map (
            O => \N__15083\,
            I => \N__15019\
        );

    \I__3154\ : InMux
    port map (
            O => \N__15082\,
            I => \N__15014\
        );

    \I__3153\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15014\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__15074\,
            I => \N__15011\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15071\,
            I => \N__15008\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__15068\,
            I => \N__15005\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__15065\,
            I => \N__15002\
        );

    \I__3148\ : InMux
    port map (
            O => \N__15064\,
            I => \N__14996\
        );

    \I__3147\ : Span4Mux_v
    port map (
            O => \N__15061\,
            I => \N__14991\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__15058\,
            I => \N__14991\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__15055\,
            I => \N__14984\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__15050\,
            I => \N__14984\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__15047\,
            I => \N__14984\
        );

    \I__3142\ : InMux
    port map (
            O => \N__15046\,
            I => \N__14977\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15045\,
            I => \N__14977\
        );

    \I__3140\ : InMux
    port map (
            O => \N__15044\,
            I => \N__14977\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__15041\,
            I => \N__14964\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__15038\,
            I => \N__14964\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__15033\,
            I => \N__14964\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__15026\,
            I => \N__14964\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__15019\,
            I => \N__14964\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__15014\,
            I => \N__14964\
        );

    \I__3133\ : Span4Mux_v
    port map (
            O => \N__15011\,
            I => \N__14961\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__15008\,
            I => \N__14958\
        );

    \I__3131\ : Span4Mux_v
    port map (
            O => \N__15005\,
            I => \N__14953\
        );

    \I__3130\ : Span4Mux_v
    port map (
            O => \N__15002\,
            I => \N__14953\
        );

    \I__3129\ : InMux
    port map (
            O => \N__15001\,
            I => \N__14950\
        );

    \I__3128\ : InMux
    port map (
            O => \N__15000\,
            I => \N__14947\
        );

    \I__3127\ : InMux
    port map (
            O => \N__14999\,
            I => \N__14944\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__14996\,
            I => \N__14941\
        );

    \I__3125\ : Span4Mux_h
    port map (
            O => \N__14991\,
            I => \N__14936\
        );

    \I__3124\ : Span4Mux_v
    port map (
            O => \N__14984\,
            I => \N__14936\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__14977\,
            I => \N__14931\
        );

    \I__3122\ : Span4Mux_v
    port map (
            O => \N__14964\,
            I => \N__14931\
        );

    \I__3121\ : Span4Mux_h
    port map (
            O => \N__14961\,
            I => \N__14920\
        );

    \I__3120\ : Span4Mux_h
    port map (
            O => \N__14958\,
            I => \N__14920\
        );

    \I__3119\ : Span4Mux_h
    port map (
            O => \N__14953\,
            I => \N__14920\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__14950\,
            I => \N__14920\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__14947\,
            I => \N__14920\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__14944\,
            I => \this_vga_signals.M_vaddress_qZ0Z_4\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__14941\,
            I => \this_vga_signals.M_vaddress_qZ0Z_4\
        );

    \I__3114\ : Odrv4
    port map (
            O => \N__14936\,
            I => \this_vga_signals.M_vaddress_qZ0Z_4\
        );

    \I__3113\ : Odrv4
    port map (
            O => \N__14931\,
            I => \this_vga_signals.M_vaddress_qZ0Z_4\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__14920\,
            I => \this_vga_signals.M_vaddress_qZ0Z_4\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__14909\,
            I => \this_vga_signals.g0_1_N_5L7_ns_cascade_\
        );

    \I__3110\ : InMux
    port map (
            O => \N__14906\,
            I => \N__14903\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__14903\,
            I => \N__14900\
        );

    \I__3108\ : Span4Mux_h
    port map (
            O => \N__14900\,
            I => \N__14897\
        );

    \I__3107\ : Odrv4
    port map (
            O => \N__14897\,
            I => \this_vga_signals.g0_1_1_0\
        );

    \I__3106\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14890\
        );

    \I__3105\ : InMux
    port map (
            O => \N__14893\,
            I => \N__14887\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__14890\,
            I => \this_vga_signals.N_355_0\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__14887\,
            I => \this_vga_signals.N_355_0\
        );

    \I__3102\ : InMux
    port map (
            O => \N__14882\,
            I => \N__14879\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__14879\,
            I => \this_vga_signals.g1_4\
        );

    \I__3100\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14867\
        );

    \I__3099\ : InMux
    port map (
            O => \N__14875\,
            I => \N__14862\
        );

    \I__3098\ : InMux
    port map (
            O => \N__14874\,
            I => \N__14862\
        );

    \I__3097\ : InMux
    port map (
            O => \N__14873\,
            I => \N__14857\
        );

    \I__3096\ : InMux
    port map (
            O => \N__14872\,
            I => \N__14857\
        );

    \I__3095\ : InMux
    port map (
            O => \N__14871\,
            I => \N__14854\
        );

    \I__3094\ : InMux
    port map (
            O => \N__14870\,
            I => \N__14851\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__14867\,
            I => \N__14846\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__14862\,
            I => \N__14846\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__14857\,
            I => \N__14843\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__14854\,
            I => \N__14840\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__14851\,
            I => \this_vga_signals.M_vaddress_qZ0Z_7\
        );

    \I__3088\ : Odrv4
    port map (
            O => \N__14846\,
            I => \this_vga_signals.M_vaddress_qZ0Z_7\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__14843\,
            I => \this_vga_signals.M_vaddress_qZ0Z_7\
        );

    \I__3086\ : Odrv12
    port map (
            O => \N__14840\,
            I => \this_vga_signals.M_vaddress_qZ0Z_7\
        );

    \I__3085\ : InMux
    port map (
            O => \N__14831\,
            I => \N__14819\
        );

    \I__3084\ : InMux
    port map (
            O => \N__14830\,
            I => \N__14816\
        );

    \I__3083\ : InMux
    port map (
            O => \N__14829\,
            I => \N__14813\
        );

    \I__3082\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14810\
        );

    \I__3081\ : InMux
    port map (
            O => \N__14827\,
            I => \N__14801\
        );

    \I__3080\ : InMux
    port map (
            O => \N__14826\,
            I => \N__14801\
        );

    \I__3079\ : InMux
    port map (
            O => \N__14825\,
            I => \N__14801\
        );

    \I__3078\ : InMux
    port map (
            O => \N__14824\,
            I => \N__14801\
        );

    \I__3077\ : InMux
    port map (
            O => \N__14823\,
            I => \N__14797\
        );

    \I__3076\ : InMux
    port map (
            O => \N__14822\,
            I => \N__14794\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__14819\,
            I => \N__14791\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__14816\,
            I => \N__14782\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__14813\,
            I => \N__14782\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__14810\,
            I => \N__14782\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__14801\,
            I => \N__14782\
        );

    \I__3070\ : InMux
    port map (
            O => \N__14800\,
            I => \N__14779\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__14797\,
            I => \this_vga_signals.M_vaddress_qZ0Z_8\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__14794\,
            I => \this_vga_signals.M_vaddress_qZ0Z_8\
        );

    \I__3067\ : Odrv4
    port map (
            O => \N__14791\,
            I => \this_vga_signals.M_vaddress_qZ0Z_8\
        );

    \I__3066\ : Odrv4
    port map (
            O => \N__14782\,
            I => \this_vga_signals.M_vaddress_qZ0Z_8\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__14779\,
            I => \this_vga_signals.M_vaddress_qZ0Z_8\
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__14768\,
            I => \N__14762\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__14767\,
            I => \N__14759\
        );

    \I__3062\ : InMux
    port map (
            O => \N__14766\,
            I => \N__14750\
        );

    \I__3061\ : InMux
    port map (
            O => \N__14765\,
            I => \N__14746\
        );

    \I__3060\ : InMux
    port map (
            O => \N__14762\,
            I => \N__14743\
        );

    \I__3059\ : InMux
    port map (
            O => \N__14759\,
            I => \N__14738\
        );

    \I__3058\ : InMux
    port map (
            O => \N__14758\,
            I => \N__14738\
        );

    \I__3057\ : InMux
    port map (
            O => \N__14757\,
            I => \N__14735\
        );

    \I__3056\ : CascadeMux
    port map (
            O => \N__14756\,
            I => \N__14732\
        );

    \I__3055\ : CascadeMux
    port map (
            O => \N__14755\,
            I => \N__14729\
        );

    \I__3054\ : InMux
    port map (
            O => \N__14754\,
            I => \N__14724\
        );

    \I__3053\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14724\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__14750\,
            I => \N__14720\
        );

    \I__3051\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14717\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__14746\,
            I => \N__14708\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__14743\,
            I => \N__14708\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__14738\,
            I => \N__14708\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__14735\,
            I => \N__14708\
        );

    \I__3046\ : InMux
    port map (
            O => \N__14732\,
            I => \N__14702\
        );

    \I__3045\ : InMux
    port map (
            O => \N__14729\,
            I => \N__14702\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__14724\,
            I => \N__14699\
        );

    \I__3043\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14696\
        );

    \I__3042\ : Span4Mux_v
    port map (
            O => \N__14720\,
            I => \N__14689\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__14717\,
            I => \N__14689\
        );

    \I__3040\ : Span4Mux_v
    port map (
            O => \N__14708\,
            I => \N__14689\
        );

    \I__3039\ : InMux
    port map (
            O => \N__14707\,
            I => \N__14686\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__14702\,
            I => \N__14683\
        );

    \I__3037\ : Odrv4
    port map (
            O => \N__14699\,
            I => \this_vga_signals.M_vaddress_qZ0Z_6\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__14696\,
            I => \this_vga_signals.M_vaddress_qZ0Z_6\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__14689\,
            I => \this_vga_signals.M_vaddress_qZ0Z_6\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__14686\,
            I => \this_vga_signals.M_vaddress_qZ0Z_6\
        );

    \I__3033\ : Odrv4
    port map (
            O => \N__14683\,
            I => \this_vga_signals.M_vaddress_qZ0Z_6\
        );

    \I__3032\ : InMux
    port map (
            O => \N__14672\,
            I => \N__14661\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__14671\,
            I => \N__14657\
        );

    \I__3030\ : InMux
    port map (
            O => \N__14670\,
            I => \N__14653\
        );

    \I__3029\ : InMux
    port map (
            O => \N__14669\,
            I => \N__14650\
        );

    \I__3028\ : InMux
    port map (
            O => \N__14668\,
            I => \N__14645\
        );

    \I__3027\ : InMux
    port map (
            O => \N__14667\,
            I => \N__14645\
        );

    \I__3026\ : InMux
    port map (
            O => \N__14666\,
            I => \N__14640\
        );

    \I__3025\ : InMux
    port map (
            O => \N__14665\,
            I => \N__14640\
        );

    \I__3024\ : InMux
    port map (
            O => \N__14664\,
            I => \N__14637\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__14661\,
            I => \N__14634\
        );

    \I__3022\ : InMux
    port map (
            O => \N__14660\,
            I => \N__14629\
        );

    \I__3021\ : InMux
    port map (
            O => \N__14657\,
            I => \N__14629\
        );

    \I__3020\ : InMux
    port map (
            O => \N__14656\,
            I => \N__14626\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__14653\,
            I => \this_vga_signals.CO0\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__14650\,
            I => \this_vga_signals.CO0\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__14645\,
            I => \this_vga_signals.CO0\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__14640\,
            I => \this_vga_signals.CO0\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__14637\,
            I => \this_vga_signals.CO0\
        );

    \I__3014\ : Odrv4
    port map (
            O => \N__14634\,
            I => \this_vga_signals.CO0\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__14629\,
            I => \this_vga_signals.CO0\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__14626\,
            I => \this_vga_signals.CO0\
        );

    \I__3011\ : InMux
    port map (
            O => \N__14609\,
            I => \N__14606\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__14606\,
            I => \N__14603\
        );

    \I__3009\ : Span4Mux_h
    port map (
            O => \N__14603\,
            I => \N__14600\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__14600\,
            I => \this_vga_signals.if_i2_mux\
        );

    \I__3007\ : InMux
    port map (
            O => \N__14597\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_4\
        );

    \I__3006\ : InMux
    port map (
            O => \N__14594\,
            I => \N__14587\
        );

    \I__3005\ : InMux
    port map (
            O => \N__14593\,
            I => \N__14587\
        );

    \I__3004\ : InMux
    port map (
            O => \N__14592\,
            I => \N__14584\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__14587\,
            I => \N__14581\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__14584\,
            I => \N__14578\
        );

    \I__3001\ : Span4Mux_h
    port map (
            O => \N__14581\,
            I => \N__14575\
        );

    \I__3000\ : Odrv4
    port map (
            O => \N__14578\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNEZ0\
        );

    \I__2999\ : Odrv4
    port map (
            O => \N__14575\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNEZ0\
        );

    \I__2998\ : InMux
    port map (
            O => \N__14570\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_5\
        );

    \I__2997\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14558\
        );

    \I__2996\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14558\
        );

    \I__2995\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14558\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__14558\,
            I => \N__14555\
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__14555\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_6_c_RNISQOEZ0\
        );

    \I__2992\ : InMux
    port map (
            O => \N__14552\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_6\
        );

    \I__2991\ : InMux
    port map (
            O => \N__14549\,
            I => \bfn_23_10_0_\
        );

    \I__2990\ : InMux
    port map (
            O => \N__14546\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_8\
        );

    \I__2989\ : InMux
    port map (
            O => \N__14543\,
            I => \N__14540\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__14540\,
            I => \N__14536\
        );

    \I__2987\ : InMux
    port map (
            O => \N__14539\,
            I => \N__14533\
        );

    \I__2986\ : Odrv4
    port map (
            O => \N__14536\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01REZ0\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__14533\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01REZ0\
        );

    \I__2984\ : InMux
    port map (
            O => \N__14528\,
            I => \N__14524\
        );

    \I__2983\ : InMux
    port map (
            O => \N__14527\,
            I => \N__14521\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__14524\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPEZ0\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__14521\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPEZ0\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__14516\,
            I => \N__14512\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__14515\,
            I => \N__14489\
        );

    \I__2978\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14486\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__14511\,
            I => \N__14483\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__14510\,
            I => \N__14478\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__14509\,
            I => \N__14472\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__14508\,
            I => \N__14468\
        );

    \I__2973\ : InMux
    port map (
            O => \N__14507\,
            I => \N__14465\
        );

    \I__2972\ : InMux
    port map (
            O => \N__14506\,
            I => \N__14462\
        );

    \I__2971\ : InMux
    port map (
            O => \N__14505\,
            I => \N__14459\
        );

    \I__2970\ : InMux
    port map (
            O => \N__14504\,
            I => \N__14454\
        );

    \I__2969\ : InMux
    port map (
            O => \N__14503\,
            I => \N__14454\
        );

    \I__2968\ : InMux
    port map (
            O => \N__14502\,
            I => \N__14449\
        );

    \I__2967\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14449\
        );

    \I__2966\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14445\
        );

    \I__2965\ : InMux
    port map (
            O => \N__14499\,
            I => \N__14442\
        );

    \I__2964\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14437\
        );

    \I__2963\ : InMux
    port map (
            O => \N__14497\,
            I => \N__14437\
        );

    \I__2962\ : InMux
    port map (
            O => \N__14496\,
            I => \N__14427\
        );

    \I__2961\ : InMux
    port map (
            O => \N__14495\,
            I => \N__14427\
        );

    \I__2960\ : InMux
    port map (
            O => \N__14494\,
            I => \N__14427\
        );

    \I__2959\ : InMux
    port map (
            O => \N__14493\,
            I => \N__14427\
        );

    \I__2958\ : InMux
    port map (
            O => \N__14492\,
            I => \N__14422\
        );

    \I__2957\ : InMux
    port map (
            O => \N__14489\,
            I => \N__14422\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__14486\,
            I => \N__14419\
        );

    \I__2955\ : InMux
    port map (
            O => \N__14483\,
            I => \N__14416\
        );

    \I__2954\ : InMux
    port map (
            O => \N__14482\,
            I => \N__14413\
        );

    \I__2953\ : InMux
    port map (
            O => \N__14481\,
            I => \N__14406\
        );

    \I__2952\ : InMux
    port map (
            O => \N__14478\,
            I => \N__14406\
        );

    \I__2951\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14406\
        );

    \I__2950\ : InMux
    port map (
            O => \N__14476\,
            I => \N__14403\
        );

    \I__2949\ : InMux
    port map (
            O => \N__14475\,
            I => \N__14400\
        );

    \I__2948\ : InMux
    port map (
            O => \N__14472\,
            I => \N__14397\
        );

    \I__2947\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14394\
        );

    \I__2946\ : InMux
    port map (
            O => \N__14468\,
            I => \N__14391\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__14465\,
            I => \N__14388\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__14462\,
            I => \N__14385\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__14459\,
            I => \N__14382\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__14454\,
            I => \N__14377\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__14449\,
            I => \N__14377\
        );

    \I__2940\ : InMux
    port map (
            O => \N__14448\,
            I => \N__14374\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__14445\,
            I => \N__14367\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__14442\,
            I => \N__14367\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__14437\,
            I => \N__14367\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__14436\,
            I => \N__14364\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__14427\,
            I => \N__14351\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__14422\,
            I => \N__14351\
        );

    \I__2933\ : Span4Mux_h
    port map (
            O => \N__14419\,
            I => \N__14351\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__14416\,
            I => \N__14351\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__14413\,
            I => \N__14351\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__14406\,
            I => \N__14351\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__14403\,
            I => \N__14340\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__14400\,
            I => \N__14340\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__14397\,
            I => \N__14340\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__14394\,
            I => \N__14340\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__14391\,
            I => \N__14340\
        );

    \I__2924\ : Span4Mux_v
    port map (
            O => \N__14388\,
            I => \N__14336\
        );

    \I__2923\ : Span4Mux_v
    port map (
            O => \N__14385\,
            I => \N__14329\
        );

    \I__2922\ : Span4Mux_v
    port map (
            O => \N__14382\,
            I => \N__14329\
        );

    \I__2921\ : Span4Mux_h
    port map (
            O => \N__14377\,
            I => \N__14329\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__14374\,
            I => \N__14324\
        );

    \I__2919\ : Span4Mux_v
    port map (
            O => \N__14367\,
            I => \N__14324\
        );

    \I__2918\ : InMux
    port map (
            O => \N__14364\,
            I => \N__14321\
        );

    \I__2917\ : Span4Mux_v
    port map (
            O => \N__14351\,
            I => \N__14316\
        );

    \I__2916\ : Span4Mux_v
    port map (
            O => \N__14340\,
            I => \N__14316\
        );

    \I__2915\ : InMux
    port map (
            O => \N__14339\,
            I => \N__14313\
        );

    \I__2914\ : Span4Mux_h
    port map (
            O => \N__14336\,
            I => \N__14310\
        );

    \I__2913\ : Span4Mux_h
    port map (
            O => \N__14329\,
            I => \N__14307\
        );

    \I__2912\ : Span4Mux_h
    port map (
            O => \N__14324\,
            I => \N__14302\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__14321\,
            I => \N__14302\
        );

    \I__2910\ : Span4Mux_h
    port map (
            O => \N__14316\,
            I => \N__14299\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__14313\,
            I => \this_vga_signals.M_vaddress_qZ0Z_3\
        );

    \I__2908\ : Odrv4
    port map (
            O => \N__14310\,
            I => \this_vga_signals.M_vaddress_qZ0Z_3\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__14307\,
            I => \this_vga_signals.M_vaddress_qZ0Z_3\
        );

    \I__2906\ : Odrv4
    port map (
            O => \N__14302\,
            I => \this_vga_signals.M_vaddress_qZ0Z_3\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__14299\,
            I => \this_vga_signals.M_vaddress_qZ0Z_3\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__14288\,
            I => \this_vga_signals.N_1253_0_cascade_\
        );

    \I__2903\ : CEMux
    port map (
            O => \N__14285\,
            I => \N__14282\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__14282\,
            I => \N__14278\
        );

    \I__2901\ : CEMux
    port map (
            O => \N__14281\,
            I => \N__14275\
        );

    \I__2900\ : Span4Mux_v
    port map (
            O => \N__14278\,
            I => \N__14270\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__14275\,
            I => \N__14270\
        );

    \I__2898\ : Span4Mux_v
    port map (
            O => \N__14270\,
            I => \N__14267\
        );

    \I__2897\ : Span4Mux_v
    port map (
            O => \N__14267\,
            I => \N__14264\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__14264\,
            I => \this_vram.mem_WE_2\
        );

    \I__2895\ : InMux
    port map (
            O => \N__14261\,
            I => \N__14258\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__14258\,
            I => \N__14255\
        );

    \I__2893\ : Span12Mux_h
    port map (
            O => \N__14255\,
            I => \N__14252\
        );

    \I__2892\ : Odrv12
    port map (
            O => \N__14252\,
            I => port_address_c_5
        );

    \I__2891\ : InMux
    port map (
            O => \N__14249\,
            I => \N__14246\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__14246\,
            I => \N__14243\
        );

    \I__2889\ : Span12Mux_v
    port map (
            O => \N__14243\,
            I => \N__14240\
        );

    \I__2888\ : Odrv12
    port map (
            O => \N__14240\,
            I => port_address_c_2
        );

    \I__2887\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14234\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__14234\,
            I => \N__14231\
        );

    \I__2885\ : Span4Mux_v
    port map (
            O => \N__14231\,
            I => \N__14228\
        );

    \I__2884\ : Sp12to4
    port map (
            O => \N__14228\,
            I => \N__14225\
        );

    \I__2883\ : Odrv12
    port map (
            O => \N__14225\,
            I => port_address_c_6
        );

    \I__2882\ : InMux
    port map (
            O => \N__14222\,
            I => \N__14219\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__14219\,
            I => \N__14216\
        );

    \I__2880\ : Span4Mux_v
    port map (
            O => \N__14216\,
            I => \N__14213\
        );

    \I__2879\ : Odrv4
    port map (
            O => \N__14213\,
            I => \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_3Z0Z_0\
        );

    \I__2878\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14207\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__14207\,
            I => \N__14203\
        );

    \I__2876\ : InMux
    port map (
            O => \N__14206\,
            I => \N__14200\
        );

    \I__2875\ : Span4Mux_h
    port map (
            O => \N__14203\,
            I => \N__14196\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__14200\,
            I => \N__14193\
        );

    \I__2873\ : InMux
    port map (
            O => \N__14199\,
            I => \N__14190\
        );

    \I__2872\ : Span4Mux_v
    port map (
            O => \N__14196\,
            I => \N__14184\
        );

    \I__2871\ : Span4Mux_h
    port map (
            O => \N__14193\,
            I => \N__14184\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__14190\,
            I => \N__14181\
        );

    \I__2869\ : InMux
    port map (
            O => \N__14189\,
            I => \N__14178\
        );

    \I__2868\ : Span4Mux_v
    port map (
            O => \N__14184\,
            I => \N__14172\
        );

    \I__2867\ : Span4Mux_h
    port map (
            O => \N__14181\,
            I => \N__14172\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__14178\,
            I => \N__14169\
        );

    \I__2865\ : InMux
    port map (
            O => \N__14177\,
            I => \N__14166\
        );

    \I__2864\ : Span4Mux_v
    port map (
            O => \N__14172\,
            I => \N__14160\
        );

    \I__2863\ : Span4Mux_h
    port map (
            O => \N__14169\,
            I => \N__14160\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__14166\,
            I => \N__14157\
        );

    \I__2861\ : InMux
    port map (
            O => \N__14165\,
            I => \N__14154\
        );

    \I__2860\ : Span4Mux_v
    port map (
            O => \N__14160\,
            I => \N__14147\
        );

    \I__2859\ : Span4Mux_h
    port map (
            O => \N__14157\,
            I => \N__14147\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__14154\,
            I => \N__14144\
        );

    \I__2857\ : InMux
    port map (
            O => \N__14153\,
            I => \N__14141\
        );

    \I__2856\ : InMux
    port map (
            O => \N__14152\,
            I => \N__14138\
        );

    \I__2855\ : Span4Mux_v
    port map (
            O => \N__14147\,
            I => \N__14133\
        );

    \I__2854\ : Span4Mux_h
    port map (
            O => \N__14144\,
            I => \N__14133\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__14141\,
            I => \N__14130\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__14138\,
            I => \N__14127\
        );

    \I__2851\ : Span4Mux_v
    port map (
            O => \N__14133\,
            I => \N__14119\
        );

    \I__2850\ : Span4Mux_h
    port map (
            O => \N__14130\,
            I => \N__14119\
        );

    \I__2849\ : Span4Mux_h
    port map (
            O => \N__14127\,
            I => \N__14119\
        );

    \I__2848\ : InMux
    port map (
            O => \N__14126\,
            I => \N__14116\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__14119\,
            I => \M_current_data_qZ0Z_1\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__14116\,
            I => \M_current_data_qZ0Z_1\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__14111\,
            I => \N__14107\
        );

    \I__2844\ : InMux
    port map (
            O => \N__14110\,
            I => \N__14104\
        );

    \I__2843\ : InMux
    port map (
            O => \N__14107\,
            I => \N__14101\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__14104\,
            I => \N__14094\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__14101\,
            I => \N__14094\
        );

    \I__2840\ : InMux
    port map (
            O => \N__14100\,
            I => \N__14089\
        );

    \I__2839\ : InMux
    port map (
            O => \N__14099\,
            I => \N__14086\
        );

    \I__2838\ : Span4Mux_h
    port map (
            O => \N__14094\,
            I => \N__14083\
        );

    \I__2837\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14077\
        );

    \I__2836\ : InMux
    port map (
            O => \N__14092\,
            I => \N__14077\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__14089\,
            I => \N__14072\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__14086\,
            I => \N__14072\
        );

    \I__2833\ : Span4Mux_v
    port map (
            O => \N__14083\,
            I => \N__14069\
        );

    \I__2832\ : InMux
    port map (
            O => \N__14082\,
            I => \N__14066\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__14077\,
            I => \N__14063\
        );

    \I__2830\ : Span4Mux_h
    port map (
            O => \N__14072\,
            I => \N__14058\
        );

    \I__2829\ : Span4Mux_h
    port map (
            O => \N__14069\,
            I => \N__14058\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__14066\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__14063\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa\
        );

    \I__2826\ : Odrv4
    port map (
            O => \N__14058\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa\
        );

    \I__2825\ : InMux
    port map (
            O => \N__14051\,
            I => \N__14047\
        );

    \I__2824\ : InMux
    port map (
            O => \N__14050\,
            I => \N__14044\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__14047\,
            I => \N__14041\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__14044\,
            I => \this_vga_signals.M_vaddress_qZ0Z_0\
        );

    \I__2821\ : Odrv4
    port map (
            O => \N__14041\,
            I => \this_vga_signals.M_vaddress_qZ0Z_0\
        );

    \I__2820\ : InMux
    port map (
            O => \N__14036\,
            I => \N__14033\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__14033\,
            I => \N__14024\
        );

    \I__2818\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14021\
        );

    \I__2817\ : InMux
    port map (
            O => \N__14031\,
            I => \N__14017\
        );

    \I__2816\ : InMux
    port map (
            O => \N__14030\,
            I => \N__14010\
        );

    \I__2815\ : InMux
    port map (
            O => \N__14029\,
            I => \N__14010\
        );

    \I__2814\ : InMux
    port map (
            O => \N__14028\,
            I => \N__14010\
        );

    \I__2813\ : InMux
    port map (
            O => \N__14027\,
            I => \N__14007\
        );

    \I__2812\ : Span4Mux_v
    port map (
            O => \N__14024\,
            I => \N__14004\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__14021\,
            I => \N__14001\
        );

    \I__2810\ : InMux
    port map (
            O => \N__14020\,
            I => \N__13998\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__14017\,
            I => \N__13991\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__14010\,
            I => \N__13991\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__14007\,
            I => \N__13991\
        );

    \I__2806\ : Span4Mux_h
    port map (
            O => \N__14004\,
            I => \N__13986\
        );

    \I__2805\ : Span4Mux_h
    port map (
            O => \N__14001\,
            I => \N__13986\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__13998\,
            I => \this_vga_signals.M_vaddress_qZ0Z_1\
        );

    \I__2803\ : Odrv12
    port map (
            O => \N__13991\,
            I => \this_vga_signals.M_vaddress_qZ0Z_1\
        );

    \I__2802\ : Odrv4
    port map (
            O => \N__13986\,
            I => \this_vga_signals.M_vaddress_qZ0Z_1\
        );

    \I__2801\ : InMux
    port map (
            O => \N__13979\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_0\
        );

    \I__2800\ : CascadeMux
    port map (
            O => \N__13976\,
            I => \N__13969\
        );

    \I__2799\ : InMux
    port map (
            O => \N__13975\,
            I => \N__13966\
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__13974\,
            I => \N__13955\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__13973\,
            I => \N__13952\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__13972\,
            I => \N__13949\
        );

    \I__2795\ : InMux
    port map (
            O => \N__13969\,
            I => \N__13945\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__13966\,
            I => \N__13941\
        );

    \I__2793\ : InMux
    port map (
            O => \N__13965\,
            I => \N__13936\
        );

    \I__2792\ : InMux
    port map (
            O => \N__13964\,
            I => \N__13936\
        );

    \I__2791\ : InMux
    port map (
            O => \N__13963\,
            I => \N__13933\
        );

    \I__2790\ : InMux
    port map (
            O => \N__13962\,
            I => \N__13929\
        );

    \I__2789\ : InMux
    port map (
            O => \N__13961\,
            I => \N__13926\
        );

    \I__2788\ : InMux
    port map (
            O => \N__13960\,
            I => \N__13915\
        );

    \I__2787\ : InMux
    port map (
            O => \N__13959\,
            I => \N__13915\
        );

    \I__2786\ : InMux
    port map (
            O => \N__13958\,
            I => \N__13915\
        );

    \I__2785\ : InMux
    port map (
            O => \N__13955\,
            I => \N__13915\
        );

    \I__2784\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13915\
        );

    \I__2783\ : InMux
    port map (
            O => \N__13949\,
            I => \N__13910\
        );

    \I__2782\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13910\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__13945\,
            I => \N__13907\
        );

    \I__2780\ : InMux
    port map (
            O => \N__13944\,
            I => \N__13904\
        );

    \I__2779\ : Span4Mux_v
    port map (
            O => \N__13941\,
            I => \N__13901\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__13936\,
            I => \N__13896\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__13933\,
            I => \N__13896\
        );

    \I__2776\ : InMux
    port map (
            O => \N__13932\,
            I => \N__13891\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__13929\,
            I => \N__13882\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__13926\,
            I => \N__13882\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__13915\,
            I => \N__13882\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__13910\,
            I => \N__13882\
        );

    \I__2771\ : Span12Mux_h
    port map (
            O => \N__13907\,
            I => \N__13879\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__13904\,
            I => \N__13871\
        );

    \I__2769\ : Span4Mux_h
    port map (
            O => \N__13901\,
            I => \N__13871\
        );

    \I__2768\ : Span4Mux_v
    port map (
            O => \N__13896\,
            I => \N__13871\
        );

    \I__2767\ : InMux
    port map (
            O => \N__13895\,
            I => \N__13866\
        );

    \I__2766\ : InMux
    port map (
            O => \N__13894\,
            I => \N__13866\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__13891\,
            I => \N__13861\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__13882\,
            I => \N__13861\
        );

    \I__2763\ : Span12Mux_v
    port map (
            O => \N__13879\,
            I => \N__13858\
        );

    \I__2762\ : InMux
    port map (
            O => \N__13878\,
            I => \N__13855\
        );

    \I__2761\ : Sp12to4
    port map (
            O => \N__13871\,
            I => \N__13850\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__13866\,
            I => \N__13850\
        );

    \I__2759\ : Span4Mux_h
    port map (
            O => \N__13861\,
            I => \N__13847\
        );

    \I__2758\ : Odrv12
    port map (
            O => \N__13858\,
            I => \this_vga_signals.M_vaddress_qZ0Z_2\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__13855\,
            I => \this_vga_signals.M_vaddress_qZ0Z_2\
        );

    \I__2756\ : Odrv12
    port map (
            O => \N__13850\,
            I => \this_vga_signals.M_vaddress_qZ0Z_2\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__13847\,
            I => \this_vga_signals.M_vaddress_qZ0Z_2\
        );

    \I__2754\ : InMux
    port map (
            O => \N__13838\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_1\
        );

    \I__2753\ : InMux
    port map (
            O => \N__13835\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_2\
        );

    \I__2752\ : InMux
    port map (
            O => \N__13832\,
            I => \this_vga_signals.un1_M_vaddress_q_cry_3\
        );

    \I__2751\ : CascadeMux
    port map (
            O => \N__13829\,
            I => \N__13825\
        );

    \I__2750\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13820\
        );

    \I__2749\ : InMux
    port map (
            O => \N__13825\,
            I => \N__13820\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__13820\,
            I => \this_vga_signals.N_9_0\
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__13817\,
            I => \N__13812\
        );

    \I__2746\ : InMux
    port map (
            O => \N__13816\,
            I => \N__13806\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__13815\,
            I => \N__13801\
        );

    \I__2744\ : InMux
    port map (
            O => \N__13812\,
            I => \N__13798\
        );

    \I__2743\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13795\
        );

    \I__2742\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13792\
        );

    \I__2741\ : InMux
    port map (
            O => \N__13809\,
            I => \N__13789\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__13806\,
            I => \N__13786\
        );

    \I__2739\ : InMux
    port map (
            O => \N__13805\,
            I => \N__13783\
        );

    \I__2738\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13778\
        );

    \I__2737\ : InMux
    port map (
            O => \N__13801\,
            I => \N__13778\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__13798\,
            I => \this_vga_signals.M_vaddress_q_6_repZ0Z1\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__13795\,
            I => \this_vga_signals.M_vaddress_q_6_repZ0Z1\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__13792\,
            I => \this_vga_signals.M_vaddress_q_6_repZ0Z1\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__13789\,
            I => \this_vga_signals.M_vaddress_q_6_repZ0Z1\
        );

    \I__2732\ : Odrv4
    port map (
            O => \N__13786\,
            I => \this_vga_signals.M_vaddress_q_6_repZ0Z1\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__13783\,
            I => \this_vga_signals.M_vaddress_q_6_repZ0Z1\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__13778\,
            I => \this_vga_signals.M_vaddress_q_6_repZ0Z1\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__13763\,
            I => \N__13756\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__13762\,
            I => \N__13753\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__13761\,
            I => \N__13749\
        );

    \I__2726\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13744\
        );

    \I__2725\ : InMux
    port map (
            O => \N__13759\,
            I => \N__13741\
        );

    \I__2724\ : InMux
    port map (
            O => \N__13756\,
            I => \N__13734\
        );

    \I__2723\ : InMux
    port map (
            O => \N__13753\,
            I => \N__13734\
        );

    \I__2722\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13734\
        );

    \I__2721\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13731\
        );

    \I__2720\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13728\
        );

    \I__2719\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13725\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__13744\,
            I => \N__13720\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__13741\,
            I => \N__13720\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__13734\,
            I => \N__13717\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__13731\,
            I => \this_vga_signals.M_vaddress_q_7_repZ0Z1\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__13728\,
            I => \this_vga_signals.M_vaddress_q_7_repZ0Z1\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__13725\,
            I => \this_vga_signals.M_vaddress_q_7_repZ0Z1\
        );

    \I__2712\ : Odrv12
    port map (
            O => \N__13720\,
            I => \this_vga_signals.M_vaddress_q_7_repZ0Z1\
        );

    \I__2711\ : Odrv4
    port map (
            O => \N__13717\,
            I => \this_vga_signals.M_vaddress_q_7_repZ0Z1\
        );

    \I__2710\ : InMux
    port map (
            O => \N__13706\,
            I => \N__13696\
        );

    \I__2709\ : InMux
    port map (
            O => \N__13705\,
            I => \N__13696\
        );

    \I__2708\ : InMux
    port map (
            O => \N__13704\,
            I => \N__13696\
        );

    \I__2707\ : InMux
    port map (
            O => \N__13703\,
            I => \N__13693\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__13696\,
            I => \N__13688\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__13693\,
            I => \N__13688\
        );

    \I__2704\ : Odrv4
    port map (
            O => \N__13688\,
            I => \this_vga_signals.N_15_0\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__13685\,
            I => \this_vga_signals.N_15_0_0_cascade_\
        );

    \I__2702\ : InMux
    port map (
            O => \N__13682\,
            I => \N__13679\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__13679\,
            I => \N__13674\
        );

    \I__2700\ : InMux
    port map (
            O => \N__13678\,
            I => \N__13670\
        );

    \I__2699\ : InMux
    port map (
            O => \N__13677\,
            I => \N__13666\
        );

    \I__2698\ : Span4Mux_h
    port map (
            O => \N__13674\,
            I => \N__13663\
        );

    \I__2697\ : InMux
    port map (
            O => \N__13673\,
            I => \N__13660\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__13670\,
            I => \N__13648\
        );

    \I__2695\ : InMux
    port map (
            O => \N__13669\,
            I => \N__13645\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__13666\,
            I => \N__13640\
        );

    \I__2693\ : Span4Mux_v
    port map (
            O => \N__13663\,
            I => \N__13640\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__13660\,
            I => \N__13637\
        );

    \I__2691\ : InMux
    port map (
            O => \N__13659\,
            I => \N__13628\
        );

    \I__2690\ : InMux
    port map (
            O => \N__13658\,
            I => \N__13628\
        );

    \I__2689\ : InMux
    port map (
            O => \N__13657\,
            I => \N__13628\
        );

    \I__2688\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13628\
        );

    \I__2687\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13617\
        );

    \I__2686\ : InMux
    port map (
            O => \N__13654\,
            I => \N__13617\
        );

    \I__2685\ : InMux
    port map (
            O => \N__13653\,
            I => \N__13617\
        );

    \I__2684\ : InMux
    port map (
            O => \N__13652\,
            I => \N__13617\
        );

    \I__2683\ : InMux
    port map (
            O => \N__13651\,
            I => \N__13617\
        );

    \I__2682\ : Odrv12
    port map (
            O => \N__13648\,
            I => \this_vga_signals.M_haddress_qZ0Z_9\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__13645\,
            I => \this_vga_signals.M_haddress_qZ0Z_9\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__13640\,
            I => \this_vga_signals.M_haddress_qZ0Z_9\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__13637\,
            I => \this_vga_signals.M_haddress_qZ0Z_9\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__13628\,
            I => \this_vga_signals.M_haddress_qZ0Z_9\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__13617\,
            I => \this_vga_signals.M_haddress_qZ0Z_9\
        );

    \I__2676\ : InMux
    port map (
            O => \N__13604\,
            I => \N__13601\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__13601\,
            I => \N__13596\
        );

    \I__2674\ : InMux
    port map (
            O => \N__13600\,
            I => \N__13592\
        );

    \I__2673\ : InMux
    port map (
            O => \N__13599\,
            I => \N__13588\
        );

    \I__2672\ : Span4Mux_h
    port map (
            O => \N__13596\,
            I => \N__13585\
        );

    \I__2671\ : InMux
    port map (
            O => \N__13595\,
            I => \N__13582\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__13592\,
            I => \N__13570\
        );

    \I__2669\ : InMux
    port map (
            O => \N__13591\,
            I => \N__13567\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__13588\,
            I => \N__13562\
        );

    \I__2667\ : Span4Mux_v
    port map (
            O => \N__13585\,
            I => \N__13562\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__13582\,
            I => \N__13559\
        );

    \I__2665\ : InMux
    port map (
            O => \N__13581\,
            I => \N__13552\
        );

    \I__2664\ : InMux
    port map (
            O => \N__13580\,
            I => \N__13552\
        );

    \I__2663\ : InMux
    port map (
            O => \N__13579\,
            I => \N__13552\
        );

    \I__2662\ : InMux
    port map (
            O => \N__13578\,
            I => \N__13547\
        );

    \I__2661\ : InMux
    port map (
            O => \N__13577\,
            I => \N__13547\
        );

    \I__2660\ : InMux
    port map (
            O => \N__13576\,
            I => \N__13542\
        );

    \I__2659\ : InMux
    port map (
            O => \N__13575\,
            I => \N__13542\
        );

    \I__2658\ : InMux
    port map (
            O => \N__13574\,
            I => \N__13537\
        );

    \I__2657\ : InMux
    port map (
            O => \N__13573\,
            I => \N__13537\
        );

    \I__2656\ : Odrv12
    port map (
            O => \N__13570\,
            I => \this_vga_signals.M_haddress_qZ0Z_8\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__13567\,
            I => \this_vga_signals.M_haddress_qZ0Z_8\
        );

    \I__2654\ : Odrv4
    port map (
            O => \N__13562\,
            I => \this_vga_signals.M_haddress_qZ0Z_8\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__13559\,
            I => \this_vga_signals.M_haddress_qZ0Z_8\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__13552\,
            I => \this_vga_signals.M_haddress_qZ0Z_8\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__13547\,
            I => \this_vga_signals.M_haddress_qZ0Z_8\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__13542\,
            I => \this_vga_signals.M_haddress_qZ0Z_8\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__13537\,
            I => \this_vga_signals.M_haddress_qZ0Z_8\
        );

    \I__2648\ : CascadeMux
    port map (
            O => \N__13520\,
            I => \N__13517\
        );

    \I__2647\ : InMux
    port map (
            O => \N__13517\,
            I => \N__13511\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__13516\,
            I => \N__13508\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__13515\,
            I => \N__13504\
        );

    \I__2644\ : CascadeMux
    port map (
            O => \N__13514\,
            I => \N__13498\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__13511\,
            I => \N__13494\
        );

    \I__2642\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13490\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__13507\,
            I => \N__13487\
        );

    \I__2640\ : InMux
    port map (
            O => \N__13504\,
            I => \N__13484\
        );

    \I__2639\ : CascadeMux
    port map (
            O => \N__13503\,
            I => \N__13480\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__13502\,
            I => \N__13477\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__13501\,
            I => \N__13472\
        );

    \I__2636\ : InMux
    port map (
            O => \N__13498\,
            I => \N__13465\
        );

    \I__2635\ : InMux
    port map (
            O => \N__13497\,
            I => \N__13465\
        );

    \I__2634\ : Span4Mux_h
    port map (
            O => \N__13494\,
            I => \N__13462\
        );

    \I__2633\ : InMux
    port map (
            O => \N__13493\,
            I => \N__13459\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__13490\,
            I => \N__13456\
        );

    \I__2631\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13453\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__13484\,
            I => \N__13450\
        );

    \I__2629\ : InMux
    port map (
            O => \N__13483\,
            I => \N__13445\
        );

    \I__2628\ : InMux
    port map (
            O => \N__13480\,
            I => \N__13445\
        );

    \I__2627\ : InMux
    port map (
            O => \N__13477\,
            I => \N__13436\
        );

    \I__2626\ : InMux
    port map (
            O => \N__13476\,
            I => \N__13436\
        );

    \I__2625\ : InMux
    port map (
            O => \N__13475\,
            I => \N__13436\
        );

    \I__2624\ : InMux
    port map (
            O => \N__13472\,
            I => \N__13436\
        );

    \I__2623\ : InMux
    port map (
            O => \N__13471\,
            I => \N__13431\
        );

    \I__2622\ : InMux
    port map (
            O => \N__13470\,
            I => \N__13431\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__13465\,
            I => \N__13426\
        );

    \I__2620\ : Span4Mux_v
    port map (
            O => \N__13462\,
            I => \N__13426\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__13459\,
            I => \this_vga_signals.M_haddress_qZ0Z_10\
        );

    \I__2618\ : Odrv12
    port map (
            O => \N__13456\,
            I => \this_vga_signals.M_haddress_qZ0Z_10\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__13453\,
            I => \this_vga_signals.M_haddress_qZ0Z_10\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__13450\,
            I => \this_vga_signals.M_haddress_qZ0Z_10\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__13445\,
            I => \this_vga_signals.M_haddress_qZ0Z_10\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__13436\,
            I => \this_vga_signals.M_haddress_qZ0Z_10\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__13431\,
            I => \this_vga_signals.M_haddress_qZ0Z_10\
        );

    \I__2612\ : Odrv4
    port map (
            O => \N__13426\,
            I => \this_vga_signals.M_haddress_qZ0Z_10\
        );

    \I__2611\ : InMux
    port map (
            O => \N__13409\,
            I => \N__13406\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__13406\,
            I => \N__13399\
        );

    \I__2609\ : InMux
    port map (
            O => \N__13405\,
            I => \N__13395\
        );

    \I__2608\ : InMux
    port map (
            O => \N__13404\,
            I => \N__13392\
        );

    \I__2607\ : InMux
    port map (
            O => \N__13403\,
            I => \N__13387\
        );

    \I__2606\ : InMux
    port map (
            O => \N__13402\,
            I => \N__13387\
        );

    \I__2605\ : Span4Mux_v
    port map (
            O => \N__13399\,
            I => \N__13376\
        );

    \I__2604\ : InMux
    port map (
            O => \N__13398\,
            I => \N__13373\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__13395\,
            I => \N__13370\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__13392\,
            I => \N__13365\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__13387\,
            I => \N__13365\
        );

    \I__2600\ : InMux
    port map (
            O => \N__13386\,
            I => \N__13354\
        );

    \I__2599\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13354\
        );

    \I__2598\ : InMux
    port map (
            O => \N__13384\,
            I => \N__13354\
        );

    \I__2597\ : InMux
    port map (
            O => \N__13383\,
            I => \N__13354\
        );

    \I__2596\ : InMux
    port map (
            O => \N__13382\,
            I => \N__13354\
        );

    \I__2595\ : InMux
    port map (
            O => \N__13381\,
            I => \N__13347\
        );

    \I__2594\ : InMux
    port map (
            O => \N__13380\,
            I => \N__13347\
        );

    \I__2593\ : InMux
    port map (
            O => \N__13379\,
            I => \N__13347\
        );

    \I__2592\ : Span4Mux_h
    port map (
            O => \N__13376\,
            I => \N__13344\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__13373\,
            I => \this_vga_signals.CO0_0\
        );

    \I__2590\ : Odrv12
    port map (
            O => \N__13370\,
            I => \this_vga_signals.CO0_0\
        );

    \I__2589\ : Odrv4
    port map (
            O => \N__13365\,
            I => \this_vga_signals.CO0_0\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__13354\,
            I => \this_vga_signals.CO0_0\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__13347\,
            I => \this_vga_signals.CO0_0\
        );

    \I__2586\ : Odrv4
    port map (
            O => \N__13344\,
            I => \this_vga_signals.CO0_0\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__13331\,
            I => \N__13328\
        );

    \I__2584\ : CascadeBuf
    port map (
            O => \N__13328\,
            I => \N__13325\
        );

    \I__2583\ : CascadeMux
    port map (
            O => \N__13325\,
            I => \N__13322\
        );

    \I__2582\ : CascadeBuf
    port map (
            O => \N__13322\,
            I => \N__13319\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__13319\,
            I => \N__13316\
        );

    \I__2580\ : CascadeBuf
    port map (
            O => \N__13316\,
            I => \N__13313\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__13313\,
            I => \N__13310\
        );

    \I__2578\ : CascadeBuf
    port map (
            O => \N__13310\,
            I => \N__13307\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__13307\,
            I => \N__13304\
        );

    \I__2576\ : CascadeBuf
    port map (
            O => \N__13304\,
            I => \N__13301\
        );

    \I__2575\ : CascadeMux
    port map (
            O => \N__13301\,
            I => \N__13298\
        );

    \I__2574\ : CascadeBuf
    port map (
            O => \N__13298\,
            I => \N__13295\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__13295\,
            I => \N__13292\
        );

    \I__2572\ : CascadeBuf
    port map (
            O => \N__13292\,
            I => \N__13289\
        );

    \I__2571\ : CascadeMux
    port map (
            O => \N__13289\,
            I => \N__13286\
        );

    \I__2570\ : CascadeBuf
    port map (
            O => \N__13286\,
            I => \N__13283\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__13283\,
            I => \N__13280\
        );

    \I__2568\ : CascadeBuf
    port map (
            O => \N__13280\,
            I => \N__13277\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__13277\,
            I => \N__13274\
        );

    \I__2566\ : CascadeBuf
    port map (
            O => \N__13274\,
            I => \N__13271\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__13271\,
            I => \N__13268\
        );

    \I__2564\ : CascadeBuf
    port map (
            O => \N__13268\,
            I => \N__13265\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__13265\,
            I => \N__13262\
        );

    \I__2562\ : CascadeBuf
    port map (
            O => \N__13262\,
            I => \N__13259\
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__13259\,
            I => \N__13256\
        );

    \I__2560\ : CascadeBuf
    port map (
            O => \N__13256\,
            I => \N__13253\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__13253\,
            I => \N__13250\
        );

    \I__2558\ : CascadeBuf
    port map (
            O => \N__13250\,
            I => \N__13247\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__13247\,
            I => \N__13244\
        );

    \I__2556\ : CascadeBuf
    port map (
            O => \N__13244\,
            I => \N__13241\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__13241\,
            I => \N__13238\
        );

    \I__2554\ : InMux
    port map (
            O => \N__13238\,
            I => \N__13235\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__13235\,
            I => \N__13232\
        );

    \I__2552\ : Span4Mux_v
    port map (
            O => \N__13232\,
            I => \N__13229\
        );

    \I__2551\ : Span4Mux_v
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__2550\ : Span4Mux_v
    port map (
            O => \N__13226\,
            I => \N__13223\
        );

    \I__2549\ : Span4Mux_v
    port map (
            O => \N__13223\,
            I => \N__13220\
        );

    \I__2548\ : Odrv4
    port map (
            O => \N__13220\,
            I => \M_haddress_q_RNI8ARU_11\
        );

    \I__2547\ : InMux
    port map (
            O => \N__13217\,
            I => \N__13214\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__13214\,
            I => \N__13210\
        );

    \I__2545\ : InMux
    port map (
            O => \N__13213\,
            I => \N__13205\
        );

    \I__2544\ : Span4Mux_h
    port map (
            O => \N__13210\,
            I => \N__13202\
        );

    \I__2543\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13199\
        );

    \I__2542\ : InMux
    port map (
            O => \N__13208\,
            I => \N__13196\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__13205\,
            I => \M_state_qZ0Z_1\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__13202\,
            I => \M_state_qZ0Z_1\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__13199\,
            I => \M_state_qZ0Z_1\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__13196\,
            I => \M_state_qZ0Z_1\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__13187\,
            I => \N__13181\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__13186\,
            I => \N__13177\
        );

    \I__2535\ : InMux
    port map (
            O => \N__13185\,
            I => \N__13174\
        );

    \I__2534\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13169\
        );

    \I__2533\ : InMux
    port map (
            O => \N__13181\,
            I => \N__13169\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__13180\,
            I => \N__13162\
        );

    \I__2531\ : InMux
    port map (
            O => \N__13177\,
            I => \N__13159\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__13174\,
            I => \N__13154\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__13169\,
            I => \N__13154\
        );

    \I__2528\ : InMux
    port map (
            O => \N__13168\,
            I => \N__13149\
        );

    \I__2527\ : InMux
    port map (
            O => \N__13167\,
            I => \N__13149\
        );

    \I__2526\ : InMux
    port map (
            O => \N__13166\,
            I => \N__13146\
        );

    \I__2525\ : InMux
    port map (
            O => \N__13165\,
            I => \N__13143\
        );

    \I__2524\ : InMux
    port map (
            O => \N__13162\,
            I => \N__13140\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__13159\,
            I => \N__13137\
        );

    \I__2522\ : Span4Mux_v
    port map (
            O => \N__13154\,
            I => \N__13134\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__13149\,
            I => \N__13129\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__13146\,
            I => \N__13129\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__13143\,
            I => \N__13124\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__13140\,
            I => \N__13124\
        );

    \I__2517\ : Span4Mux_v
    port map (
            O => \N__13137\,
            I => \N__13121\
        );

    \I__2516\ : Span4Mux_h
    port map (
            O => \N__13134\,
            I => \N__13118\
        );

    \I__2515\ : Span4Mux_v
    port map (
            O => \N__13129\,
            I => \N__13115\
        );

    \I__2514\ : Span12Mux_v
    port map (
            O => \N__13124\,
            I => \N__13110\
        );

    \I__2513\ : Sp12to4
    port map (
            O => \N__13121\,
            I => \N__13110\
        );

    \I__2512\ : Sp12to4
    port map (
            O => \N__13118\,
            I => \N__13105\
        );

    \I__2511\ : Sp12to4
    port map (
            O => \N__13115\,
            I => \N__13105\
        );

    \I__2510\ : Span12Mux_h
    port map (
            O => \N__13110\,
            I => \N__13102\
        );

    \I__2509\ : Span12Mux_h
    port map (
            O => \N__13105\,
            I => \N__13099\
        );

    \I__2508\ : Odrv12
    port map (
            O => \N__13102\,
            I => port_enb_c
        );

    \I__2507\ : Odrv12
    port map (
            O => \N__13099\,
            I => port_enb_c
        );

    \I__2506\ : InMux
    port map (
            O => \N__13094\,
            I => \N__13088\
        );

    \I__2505\ : InMux
    port map (
            O => \N__13093\,
            I => \N__13085\
        );

    \I__2504\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13082\
        );

    \I__2503\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13079\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__13088\,
            I => \N__13074\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__13085\,
            I => \N__13074\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__13082\,
            I => \M_state_qZ0Z_3\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__13079\,
            I => \M_state_qZ0Z_3\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__13074\,
            I => \M_state_qZ0Z_3\
        );

    \I__2497\ : InMux
    port map (
            O => \N__13067\,
            I => \N__13059\
        );

    \I__2496\ : InMux
    port map (
            O => \N__13066\,
            I => \N__13056\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13065\,
            I => \N__13053\
        );

    \I__2494\ : InMux
    port map (
            O => \N__13064\,
            I => \N__13047\
        );

    \I__2493\ : InMux
    port map (
            O => \N__13063\,
            I => \N__13047\
        );

    \I__2492\ : InMux
    port map (
            O => \N__13062\,
            I => \N__13042\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__13059\,
            I => \N__13039\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__13056\,
            I => \N__13034\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__13053\,
            I => \N__13034\
        );

    \I__2488\ : InMux
    port map (
            O => \N__13052\,
            I => \N__13031\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__13047\,
            I => \N__13028\
        );

    \I__2486\ : InMux
    port map (
            O => \N__13046\,
            I => \N__13023\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13045\,
            I => \N__13023\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__13042\,
            I => \N__13018\
        );

    \I__2483\ : Span4Mux_h
    port map (
            O => \N__13039\,
            I => \N__13018\
        );

    \I__2482\ : Span4Mux_h
    port map (
            O => \N__13034\,
            I => \N__13015\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__13031\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__13028\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__13023\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__2478\ : Odrv4
    port map (
            O => \N__13018\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__13015\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__2476\ : InMux
    port map (
            O => \N__13004\,
            I => \N__12998\
        );

    \I__2475\ : InMux
    port map (
            O => \N__13003\,
            I => \N__12998\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__12998\,
            I => \this_vga_signals.M_vaddress_q_fastZ0Z_5\
        );

    \I__2473\ : InMux
    port map (
            O => \N__12995\,
            I => \N__12991\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__12994\,
            I => \N__12985\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__12991\,
            I => \N__12982\
        );

    \I__2470\ : InMux
    port map (
            O => \N__12990\,
            I => \N__12975\
        );

    \I__2469\ : InMux
    port map (
            O => \N__12989\,
            I => \N__12975\
        );

    \I__2468\ : InMux
    port map (
            O => \N__12988\,
            I => \N__12975\
        );

    \I__2467\ : InMux
    port map (
            O => \N__12985\,
            I => \N__12972\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__12982\,
            I => \this_vga_signals.M_vaddress_q_fastZ0Z_9\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__12975\,
            I => \this_vga_signals.M_vaddress_q_fastZ0Z_9\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__12972\,
            I => \this_vga_signals.M_vaddress_q_fastZ0Z_9\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__12965\,
            I => \N__12958\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__12964\,
            I => \N__12955\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__12963\,
            I => \N__12952\
        );

    \I__2460\ : InMux
    port map (
            O => \N__12962\,
            I => \N__12949\
        );

    \I__2459\ : InMux
    port map (
            O => \N__12961\,
            I => \N__12940\
        );

    \I__2458\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12940\
        );

    \I__2457\ : InMux
    port map (
            O => \N__12955\,
            I => \N__12940\
        );

    \I__2456\ : InMux
    port map (
            O => \N__12952\,
            I => \N__12940\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__12949\,
            I => \this_vga_signals.M_vaddress_q_fastZ0Z_8\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__12940\,
            I => \this_vga_signals.M_vaddress_q_fastZ0Z_8\
        );

    \I__2453\ : InMux
    port map (
            O => \N__12935\,
            I => \N__12931\
        );

    \I__2452\ : InMux
    port map (
            O => \N__12934\,
            I => \N__12928\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__12931\,
            I => \this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__12928\,
            I => \this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8\
        );

    \I__2449\ : CascadeMux
    port map (
            O => \N__12923\,
            I => \this_vga_signals.N_353_0_cascade_\
        );

    \I__2448\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12912\
        );

    \I__2447\ : InMux
    port map (
            O => \N__12919\,
            I => \N__12912\
        );

    \I__2446\ : InMux
    port map (
            O => \N__12918\,
            I => \N__12907\
        );

    \I__2445\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12907\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__12912\,
            I => \this_vga_signals.mult1_un40_sum_m_bm_2\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__12907\,
            I => \this_vga_signals.mult1_un40_sum_m_bm_2\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__12902\,
            I => \this_vga_signals.mult1_un40_sum_0_axbxc3_5_1_0_cascade_\
        );

    \I__2441\ : InMux
    port map (
            O => \N__12899\,
            I => \N__12896\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__12896\,
            I => \this_vga_signals.mult1_un40_sum_0_axbxc3_5_3\
        );

    \I__2439\ : InMux
    port map (
            O => \N__12893\,
            I => \N__12887\
        );

    \I__2438\ : InMux
    port map (
            O => \N__12892\,
            I => \N__12887\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__12887\,
            I => \N__12883\
        );

    \I__2436\ : InMux
    port map (
            O => \N__12886\,
            I => \N__12878\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__12883\,
            I => \N__12875\
        );

    \I__2434\ : InMux
    port map (
            O => \N__12882\,
            I => \N__12870\
        );

    \I__2433\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12870\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__12878\,
            I => \this_vga_signals.mult1_un40_sum0_3\
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__12875\,
            I => \this_vga_signals.mult1_un40_sum0_3\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__12870\,
            I => \this_vga_signals.mult1_un40_sum0_3\
        );

    \I__2429\ : InMux
    port map (
            O => \N__12863\,
            I => \N__12852\
        );

    \I__2428\ : InMux
    port map (
            O => \N__12862\,
            I => \N__12852\
        );

    \I__2427\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12845\
        );

    \I__2426\ : InMux
    port map (
            O => \N__12860\,
            I => \N__12845\
        );

    \I__2425\ : InMux
    port map (
            O => \N__12859\,
            I => \N__12845\
        );

    \I__2424\ : InMux
    port map (
            O => \N__12858\,
            I => \N__12840\
        );

    \I__2423\ : InMux
    port map (
            O => \N__12857\,
            I => \N__12840\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__12852\,
            I => \this_vga_signals.M_vaddress_q_5_repZ0Z1\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__12845\,
            I => \this_vga_signals.M_vaddress_q_5_repZ0Z1\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__12840\,
            I => \this_vga_signals.M_vaddress_q_5_repZ0Z1\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__12833\,
            I => \N__12830\
        );

    \I__2418\ : InMux
    port map (
            O => \N__12830\,
            I => \N__12827\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__12827\,
            I => \N__12824\
        );

    \I__2416\ : Span4Mux_v
    port map (
            O => \N__12824\,
            I => \N__12821\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__12821\,
            I => \this_vga_signals.mult1_un40_sum_0_axb1\
        );

    \I__2414\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12815\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__12815\,
            I => \this_vga_signals.mult1_un40_sum_m_1_1\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__12812\,
            I => \this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8_cascade_\
        );

    \I__2411\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12805\
        );

    \I__2410\ : CascadeMux
    port map (
            O => \N__12808\,
            I => \N__12801\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__12805\,
            I => \N__12798\
        );

    \I__2408\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12795\
        );

    \I__2407\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12792\
        );

    \I__2406\ : Span4Mux_v
    port map (
            O => \N__12798\,
            I => \N__12787\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__12795\,
            I => \N__12787\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__12792\,
            I => \this_vga_signals.mult1_un40_sum_m_0_1\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__12787\,
            I => \this_vga_signals.mult1_un40_sum_m_0_1\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__12782\,
            I => \N__12779\
        );

    \I__2401\ : InMux
    port map (
            O => \N__12779\,
            I => \N__12775\
        );

    \I__2400\ : InMux
    port map (
            O => \N__12778\,
            I => \N__12772\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__12775\,
            I => \this_vga_signals.M_vaddress_q_fastZ0Z_6\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__12772\,
            I => \this_vga_signals.M_vaddress_q_fastZ0Z_6\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__12767\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_2_0_cascade_\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__12764\,
            I => \N__12760\
        );

    \I__2395\ : InMux
    port map (
            O => \N__12763\,
            I => \N__12757\
        );

    \I__2394\ : InMux
    port map (
            O => \N__12760\,
            I => \N__12754\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__12757\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_2\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__12754\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_2\
        );

    \I__2391\ : CascadeMux
    port map (
            O => \N__12749\,
            I => \N__12746\
        );

    \I__2390\ : InMux
    port map (
            O => \N__12746\,
            I => \N__12743\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__12743\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc3_a4_1_0\
        );

    \I__2388\ : InMux
    port map (
            O => \N__12740\,
            I => \N__12734\
        );

    \I__2387\ : InMux
    port map (
            O => \N__12739\,
            I => \N__12731\
        );

    \I__2386\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12726\
        );

    \I__2385\ : InMux
    port map (
            O => \N__12737\,
            I => \N__12726\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__12734\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__12731\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__12726\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0\
        );

    \I__2381\ : InMux
    port map (
            O => \N__12719\,
            I => \N__12714\
        );

    \I__2380\ : InMux
    port map (
            O => \N__12718\,
            I => \N__12711\
        );

    \I__2379\ : InMux
    port map (
            O => \N__12717\,
            I => \N__12708\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__12714\,
            I => \this_vga_signals.if_m5_0_s\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__12711\,
            I => \this_vga_signals.if_m5_0_s\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__12708\,
            I => \this_vga_signals.if_m5_0_s\
        );

    \I__2375\ : InMux
    port map (
            O => \N__12701\,
            I => \N__12696\
        );

    \I__2374\ : InMux
    port map (
            O => \N__12700\,
            I => \N__12693\
        );

    \I__2373\ : InMux
    port map (
            O => \N__12699\,
            I => \N__12690\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__12696\,
            I => \this_vga_signals.if_m1_0\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__12693\,
            I => \this_vga_signals.if_m1_0\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__12690\,
            I => \this_vga_signals.if_m1_0\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__12683\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\
        );

    \I__2368\ : CascadeMux
    port map (
            O => \N__12680\,
            I => \this_vga_signals.if_N_2_2_cascade_\
        );

    \I__2367\ : InMux
    port map (
            O => \N__12677\,
            I => \N__12674\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__12674\,
            I => \N__12670\
        );

    \I__2365\ : InMux
    port map (
            O => \N__12673\,
            I => \N__12667\
        );

    \I__2364\ : Span4Mux_v
    port map (
            O => \N__12670\,
            I => \N__12664\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__12667\,
            I => \this_vga_signals.mult1_un54_sum_axb1_3\
        );

    \I__2362\ : Odrv4
    port map (
            O => \N__12664\,
            I => \this_vga_signals.mult1_un54_sum_axb1_3\
        );

    \I__2361\ : InMux
    port map (
            O => \N__12659\,
            I => \N__12656\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__12656\,
            I => \N__12653\
        );

    \I__2359\ : Span4Mux_h
    port map (
            O => \N__12653\,
            I => \N__12650\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__12650\,
            I => \this_vga_signals.mult1_un61_sum_c3_1_0\
        );

    \I__2357\ : InMux
    port map (
            O => \N__12647\,
            I => \N__12642\
        );

    \I__2356\ : InMux
    port map (
            O => \N__12646\,
            I => \N__12637\
        );

    \I__2355\ : InMux
    port map (
            O => \N__12645\,
            I => \N__12637\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__12642\,
            I => \M_state_qZ0Z_2\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__12637\,
            I => \M_state_qZ0Z_2\
        );

    \I__2352\ : InMux
    port map (
            O => \N__12632\,
            I => \N__12624\
        );

    \I__2351\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12615\
        );

    \I__2350\ : InMux
    port map (
            O => \N__12630\,
            I => \N__12615\
        );

    \I__2349\ : InMux
    port map (
            O => \N__12629\,
            I => \N__12612\
        );

    \I__2348\ : InMux
    port map (
            O => \N__12628\,
            I => \N__12609\
        );

    \I__2347\ : InMux
    port map (
            O => \N__12627\,
            I => \N__12602\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__12624\,
            I => \N__12599\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__12623\,
            I => \N__12595\
        );

    \I__2344\ : InMux
    port map (
            O => \N__12622\,
            I => \N__12588\
        );

    \I__2343\ : InMux
    port map (
            O => \N__12621\,
            I => \N__12588\
        );

    \I__2342\ : InMux
    port map (
            O => \N__12620\,
            I => \N__12581\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__12615\,
            I => \N__12576\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__12612\,
            I => \N__12576\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__12609\,
            I => \N__12573\
        );

    \I__2338\ : InMux
    port map (
            O => \N__12608\,
            I => \N__12568\
        );

    \I__2337\ : InMux
    port map (
            O => \N__12607\,
            I => \N__12568\
        );

    \I__2336\ : InMux
    port map (
            O => \N__12606\,
            I => \N__12565\
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__12605\,
            I => \N__12560\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__12602\,
            I => \N__12549\
        );

    \I__2333\ : Span12Mux_h
    port map (
            O => \N__12599\,
            I => \N__12549\
        );

    \I__2332\ : InMux
    port map (
            O => \N__12598\,
            I => \N__12546\
        );

    \I__2331\ : InMux
    port map (
            O => \N__12595\,
            I => \N__12541\
        );

    \I__2330\ : InMux
    port map (
            O => \N__12594\,
            I => \N__12541\
        );

    \I__2329\ : InMux
    port map (
            O => \N__12593\,
            I => \N__12538\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__12588\,
            I => \N__12535\
        );

    \I__2327\ : InMux
    port map (
            O => \N__12587\,
            I => \N__12526\
        );

    \I__2326\ : InMux
    port map (
            O => \N__12586\,
            I => \N__12526\
        );

    \I__2325\ : InMux
    port map (
            O => \N__12585\,
            I => \N__12526\
        );

    \I__2324\ : InMux
    port map (
            O => \N__12584\,
            I => \N__12526\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__12581\,
            I => \N__12519\
        );

    \I__2322\ : Span4Mux_v
    port map (
            O => \N__12576\,
            I => \N__12519\
        );

    \I__2321\ : Span4Mux_v
    port map (
            O => \N__12573\,
            I => \N__12519\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__12568\,
            I => \N__12514\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__12565\,
            I => \N__12514\
        );

    \I__2318\ : InMux
    port map (
            O => \N__12564\,
            I => \N__12509\
        );

    \I__2317\ : InMux
    port map (
            O => \N__12563\,
            I => \N__12509\
        );

    \I__2316\ : InMux
    port map (
            O => \N__12560\,
            I => \N__12502\
        );

    \I__2315\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12502\
        );

    \I__2314\ : InMux
    port map (
            O => \N__12558\,
            I => \N__12502\
        );

    \I__2313\ : InMux
    port map (
            O => \N__12557\,
            I => \N__12495\
        );

    \I__2312\ : InMux
    port map (
            O => \N__12556\,
            I => \N__12495\
        );

    \I__2311\ : InMux
    port map (
            O => \N__12555\,
            I => \N__12495\
        );

    \I__2310\ : InMux
    port map (
            O => \N__12554\,
            I => \N__12492\
        );

    \I__2309\ : Odrv12
    port map (
            O => \N__12549\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__12546\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__12541\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__12538\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2305\ : Odrv4
    port map (
            O => \N__12535\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__12526\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2303\ : Odrv4
    port map (
            O => \N__12519\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__12514\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__12509\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__12502\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__12495\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__12492\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2297\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12464\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__12464\,
            I => \N__12461\
        );

    \I__2295\ : Sp12to4
    port map (
            O => \N__12461\,
            I => \N__12458\
        );

    \I__2294\ : Span12Mux_v
    port map (
            O => \N__12458\,
            I => \N__12451\
        );

    \I__2293\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12446\
        );

    \I__2292\ : InMux
    port map (
            O => \N__12456\,
            I => \N__12446\
        );

    \I__2291\ : InMux
    port map (
            O => \N__12455\,
            I => \N__12443\
        );

    \I__2290\ : InMux
    port map (
            O => \N__12454\,
            I => \N__12440\
        );

    \I__2289\ : Odrv12
    port map (
            O => \N__12451\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__12446\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__12443\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__12440\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__12431\,
            I => \N__12428\
        );

    \I__2284\ : InMux
    port map (
            O => \N__12428\,
            I => \N__12424\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__12427\,
            I => \N__12421\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__12424\,
            I => \N__12417\
        );

    \I__2281\ : InMux
    port map (
            O => \N__12421\,
            I => \N__12413\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__12420\,
            I => \N__12409\
        );

    \I__2279\ : Span4Mux_v
    port map (
            O => \N__12417\,
            I => \N__12406\
        );

    \I__2278\ : InMux
    port map (
            O => \N__12416\,
            I => \N__12403\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__12413\,
            I => \N__12400\
        );

    \I__2276\ : InMux
    port map (
            O => \N__12412\,
            I => \N__12393\
        );

    \I__2275\ : InMux
    port map (
            O => \N__12409\,
            I => \N__12393\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__12406\,
            I => \N__12388\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__12403\,
            I => \N__12388\
        );

    \I__2272\ : Span4Mux_v
    port map (
            O => \N__12400\,
            I => \N__12385\
        );

    \I__2271\ : InMux
    port map (
            O => \N__12399\,
            I => \N__12380\
        );

    \I__2270\ : InMux
    port map (
            O => \N__12398\,
            I => \N__12380\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__12393\,
            I => \N__12377\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__12388\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_1\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__12385\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_1\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__12380\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_1\
        );

    \I__2265\ : Odrv4
    port map (
            O => \N__12377\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_1\
        );

    \I__2264\ : InMux
    port map (
            O => \N__12368\,
            I => \N__12364\
        );

    \I__2263\ : InMux
    port map (
            O => \N__12367\,
            I => \N__12359\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__12364\,
            I => \N__12349\
        );

    \I__2261\ : InMux
    port map (
            O => \N__12363\,
            I => \N__12343\
        );

    \I__2260\ : InMux
    port map (
            O => \N__12362\,
            I => \N__12343\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__12359\,
            I => \N__12340\
        );

    \I__2258\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12337\
        );

    \I__2257\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12332\
        );

    \I__2256\ : InMux
    port map (
            O => \N__12356\,
            I => \N__12332\
        );

    \I__2255\ : InMux
    port map (
            O => \N__12355\,
            I => \N__12329\
        );

    \I__2254\ : InMux
    port map (
            O => \N__12354\,
            I => \N__12324\
        );

    \I__2253\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12324\
        );

    \I__2252\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12319\
        );

    \I__2251\ : Span4Mux_v
    port map (
            O => \N__12349\,
            I => \N__12306\
        );

    \I__2250\ : InMux
    port map (
            O => \N__12348\,
            I => \N__12303\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__12343\,
            I => \N__12298\
        );

    \I__2248\ : Span4Mux_v
    port map (
            O => \N__12340\,
            I => \N__12298\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__12337\,
            I => \N__12295\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__12332\,
            I => \N__12292\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__12329\,
            I => \N__12279\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__12324\,
            I => \N__12279\
        );

    \I__2243\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12274\
        );

    \I__2242\ : InMux
    port map (
            O => \N__12322\,
            I => \N__12274\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__12319\,
            I => \N__12271\
        );

    \I__2240\ : InMux
    port map (
            O => \N__12318\,
            I => \N__12266\
        );

    \I__2239\ : InMux
    port map (
            O => \N__12317\,
            I => \N__12266\
        );

    \I__2238\ : InMux
    port map (
            O => \N__12316\,
            I => \N__12259\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12315\,
            I => \N__12259\
        );

    \I__2236\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12259\
        );

    \I__2235\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12256\
        );

    \I__2234\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12247\
        );

    \I__2233\ : InMux
    port map (
            O => \N__12311\,
            I => \N__12247\
        );

    \I__2232\ : InMux
    port map (
            O => \N__12310\,
            I => \N__12247\
        );

    \I__2231\ : InMux
    port map (
            O => \N__12309\,
            I => \N__12247\
        );

    \I__2230\ : Span4Mux_v
    port map (
            O => \N__12306\,
            I => \N__12236\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__12303\,
            I => \N__12236\
        );

    \I__2228\ : Span4Mux_h
    port map (
            O => \N__12298\,
            I => \N__12236\
        );

    \I__2227\ : Span4Mux_v
    port map (
            O => \N__12295\,
            I => \N__12236\
        );

    \I__2226\ : Span4Mux_v
    port map (
            O => \N__12292\,
            I => \N__12236\
        );

    \I__2225\ : InMux
    port map (
            O => \N__12291\,
            I => \N__12229\
        );

    \I__2224\ : InMux
    port map (
            O => \N__12290\,
            I => \N__12229\
        );

    \I__2223\ : InMux
    port map (
            O => \N__12289\,
            I => \N__12229\
        );

    \I__2222\ : InMux
    port map (
            O => \N__12288\,
            I => \N__12226\
        );

    \I__2221\ : InMux
    port map (
            O => \N__12287\,
            I => \N__12217\
        );

    \I__2220\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12217\
        );

    \I__2219\ : InMux
    port map (
            O => \N__12285\,
            I => \N__12217\
        );

    \I__2218\ : InMux
    port map (
            O => \N__12284\,
            I => \N__12217\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__12279\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__12274\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2215\ : Odrv4
    port map (
            O => \N__12271\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__12266\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__12259\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__12256\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__12247\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__12236\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__12229\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__12226\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__12217\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__12194\,
            I => \N__12191\
        );

    \I__2205\ : CascadeBuf
    port map (
            O => \N__12191\,
            I => \N__12188\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__12188\,
            I => \N__12185\
        );

    \I__2203\ : CascadeBuf
    port map (
            O => \N__12185\,
            I => \N__12182\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__12182\,
            I => \N__12179\
        );

    \I__2201\ : CascadeBuf
    port map (
            O => \N__12179\,
            I => \N__12176\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__12176\,
            I => \N__12173\
        );

    \I__2199\ : CascadeBuf
    port map (
            O => \N__12173\,
            I => \N__12170\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__12170\,
            I => \N__12167\
        );

    \I__2197\ : CascadeBuf
    port map (
            O => \N__12167\,
            I => \N__12164\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__12164\,
            I => \N__12161\
        );

    \I__2195\ : CascadeBuf
    port map (
            O => \N__12161\,
            I => \N__12158\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__12158\,
            I => \N__12155\
        );

    \I__2193\ : CascadeBuf
    port map (
            O => \N__12155\,
            I => \N__12152\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__12152\,
            I => \N__12149\
        );

    \I__2191\ : CascadeBuf
    port map (
            O => \N__12149\,
            I => \N__12146\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__12146\,
            I => \N__12143\
        );

    \I__2189\ : CascadeBuf
    port map (
            O => \N__12143\,
            I => \N__12140\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__12140\,
            I => \N__12137\
        );

    \I__2187\ : CascadeBuf
    port map (
            O => \N__12137\,
            I => \N__12134\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__12134\,
            I => \N__12131\
        );

    \I__2185\ : CascadeBuf
    port map (
            O => \N__12131\,
            I => \N__12128\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__12128\,
            I => \N__12125\
        );

    \I__2183\ : CascadeBuf
    port map (
            O => \N__12125\,
            I => \N__12122\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__12122\,
            I => \N__12119\
        );

    \I__2181\ : CascadeBuf
    port map (
            O => \N__12119\,
            I => \N__12116\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__12116\,
            I => \N__12113\
        );

    \I__2179\ : CascadeBuf
    port map (
            O => \N__12113\,
            I => \N__12110\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__12110\,
            I => \N__12107\
        );

    \I__2177\ : CascadeBuf
    port map (
            O => \N__12107\,
            I => \N__12104\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__12104\,
            I => \N__12101\
        );

    \I__2175\ : InMux
    port map (
            O => \N__12101\,
            I => \N__12098\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__12098\,
            I => \N__12095\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__12095\,
            I => \N__12092\
        );

    \I__2172\ : Span4Mux_h
    port map (
            O => \N__12092\,
            I => \N__12089\
        );

    \I__2171\ : Sp12to4
    port map (
            O => \N__12089\,
            I => \N__12086\
        );

    \I__2170\ : Odrv12
    port map (
            O => \N__12086\,
            I => this_vga_signals_un14_address_if_generate_plus_mult1_un54_sum_i_3
        );

    \I__2169\ : InMux
    port map (
            O => \N__12083\,
            I => \N__12079\
        );

    \I__2168\ : InMux
    port map (
            O => \N__12082\,
            I => \N__12076\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__12079\,
            I => \N__12073\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__12076\,
            I => \N__12068\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__12073\,
            I => \N__12068\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__12068\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_4\
        );

    \I__2163\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12062\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__12062\,
            I => \this_vga_signals.M_vaddress_q_fastZ0Z_7\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__12059\,
            I => \this_vga_signals.mult1_un40_sum_m_am_x_2_cascade_\
        );

    \I__2160\ : InMux
    port map (
            O => \N__12056\,
            I => \N__12052\
        );

    \I__2159\ : InMux
    port map (
            O => \N__12055\,
            I => \N__12049\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__12052\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_2\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__12049\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_2\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12044\,
            I => \N__12040\
        );

    \I__2155\ : InMux
    port map (
            O => \N__12043\,
            I => \N__12037\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__12040\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_3\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__12037\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_3\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__12032\,
            I => \this_vga_signals.mult1_un40_sum_m_x1_3_cascade_\
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__12029\,
            I => \this_vga_signals.mult1_un40_sum_m_ns_3_cascade_\
        );

    \I__2150\ : InMux
    port map (
            O => \N__12026\,
            I => \N__12023\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__12023\,
            I => \this_vga_signals.N_6_i\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__12020\,
            I => \N__12016\
        );

    \I__2147\ : InMux
    port map (
            O => \N__12019\,
            I => \N__12012\
        );

    \I__2146\ : InMux
    port map (
            O => \N__12016\,
            I => \N__12007\
        );

    \I__2145\ : InMux
    port map (
            O => \N__12015\,
            I => \N__12007\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__12012\,
            I => \N__12004\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__12007\,
            I => \this_vga_signals.mult1_un40_sum_m_am_2\
        );

    \I__2142\ : Odrv4
    port map (
            O => \N__12004\,
            I => \this_vga_signals.mult1_un40_sum_m_am_2\
        );

    \I__2141\ : InMux
    port map (
            O => \N__11999\,
            I => \N__11996\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__11996\,
            I => \N__11992\
        );

    \I__2139\ : InMux
    port map (
            O => \N__11995\,
            I => \N__11989\
        );

    \I__2138\ : Span4Mux_h
    port map (
            O => \N__11992\,
            I => \N__11986\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__11989\,
            I => \this_vga_signals.mult1_un40_sum1_3\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__11986\,
            I => \this_vga_signals.mult1_un40_sum1_3\
        );

    \I__2135\ : InMux
    port map (
            O => \N__11981\,
            I => \N__11978\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__11978\,
            I => \this_vga_signals.N_6_i_0\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__11975\,
            I => \this_vga_signals.mult1_un40_sum1_3_cascade_\
        );

    \I__2132\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11969\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__11969\,
            I => \this_vga_signals.g0_4_0\
        );

    \I__2130\ : CascadeMux
    port map (
            O => \N__11966\,
            I => \N__11963\
        );

    \I__2129\ : InMux
    port map (
            O => \N__11963\,
            I => \N__11959\
        );

    \I__2128\ : InMux
    port map (
            O => \N__11962\,
            I => \N__11955\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__11959\,
            I => \N__11952\
        );

    \I__2126\ : InMux
    port map (
            O => \N__11958\,
            I => \N__11949\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__11955\,
            I => \N__11942\
        );

    \I__2124\ : Span4Mux_h
    port map (
            O => \N__11952\,
            I => \N__11942\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__11949\,
            I => \N__11942\
        );

    \I__2122\ : Span4Mux_v
    port map (
            O => \N__11942\,
            I => \N__11936\
        );

    \I__2121\ : InMux
    port map (
            O => \N__11941\,
            I => \N__11933\
        );

    \I__2120\ : InMux
    port map (
            O => \N__11940\,
            I => \N__11930\
        );

    \I__2119\ : InMux
    port map (
            O => \N__11939\,
            I => \N__11927\
        );

    \I__2118\ : Sp12to4
    port map (
            O => \N__11936\,
            I => \N__11924\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__11933\,
            I => \N__11917\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__11930\,
            I => \N__11917\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__11927\,
            I => \N__11917\
        );

    \I__2114\ : Span12Mux_h
    port map (
            O => \N__11924\,
            I => \N__11914\
        );

    \I__2113\ : Span12Mux_v
    port map (
            O => \N__11917\,
            I => \N__11911\
        );

    \I__2112\ : Odrv12
    port map (
            O => \N__11914\,
            I => \M_this_vram_read_data_1\
        );

    \I__2111\ : Odrv12
    port map (
            O => \N__11911\,
            I => \M_this_vram_read_data_1\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__11906\,
            I => \this_vga_signals.g0_1_1_1_cascade_\
        );

    \I__2109\ : InMux
    port map (
            O => \N__11903\,
            I => \N__11900\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__11900\,
            I => \this_vga_signals.g0_3_0_0\
        );

    \I__2107\ : InMux
    port map (
            O => \N__11897\,
            I => \N__11893\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__11896\,
            I => \N__11890\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__11893\,
            I => \N__11887\
        );

    \I__2104\ : InMux
    port map (
            O => \N__11890\,
            I => \N__11884\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__11887\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_1_1\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__11884\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_1_1\
        );

    \I__2101\ : InMux
    port map (
            O => \N__11879\,
            I => \N__11876\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__11876\,
            I => \this_vga_signals.N_2_1_0\
        );

    \I__2099\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11870\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__11870\,
            I => \this_vga_signals.g0_3_2_1\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__11867\,
            I => \this_start_data_delay.this_edge_detector.N_263_cascade_\
        );

    \I__2096\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11857\
        );

    \I__2095\ : InMux
    port map (
            O => \N__11863\,
            I => \N__11857\
        );

    \I__2094\ : InMux
    port map (
            O => \N__11862\,
            I => \N__11854\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__11857\,
            I => \M_state_qZ0Z_0\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__11854\,
            I => \M_state_qZ0Z_0\
        );

    \I__2091\ : InMux
    port map (
            O => \N__11849\,
            I => \N__11843\
        );

    \I__2090\ : InMux
    port map (
            O => \N__11848\,
            I => \N__11843\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__11843\,
            I => \N__11838\
        );

    \I__2088\ : InMux
    port map (
            O => \N__11842\,
            I => \N__11833\
        );

    \I__2087\ : InMux
    port map (
            O => \N__11841\,
            I => \N__11833\
        );

    \I__2086\ : Span4Mux_h
    port map (
            O => \N__11838\,
            I => \N__11828\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__11833\,
            I => \N__11828\
        );

    \I__2084\ : Span4Mux_v
    port map (
            O => \N__11828\,
            I => \N__11825\
        );

    \I__2083\ : Span4Mux_v
    port map (
            O => \N__11825\,
            I => \N__11822\
        );

    \I__2082\ : Span4Mux_v
    port map (
            O => \N__11822\,
            I => \N__11819\
        );

    \I__2081\ : IoSpan4Mux
    port map (
            O => \N__11819\,
            I => \N__11816\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__11816\,
            I => port_address_c_0
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__11813\,
            I => \N__11808\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__11812\,
            I => \N__11804\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__11811\,
            I => \N__11801\
        );

    \I__2076\ : InMux
    port map (
            O => \N__11808\,
            I => \N__11796\
        );

    \I__2075\ : InMux
    port map (
            O => \N__11807\,
            I => \N__11796\
        );

    \I__2074\ : InMux
    port map (
            O => \N__11804\,
            I => \N__11791\
        );

    \I__2073\ : InMux
    port map (
            O => \N__11801\,
            I => \N__11791\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__11796\,
            I => \N__11788\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__11791\,
            I => \N__11785\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__11788\,
            I => \N__11782\
        );

    \I__2069\ : Span12Mux_h
    port map (
            O => \N__11785\,
            I => \N__11779\
        );

    \I__2068\ : Sp12to4
    port map (
            O => \N__11782\,
            I => \N__11776\
        );

    \I__2067\ : Span12Mux_v
    port map (
            O => \N__11779\,
            I => \N__11773\
        );

    \I__2066\ : Span12Mux_h
    port map (
            O => \N__11776\,
            I => \N__11770\
        );

    \I__2065\ : Odrv12
    port map (
            O => \N__11773\,
            I => port_address_c_1
        );

    \I__2064\ : Odrv12
    port map (
            O => \N__11770\,
            I => port_address_c_1
        );

    \I__2063\ : InMux
    port map (
            O => \N__11765\,
            I => \N__11758\
        );

    \I__2062\ : InMux
    port map (
            O => \N__11764\,
            I => \N__11758\
        );

    \I__2061\ : InMux
    port map (
            O => \N__11763\,
            I => \N__11755\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__11758\,
            I => \this_start_data_delay.this_edge_detector.N_275\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__11755\,
            I => \this_start_data_delay.this_edge_detector.N_275\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__11750\,
            I => \this_start_data_delay.this_edge_detector.N_259_cascade_\
        );

    \I__2057\ : InMux
    port map (
            O => \N__11747\,
            I => \N__11744\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__11744\,
            I => \N__11741\
        );

    \I__2055\ : Span4Mux_s2_v
    port map (
            O => \N__11741\,
            I => \N__11738\
        );

    \I__2054\ : Sp12to4
    port map (
            O => \N__11738\,
            I => \N__11735\
        );

    \I__2053\ : Span12Mux_s6_v
    port map (
            O => \N__11735\,
            I => \N__11732\
        );

    \I__2052\ : Span12Mux_v
    port map (
            O => \N__11732\,
            I => \N__11729\
        );

    \I__2051\ : Odrv12
    port map (
            O => \N__11729\,
            I => \this_vga_signals.mult1_un61_sum_axbxc1\
        );

    \I__2050\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11723\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__11723\,
            I => \N__11720\
        );

    \I__2048\ : Span12Mux_s11_v
    port map (
            O => \N__11720\,
            I => \N__11717\
        );

    \I__2047\ : Odrv12
    port map (
            O => \N__11717\,
            I => \this_vga_signals.mult1_un68_sum_i_1_3\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__11714\,
            I => \N__11711\
        );

    \I__2045\ : InMux
    port map (
            O => \N__11711\,
            I => \N__11708\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__11708\,
            I => \N__11705\
        );

    \I__2043\ : Span4Mux_v
    port map (
            O => \N__11705\,
            I => \N__11702\
        );

    \I__2042\ : Span4Mux_v
    port map (
            O => \N__11702\,
            I => \N__11695\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__11701\,
            I => \N__11691\
        );

    \I__2040\ : InMux
    port map (
            O => \N__11700\,
            I => \N__11688\
        );

    \I__2039\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11685\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__11698\,
            I => \N__11682\
        );

    \I__2037\ : Span4Mux_v
    port map (
            O => \N__11695\,
            I => \N__11679\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__11694\,
            I => \N__11674\
        );

    \I__2035\ : InMux
    port map (
            O => \N__11691\,
            I => \N__11671\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__11688\,
            I => \N__11668\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__11685\,
            I => \N__11665\
        );

    \I__2032\ : InMux
    port map (
            O => \N__11682\,
            I => \N__11662\
        );

    \I__2031\ : Span4Mux_v
    port map (
            O => \N__11679\,
            I => \N__11659\
        );

    \I__2030\ : InMux
    port map (
            O => \N__11678\,
            I => \N__11656\
        );

    \I__2029\ : InMux
    port map (
            O => \N__11677\,
            I => \N__11651\
        );

    \I__2028\ : InMux
    port map (
            O => \N__11674\,
            I => \N__11651\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__11671\,
            I => \N__11648\
        );

    \I__2026\ : Span4Mux_h
    port map (
            O => \N__11668\,
            I => \N__11641\
        );

    \I__2025\ : Span4Mux_h
    port map (
            O => \N__11665\,
            I => \N__11641\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__11662\,
            I => \N__11641\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__11659\,
            I => \this_vga_signals.M_haddress_qZ0Z_4\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__11656\,
            I => \this_vga_signals.M_haddress_qZ0Z_4\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__11651\,
            I => \this_vga_signals.M_haddress_qZ0Z_4\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__11648\,
            I => \this_vga_signals.M_haddress_qZ0Z_4\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__11641\,
            I => \this_vga_signals.M_haddress_qZ0Z_4\
        );

    \I__2018\ : InMux
    port map (
            O => \N__11630\,
            I => \N__11627\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__11627\,
            I => \N__11624\
        );

    \I__2016\ : Span12Mux_s8_v
    port map (
            O => \N__11624\,
            I => \N__11621\
        );

    \I__2015\ : Odrv12
    port map (
            O => \N__11621\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_2\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__11618\,
            I => \N__11615\
        );

    \I__2013\ : CascadeBuf
    port map (
            O => \N__11615\,
            I => \N__11612\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__11612\,
            I => \N__11609\
        );

    \I__2011\ : CascadeBuf
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__11606\,
            I => \N__11603\
        );

    \I__2009\ : CascadeBuf
    port map (
            O => \N__11603\,
            I => \N__11600\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__11600\,
            I => \N__11597\
        );

    \I__2007\ : CascadeBuf
    port map (
            O => \N__11597\,
            I => \N__11594\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__11594\,
            I => \N__11591\
        );

    \I__2005\ : CascadeBuf
    port map (
            O => \N__11591\,
            I => \N__11588\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__11588\,
            I => \N__11585\
        );

    \I__2003\ : CascadeBuf
    port map (
            O => \N__11585\,
            I => \N__11582\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__11582\,
            I => \N__11579\
        );

    \I__2001\ : CascadeBuf
    port map (
            O => \N__11579\,
            I => \N__11576\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__11576\,
            I => \N__11573\
        );

    \I__1999\ : CascadeBuf
    port map (
            O => \N__11573\,
            I => \N__11570\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__11570\,
            I => \N__11567\
        );

    \I__1997\ : CascadeBuf
    port map (
            O => \N__11567\,
            I => \N__11564\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__11564\,
            I => \N__11561\
        );

    \I__1995\ : CascadeBuf
    port map (
            O => \N__11561\,
            I => \N__11558\
        );

    \I__1994\ : CascadeMux
    port map (
            O => \N__11558\,
            I => \N__11555\
        );

    \I__1993\ : CascadeBuf
    port map (
            O => \N__11555\,
            I => \N__11552\
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__11552\,
            I => \N__11549\
        );

    \I__1991\ : CascadeBuf
    port map (
            O => \N__11549\,
            I => \N__11546\
        );

    \I__1990\ : CascadeMux
    port map (
            O => \N__11546\,
            I => \N__11543\
        );

    \I__1989\ : CascadeBuf
    port map (
            O => \N__11543\,
            I => \N__11540\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__11540\,
            I => \N__11537\
        );

    \I__1987\ : CascadeBuf
    port map (
            O => \N__11537\,
            I => \N__11534\
        );

    \I__1986\ : CascadeMux
    port map (
            O => \N__11534\,
            I => \N__11531\
        );

    \I__1985\ : CascadeBuf
    port map (
            O => \N__11531\,
            I => \N__11528\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__11528\,
            I => \N__11525\
        );

    \I__1983\ : InMux
    port map (
            O => \N__11525\,
            I => \N__11522\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__11522\,
            I => \N__11519\
        );

    \I__1981\ : Odrv12
    port map (
            O => \N__11519\,
            I => this_vga_signals_un6_address_if_generate_plus_mult1_un68_sum_i_3
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__11516\,
            I => \N__11513\
        );

    \I__1979\ : InMux
    port map (
            O => \N__11513\,
            I => \N__11510\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__11510\,
            I => \N__11507\
        );

    \I__1977\ : Span12Mux_h
    port map (
            O => \N__11507\,
            I => \N__11504\
        );

    \I__1976\ : Odrv12
    port map (
            O => \N__11504\,
            I => \this_vga_signals.g0_14_N_8L16_sx\
        );

    \I__1975\ : InMux
    port map (
            O => \N__11501\,
            I => \N__11498\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__11498\,
            I => \this_vga_signals.mult1_un54_sum_c3_1_0_0\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__11495\,
            I => \N__11489\
        );

    \I__1972\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11486\
        );

    \I__1971\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11482\
        );

    \I__1970\ : InMux
    port map (
            O => \N__11492\,
            I => \N__11479\
        );

    \I__1969\ : InMux
    port map (
            O => \N__11489\,
            I => \N__11476\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__11486\,
            I => \N__11473\
        );

    \I__1967\ : InMux
    port map (
            O => \N__11485\,
            I => \N__11470\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__11482\,
            I => \N__11459\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__11479\,
            I => \N__11459\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__11476\,
            I => \N__11459\
        );

    \I__1963\ : Span4Mux_h
    port map (
            O => \N__11473\,
            I => \N__11459\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__11470\,
            I => \N__11459\
        );

    \I__1961\ : Span4Mux_v
    port map (
            O => \N__11459\,
            I => \N__11455\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__11458\,
            I => \N__11452\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__11455\,
            I => \N__11449\
        );

    \I__1958\ : InMux
    port map (
            O => \N__11452\,
            I => \N__11446\
        );

    \I__1957\ : Sp12to4
    port map (
            O => \N__11449\,
            I => \N__11441\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__11446\,
            I => \N__11441\
        );

    \I__1955\ : Odrv12
    port map (
            O => \N__11441\,
            I => \M_this_vram_read_data_3\
        );

    \I__1954\ : InMux
    port map (
            O => \N__11438\,
            I => \N__11434\
        );

    \I__1953\ : InMux
    port map (
            O => \N__11437\,
            I => \N__11431\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__11434\,
            I => \N__11427\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__11431\,
            I => \N__11424\
        );

    \I__1950\ : InMux
    port map (
            O => \N__11430\,
            I => \N__11421\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__11427\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__11424\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__11421\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0\
        );

    \I__1946\ : InMux
    port map (
            O => \N__11414\,
            I => \N__11410\
        );

    \I__1945\ : InMux
    port map (
            O => \N__11413\,
            I => \N__11405\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__11410\,
            I => \N__11402\
        );

    \I__1943\ : InMux
    port map (
            O => \N__11409\,
            I => \N__11397\
        );

    \I__1942\ : InMux
    port map (
            O => \N__11408\,
            I => \N__11397\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__11405\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__11402\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__11397\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__1938\ : InMux
    port map (
            O => \N__11390\,
            I => \N__11386\
        );

    \I__1937\ : InMux
    port map (
            O => \N__11389\,
            I => \N__11383\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__11386\,
            I => \this_start_data_delay.this_edge_detector.N_253_0\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__11383\,
            I => \this_start_data_delay.this_edge_detector.N_253_0\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__11378\,
            I => \N__11375\
        );

    \I__1933\ : InMux
    port map (
            O => \N__11375\,
            I => \N__11370\
        );

    \I__1932\ : InMux
    port map (
            O => \N__11374\,
            I => \N__11367\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__11373\,
            I => \N__11363\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__11370\,
            I => \N__11358\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__11367\,
            I => \N__11355\
        );

    \I__1928\ : InMux
    port map (
            O => \N__11366\,
            I => \N__11348\
        );

    \I__1927\ : InMux
    port map (
            O => \N__11363\,
            I => \N__11348\
        );

    \I__1926\ : InMux
    port map (
            O => \N__11362\,
            I => \N__11348\
        );

    \I__1925\ : InMux
    port map (
            O => \N__11361\,
            I => \N__11345\
        );

    \I__1924\ : Span4Mux_v
    port map (
            O => \N__11358\,
            I => \N__11342\
        );

    \I__1923\ : Span4Mux_v
    port map (
            O => \N__11355\,
            I => \N__11339\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__11348\,
            I => \N__11336\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__11345\,
            I => \this_vga_signals.M_haddress_qZ0Z_3\
        );

    \I__1920\ : Odrv4
    port map (
            O => \N__11342\,
            I => \this_vga_signals.M_haddress_qZ0Z_3\
        );

    \I__1919\ : Odrv4
    port map (
            O => \N__11339\,
            I => \this_vga_signals.M_haddress_qZ0Z_3\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__11336\,
            I => \this_vga_signals.M_haddress_qZ0Z_3\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__11327\,
            I => \this_start_data_delay.this_edge_detector.N_261_cascade_\
        );

    \I__1916\ : InMux
    port map (
            O => \N__11324\,
            I => \N__11321\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__11321\,
            I => \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_0Z0Z_0\
        );

    \I__1914\ : InMux
    port map (
            O => \N__11318\,
            I => \N__11315\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__11315\,
            I => \M_this_start_address_delay_out_0\
        );

    \I__1912\ : InMux
    port map (
            O => \N__11312\,
            I => \N__11308\
        );

    \I__1911\ : InMux
    port map (
            O => \N__11311\,
            I => \N__11305\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__11308\,
            I => \this_start_data_delay.this_edge_detector.N_267\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__11305\,
            I => \this_start_data_delay.this_edge_detector.N_267\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__11300\,
            I => \this_start_data_delay.this_edge_detector.N_275_cascade_\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__11297\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0_cascade_\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__11294\,
            I => \N__11291\
        );

    \I__1905\ : InMux
    port map (
            O => \N__11291\,
            I => \N__11288\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__11288\,
            I => \N__11285\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__11285\,
            I => \this_vga_signals.g0_0_0_0\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__11282\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_cascade_\
        );

    \I__1901\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11272\
        );

    \I__1900\ : InMux
    port map (
            O => \N__11278\,
            I => \N__11272\
        );

    \I__1899\ : InMux
    port map (
            O => \N__11277\,
            I => \N__11269\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__11272\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_0\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__11269\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_0\
        );

    \I__1896\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11261\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__11261\,
            I => \N__11258\
        );

    \I__1894\ : Odrv12
    port map (
            O => \N__11258\,
            I => \this_vga_signals.mult1_un54_sum_axb1_0\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__11255\,
            I => \this_vga_signals.g0_0_5_1_cascade_\
        );

    \I__1892\ : CascadeMux
    port map (
            O => \N__11252\,
            I => \N__11249\
        );

    \I__1891\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11246\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__11246\,
            I => \this_vga_signals.g0_3_1\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__11243\,
            I => \this_vga_signals.if_N_2_1_0_cascade_\
        );

    \I__1888\ : InMux
    port map (
            O => \N__11240\,
            I => \N__11236\
        );

    \I__1887\ : InMux
    port map (
            O => \N__11239\,
            I => \N__11233\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__11236\,
            I => \N__11230\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__11233\,
            I => \this_vga_signals.mult1_un54_sum_axb1_0_0_1_1\
        );

    \I__1884\ : Odrv12
    port map (
            O => \N__11230\,
            I => \this_vga_signals.mult1_un54_sum_axb1_0_0_1_1\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__11225\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d_cascade_\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__11222\,
            I => \this_vga_signals.if_N_2_1_1_cascade_\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__11219\,
            I => \this_vga_signals.mult1_un54_sum_c3_2_cascade_\
        );

    \I__1880\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11213\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__11213\,
            I => \this_vga_signals.N_3_1_0\
        );

    \I__1878\ : InMux
    port map (
            O => \N__11210\,
            I => \N__11207\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__11207\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_1_x\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__11204\,
            I => \this_vga_signals.g0_3_0_cascade_\
        );

    \I__1875\ : InMux
    port map (
            O => \N__11201\,
            I => \N__11198\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__11198\,
            I => \this_vga_signals.if_N_2_5\
        );

    \I__1873\ : InMux
    port map (
            O => \N__11195\,
            I => \N__11188\
        );

    \I__1872\ : InMux
    port map (
            O => \N__11194\,
            I => \N__11188\
        );

    \I__1871\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11185\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__11188\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__11185\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__1868\ : InMux
    port map (
            O => \N__11180\,
            I => \N__11177\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__11177\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_18\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__11174\,
            I => \this_start_data_delay.this_edge_detector.N_267_cascade_\
        );

    \I__1865\ : InMux
    port map (
            O => \N__11171\,
            I => \N__11168\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__11168\,
            I => \N__11165\
        );

    \I__1863\ : Span12Mux_s3_v
    port map (
            O => \N__11165\,
            I => \N__11162\
        );

    \I__1862\ : Span12Mux_v
    port map (
            O => \N__11162\,
            I => \N__11159\
        );

    \I__1861\ : Odrv12
    port map (
            O => \N__11159\,
            I => \this_vga_signals.if_m12_bm\
        );

    \I__1860\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11153\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__11153\,
            I => \N__11150\
        );

    \I__1858\ : Span4Mux_v
    port map (
            O => \N__11150\,
            I => \N__11147\
        );

    \I__1857\ : Span4Mux_v
    port map (
            O => \N__11147\,
            I => \N__11144\
        );

    \I__1856\ : Span4Mux_v
    port map (
            O => \N__11144\,
            I => \N__11141\
        );

    \I__1855\ : Span4Mux_v
    port map (
            O => \N__11141\,
            I => \N__11138\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__11138\,
            I => \this_vga_signals.if_m12_am\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11135\,
            I => \N__11132\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__11132\,
            I => \N__11129\
        );

    \I__1851\ : Span12Mux_s5_v
    port map (
            O => \N__11129\,
            I => \N__11126\
        );

    \I__1850\ : Span12Mux_v
    port map (
            O => \N__11126\,
            I => \N__11123\
        );

    \I__1849\ : Odrv12
    port map (
            O => \N__11123\,
            I => \this_vga_signals.if_m13_ns_1\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__11120\,
            I => \N__11117\
        );

    \I__1847\ : CascadeBuf
    port map (
            O => \N__11117\,
            I => \N__11114\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__11114\,
            I => \N__11111\
        );

    \I__1845\ : CascadeBuf
    port map (
            O => \N__11111\,
            I => \N__11108\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__11108\,
            I => \N__11105\
        );

    \I__1843\ : CascadeBuf
    port map (
            O => \N__11105\,
            I => \N__11102\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__11102\,
            I => \N__11099\
        );

    \I__1841\ : CascadeBuf
    port map (
            O => \N__11099\,
            I => \N__11096\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__11096\,
            I => \N__11093\
        );

    \I__1839\ : CascadeBuf
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__11090\,
            I => \N__11087\
        );

    \I__1837\ : CascadeBuf
    port map (
            O => \N__11087\,
            I => \N__11084\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__11084\,
            I => \N__11081\
        );

    \I__1835\ : CascadeBuf
    port map (
            O => \N__11081\,
            I => \N__11078\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__11078\,
            I => \N__11075\
        );

    \I__1833\ : CascadeBuf
    port map (
            O => \N__11075\,
            I => \N__11072\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__11072\,
            I => \N__11069\
        );

    \I__1831\ : CascadeBuf
    port map (
            O => \N__11069\,
            I => \N__11066\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__11066\,
            I => \N__11063\
        );

    \I__1829\ : CascadeBuf
    port map (
            O => \N__11063\,
            I => \N__11060\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__11060\,
            I => \N__11057\
        );

    \I__1827\ : CascadeBuf
    port map (
            O => \N__11057\,
            I => \N__11054\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__11054\,
            I => \N__11051\
        );

    \I__1825\ : CascadeBuf
    port map (
            O => \N__11051\,
            I => \N__11048\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__11048\,
            I => \N__11045\
        );

    \I__1823\ : CascadeBuf
    port map (
            O => \N__11045\,
            I => \N__11042\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__11042\,
            I => \N__11039\
        );

    \I__1821\ : CascadeBuf
    port map (
            O => \N__11039\,
            I => \N__11036\
        );

    \I__1820\ : CascadeMux
    port map (
            O => \N__11036\,
            I => \N__11033\
        );

    \I__1819\ : CascadeBuf
    port map (
            O => \N__11033\,
            I => \N__11030\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__11030\,
            I => \N__11027\
        );

    \I__1817\ : InMux
    port map (
            O => \N__11027\,
            I => \N__11024\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__11024\,
            I => \N__11021\
        );

    \I__1815\ : Odrv12
    port map (
            O => \N__11021\,
            I => if_m13_ns
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__11018\,
            I => \this_vga_signals.N_9_0_0_cascade_\
        );

    \I__1813\ : InMux
    port map (
            O => \N__11015\,
            I => \N__11012\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__11012\,
            I => \N__11009\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__11009\,
            I => \N__11006\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__11006\,
            I => \this_vga_signals.g0_4_2\
        );

    \I__1809\ : InMux
    port map (
            O => \N__11003\,
            I => \N__11000\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__11000\,
            I => \this_vga_signals.mult1_un40_sum_1_ac0_2\
        );

    \I__1807\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10994\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__10994\,
            I => \N__10991\
        );

    \I__1805\ : Span4Mux_h
    port map (
            O => \N__10991\,
            I => \N__10988\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__10988\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_15\
        );

    \I__1803\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10982\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__10982\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_18\
        );

    \I__1801\ : InMux
    port map (
            O => \N__10979\,
            I => \N__10976\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__10976\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_16\
        );

    \I__1799\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10970\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__10970\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_17\
        );

    \I__1797\ : InMux
    port map (
            O => \N__10967\,
            I => \N__10964\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__10964\,
            I => \M_state_qZ0Z_5\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__10961\,
            I => \N__10958\
        );

    \I__1794\ : InMux
    port map (
            O => \N__10958\,
            I => \N__10955\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__10955\,
            I => \this_start_data_delay.this_edge_detector.N_252_0\
        );

    \I__1792\ : InMux
    port map (
            O => \N__10952\,
            I => \N__10949\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__10949\,
            I => \N__10946\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__10946\,
            I => \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_o3_0_0\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__10943\,
            I => \this_start_data_delay.this_edge_detector.N_252_0_cascade_\
        );

    \I__1788\ : InMux
    port map (
            O => \N__10940\,
            I => \N__10936\
        );

    \I__1787\ : InMux
    port map (
            O => \N__10939\,
            I => \N__10933\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__10936\,
            I => \this_vga_signals.mult1_un40_sum_1_axb1\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__10933\,
            I => \this_vga_signals.mult1_un40_sum_1_axb1\
        );

    \I__1784\ : InMux
    port map (
            O => \N__10928\,
            I => \N__10924\
        );

    \I__1783\ : InMux
    port map (
            O => \N__10927\,
            I => \N__10921\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__10924\,
            I => \this_vga_signals.mult1_un40_sum_1_c2_0\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__10921\,
            I => \this_vga_signals.mult1_un40_sum_1_c2_0\
        );

    \I__1780\ : CascadeMux
    port map (
            O => \N__10916\,
            I => \N__10913\
        );

    \I__1779\ : InMux
    port map (
            O => \N__10913\,
            I => \N__10907\
        );

    \I__1778\ : InMux
    port map (
            O => \N__10912\,
            I => \N__10907\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__10907\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc2_0\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__10904\,
            I => \this_vga_signals.N_2_1_1_cascade_\
        );

    \I__1775\ : CascadeMux
    port map (
            O => \N__10901\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc3_a4_cascade_\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__10898\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_cascade_\
        );

    \I__1773\ : InMux
    port map (
            O => \N__10895\,
            I => \N__10892\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__10892\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_0\
        );

    \I__1771\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10886\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__10886\,
            I => \this_vga_signals.mult1_un40_sum1_0_3\
        );

    \I__1769\ : InMux
    port map (
            O => \N__10883\,
            I => \N__10875\
        );

    \I__1768\ : InMux
    port map (
            O => \N__10882\,
            I => \N__10868\
        );

    \I__1767\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10868\
        );

    \I__1766\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10863\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__10879\,
            I => \N__10855\
        );

    \I__1764\ : InMux
    port map (
            O => \N__10878\,
            I => \N__10851\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__10875\,
            I => \N__10848\
        );

    \I__1762\ : InMux
    port map (
            O => \N__10874\,
            I => \N__10843\
        );

    \I__1761\ : InMux
    port map (
            O => \N__10873\,
            I => \N__10843\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__10868\,
            I => \N__10840\
        );

    \I__1759\ : InMux
    port map (
            O => \N__10867\,
            I => \N__10835\
        );

    \I__1758\ : InMux
    port map (
            O => \N__10866\,
            I => \N__10835\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__10863\,
            I => \N__10832\
        );

    \I__1756\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10829\
        );

    \I__1755\ : InMux
    port map (
            O => \N__10861\,
            I => \N__10824\
        );

    \I__1754\ : InMux
    port map (
            O => \N__10860\,
            I => \N__10824\
        );

    \I__1753\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10815\
        );

    \I__1752\ : InMux
    port map (
            O => \N__10858\,
            I => \N__10815\
        );

    \I__1751\ : InMux
    port map (
            O => \N__10855\,
            I => \N__10815\
        );

    \I__1750\ : InMux
    port map (
            O => \N__10854\,
            I => \N__10815\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__10851\,
            I => \this_vga_signals.M_haddress_qZ0Z_7\
        );

    \I__1748\ : Odrv12
    port map (
            O => \N__10848\,
            I => \this_vga_signals.M_haddress_qZ0Z_7\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__10843\,
            I => \this_vga_signals.M_haddress_qZ0Z_7\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__10840\,
            I => \this_vga_signals.M_haddress_qZ0Z_7\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__10835\,
            I => \this_vga_signals.M_haddress_qZ0Z_7\
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__10832\,
            I => \this_vga_signals.M_haddress_qZ0Z_7\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__10829\,
            I => \this_vga_signals.M_haddress_qZ0Z_7\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__10824\,
            I => \this_vga_signals.M_haddress_qZ0Z_7\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__10815\,
            I => \this_vga_signals.M_haddress_qZ0Z_7\
        );

    \I__1740\ : InMux
    port map (
            O => \N__10796\,
            I => \N__10793\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__10793\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc3_a5\
        );

    \I__1738\ : InMux
    port map (
            O => \N__10790\,
            I => \N__10787\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__10787\,
            I => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_1\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__10784\,
            I => \this_vga_signals.g1_0_1_cascade_\
        );

    \I__1735\ : InMux
    port map (
            O => \N__10781\,
            I => \N__10778\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__10778\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_1\
        );

    \I__1733\ : InMux
    port map (
            O => \N__10775\,
            I => \N__10772\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__10772\,
            I => \this_vga_signals.g0_0_0_2\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__10769\,
            I => \N__10766\
        );

    \I__1730\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10763\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__10763\,
            I => \this_vga_signals.g0_29_1\
        );

    \I__1728\ : InMux
    port map (
            O => \N__10760\,
            I => \N__10757\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__10757\,
            I => \this_vga_signals.N_3_0_0_0\
        );

    \I__1726\ : InMux
    port map (
            O => \N__10754\,
            I => \N__10751\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__10751\,
            I => \N__10748\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__10748\,
            I => \this_vga_signals.if_N_7\
        );

    \I__1723\ : InMux
    port map (
            O => \N__10745\,
            I => \N__10735\
        );

    \I__1722\ : InMux
    port map (
            O => \N__10744\,
            I => \N__10735\
        );

    \I__1721\ : InMux
    port map (
            O => \N__10743\,
            I => \N__10735\
        );

    \I__1720\ : InMux
    port map (
            O => \N__10742\,
            I => \N__10729\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__10735\,
            I => \N__10726\
        );

    \I__1718\ : InMux
    port map (
            O => \N__10734\,
            I => \N__10723\
        );

    \I__1717\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10720\
        );

    \I__1716\ : InMux
    port map (
            O => \N__10732\,
            I => \N__10717\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__10729\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__10726\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__10723\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__10720\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__10717\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__1710\ : InMux
    port map (
            O => \N__10706\,
            I => \N__10703\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__10703\,
            I => \N__10698\
        );

    \I__1708\ : InMux
    port map (
            O => \N__10702\,
            I => \N__10695\
        );

    \I__1707\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10692\
        );

    \I__1706\ : Odrv4
    port map (
            O => \N__10698\,
            I => \this_vga_signals.mult1_un40_sum_m_2\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__10695\,
            I => \this_vga_signals.mult1_un40_sum_m_2\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__10692\,
            I => \this_vga_signals.mult1_un40_sum_m_2\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__10685\,
            I => \N__10682\
        );

    \I__1702\ : CascadeBuf
    port map (
            O => \N__10682\,
            I => \N__10679\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__10679\,
            I => \N__10676\
        );

    \I__1700\ : CascadeBuf
    port map (
            O => \N__10676\,
            I => \N__10673\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__10673\,
            I => \N__10670\
        );

    \I__1698\ : CascadeBuf
    port map (
            O => \N__10670\,
            I => \N__10667\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__10667\,
            I => \N__10664\
        );

    \I__1696\ : CascadeBuf
    port map (
            O => \N__10664\,
            I => \N__10661\
        );

    \I__1695\ : CascadeMux
    port map (
            O => \N__10661\,
            I => \N__10658\
        );

    \I__1694\ : CascadeBuf
    port map (
            O => \N__10658\,
            I => \N__10655\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__10655\,
            I => \N__10652\
        );

    \I__1692\ : CascadeBuf
    port map (
            O => \N__10652\,
            I => \N__10649\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__10649\,
            I => \N__10646\
        );

    \I__1690\ : CascadeBuf
    port map (
            O => \N__10646\,
            I => \N__10643\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__10643\,
            I => \N__10640\
        );

    \I__1688\ : CascadeBuf
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__10637\,
            I => \N__10634\
        );

    \I__1686\ : CascadeBuf
    port map (
            O => \N__10634\,
            I => \N__10631\
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__10631\,
            I => \N__10628\
        );

    \I__1684\ : CascadeBuf
    port map (
            O => \N__10628\,
            I => \N__10625\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__10625\,
            I => \N__10622\
        );

    \I__1682\ : CascadeBuf
    port map (
            O => \N__10622\,
            I => \N__10619\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__10619\,
            I => \N__10616\
        );

    \I__1680\ : CascadeBuf
    port map (
            O => \N__10616\,
            I => \N__10613\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__10613\,
            I => \N__10610\
        );

    \I__1678\ : CascadeBuf
    port map (
            O => \N__10610\,
            I => \N__10607\
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__10607\,
            I => \N__10604\
        );

    \I__1676\ : CascadeBuf
    port map (
            O => \N__10604\,
            I => \N__10601\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__10601\,
            I => \N__10598\
        );

    \I__1674\ : CascadeBuf
    port map (
            O => \N__10598\,
            I => \N__10595\
        );

    \I__1673\ : CascadeMux
    port map (
            O => \N__10595\,
            I => \N__10592\
        );

    \I__1672\ : InMux
    port map (
            O => \N__10592\,
            I => \N__10589\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__10589\,
            I => \N__10586\
        );

    \I__1670\ : Span4Mux_v
    port map (
            O => \N__10586\,
            I => \N__10583\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__10583\,
            I => \N__10580\
        );

    \I__1668\ : Sp12to4
    port map (
            O => \N__10580\,
            I => \N__10572\
        );

    \I__1667\ : InMux
    port map (
            O => \N__10579\,
            I => \N__10569\
        );

    \I__1666\ : InMux
    port map (
            O => \N__10578\,
            I => \N__10564\
        );

    \I__1665\ : InMux
    port map (
            O => \N__10577\,
            I => \N__10564\
        );

    \I__1664\ : InMux
    port map (
            O => \N__10576\,
            I => \N__10559\
        );

    \I__1663\ : InMux
    port map (
            O => \N__10575\,
            I => \N__10559\
        );

    \I__1662\ : Span12Mux_h
    port map (
            O => \N__10572\,
            I => \N__10556\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__10569\,
            I => \this_vga_signals_un6_address_if_N_5_mux_0\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__10564\,
            I => \this_vga_signals_un6_address_if_N_5_mux_0\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__10559\,
            I => \this_vga_signals_un6_address_if_N_5_mux_0\
        );

    \I__1658\ : Odrv12
    port map (
            O => \N__10556\,
            I => \this_vga_signals_un6_address_if_N_5_mux_0\
        );

    \I__1657\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10539\
        );

    \I__1656\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10539\
        );

    \I__1655\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10534\
        );

    \I__1654\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10534\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__10539\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__10534\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0\
        );

    \I__1651\ : CascadeMux
    port map (
            O => \N__10529\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0_cascade_\
        );

    \I__1650\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10519\
        );

    \I__1649\ : InMux
    port map (
            O => \N__10525\,
            I => \N__10516\
        );

    \I__1648\ : InMux
    port map (
            O => \N__10524\,
            I => \N__10509\
        );

    \I__1647\ : InMux
    port map (
            O => \N__10523\,
            I => \N__10509\
        );

    \I__1646\ : InMux
    port map (
            O => \N__10522\,
            I => \N__10509\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__10519\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__10516\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__10509\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__10502\,
            I => \N__10499\
        );

    \I__1641\ : CascadeBuf
    port map (
            O => \N__10499\,
            I => \N__10496\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__10496\,
            I => \N__10493\
        );

    \I__1639\ : CascadeBuf
    port map (
            O => \N__10493\,
            I => \N__10490\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__10490\,
            I => \N__10487\
        );

    \I__1637\ : CascadeBuf
    port map (
            O => \N__10487\,
            I => \N__10484\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__10484\,
            I => \N__10481\
        );

    \I__1635\ : CascadeBuf
    port map (
            O => \N__10481\,
            I => \N__10478\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__10478\,
            I => \N__10475\
        );

    \I__1633\ : CascadeBuf
    port map (
            O => \N__10475\,
            I => \N__10472\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__10472\,
            I => \N__10469\
        );

    \I__1631\ : CascadeBuf
    port map (
            O => \N__10469\,
            I => \N__10466\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__10466\,
            I => \N__10463\
        );

    \I__1629\ : CascadeBuf
    port map (
            O => \N__10463\,
            I => \N__10460\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__10460\,
            I => \N__10457\
        );

    \I__1627\ : CascadeBuf
    port map (
            O => \N__10457\,
            I => \N__10454\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__10454\,
            I => \N__10451\
        );

    \I__1625\ : CascadeBuf
    port map (
            O => \N__10451\,
            I => \N__10448\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__10448\,
            I => \N__10445\
        );

    \I__1623\ : CascadeBuf
    port map (
            O => \N__10445\,
            I => \N__10442\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__10442\,
            I => \N__10439\
        );

    \I__1621\ : CascadeBuf
    port map (
            O => \N__10439\,
            I => \N__10436\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__10436\,
            I => \N__10433\
        );

    \I__1619\ : CascadeBuf
    port map (
            O => \N__10433\,
            I => \N__10430\
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__10430\,
            I => \N__10427\
        );

    \I__1617\ : CascadeBuf
    port map (
            O => \N__10427\,
            I => \N__10424\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__10424\,
            I => \N__10421\
        );

    \I__1615\ : CascadeBuf
    port map (
            O => \N__10421\,
            I => \N__10418\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__10418\,
            I => \N__10415\
        );

    \I__1613\ : CascadeBuf
    port map (
            O => \N__10415\,
            I => \N__10412\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__10412\,
            I => \N__10409\
        );

    \I__1611\ : InMux
    port map (
            O => \N__10409\,
            I => \N__10406\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__10406\,
            I => \N__10403\
        );

    \I__1609\ : Span4Mux_h
    port map (
            O => \N__10403\,
            I => \N__10400\
        );

    \I__1608\ : Span4Mux_h
    port map (
            O => \N__10400\,
            I => \N__10397\
        );

    \I__1607\ : Sp12to4
    port map (
            O => \N__10397\,
            I => \N__10394\
        );

    \I__1606\ : Span12Mux_v
    port map (
            O => \N__10394\,
            I => \N__10391\
        );

    \I__1605\ : Odrv12
    port map (
            O => \N__10391\,
            I => this_vga_signals_un6_address_if_generate_plus_mult1_un47_sum_i_3
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__10388\,
            I => \N__10384\
        );

    \I__1603\ : InMux
    port map (
            O => \N__10387\,
            I => \N__10378\
        );

    \I__1602\ : InMux
    port map (
            O => \N__10384\,
            I => \N__10378\
        );

    \I__1601\ : InMux
    port map (
            O => \N__10383\,
            I => \N__10375\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__10378\,
            I => \this_vga_signals.mult1_un40_sum_m_1\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__10375\,
            I => \this_vga_signals.mult1_un40_sum_m_1\
        );

    \I__1598\ : InMux
    port map (
            O => \N__10370\,
            I => \N__10360\
        );

    \I__1597\ : InMux
    port map (
            O => \N__10369\,
            I => \N__10360\
        );

    \I__1596\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10360\
        );

    \I__1595\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10357\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__10360\,
            I => \this_vga_signals.CO1_1_0\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__10357\,
            I => \this_vga_signals.CO1_1_0\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__10352\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\
        );

    \I__1591\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10346\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__10346\,
            I => \this_vga_signals.if_m1\
        );

    \I__1589\ : InMux
    port map (
            O => \N__10343\,
            I => \N__10339\
        );

    \I__1588\ : InMux
    port map (
            O => \N__10342\,
            I => \N__10336\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__10339\,
            I => \this_vga_signals.mult1_un54_sum_axb1_2\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__10336\,
            I => \this_vga_signals.mult1_un54_sum_axb1_2\
        );

    \I__1585\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__10328\,
            I => \this_vga_signals.g1_N_2L1\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__10325\,
            I => \N__10322\
        );

    \I__1582\ : InMux
    port map (
            O => \N__10322\,
            I => \N__10319\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__10319\,
            I => \this_vga_signals.G_5_0_x2_1\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__10316\,
            I => \this_vga_signals.mult1_un54_sum_axb1_cascade_\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__10313\,
            I => \this_vga_signals.g2_4_cascade_\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__10310\,
            I => \N__10307\
        );

    \I__1577\ : InMux
    port map (
            O => \N__10307\,
            I => \N__10304\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__10304\,
            I => \this_vga_signals.if_m1_3\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__10301\,
            I => \this_vga_signals.if_m1_3_cascade_\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__10298\,
            I => \this_vga_signals.if_m8_am_cascade_\
        );

    \I__1573\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10292\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__10292\,
            I => \this_vga_signals.if_m8_bm\
        );

    \I__1571\ : InMux
    port map (
            O => \N__10289\,
            I => \N__10286\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__10286\,
            I => \this_vga_signals.g1_0_0\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__10283\,
            I => \this_vga_signals.g0_0_2_cascade_\
        );

    \I__1568\ : InMux
    port map (
            O => \N__10280\,
            I => \N__10277\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__10277\,
            I => \this_vga_signals.g0_0_3_0\
        );

    \I__1566\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10271\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__10271\,
            I => \N__10268\
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__10268\,
            I => \this_vga_signals.g3_2\
        );

    \I__1563\ : InMux
    port map (
            O => \N__10265\,
            I => \N__10262\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__10262\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_0_0_1\
        );

    \I__1561\ : InMux
    port map (
            O => \N__10259\,
            I => \this_vga_signals.un1_M_haddress_q_cry_9\
        );

    \I__1560\ : InMux
    port map (
            O => \N__10256\,
            I => \this_vga_signals.un1_M_haddress_q_cry_10\
        );

    \I__1559\ : SRMux
    port map (
            O => \N__10253\,
            I => \N__10249\
        );

    \I__1558\ : SRMux
    port map (
            O => \N__10252\,
            I => \N__10246\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__10249\,
            I => \N__10243\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__10246\,
            I => \N__10240\
        );

    \I__1555\ : Span4Mux_h
    port map (
            O => \N__10243\,
            I => \N__10237\
        );

    \I__1554\ : Span4Mux_h
    port map (
            O => \N__10240\,
            I => \N__10234\
        );

    \I__1553\ : Span4Mux_h
    port map (
            O => \N__10237\,
            I => \N__10231\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__10234\,
            I => \this_vga_signals.M_hstate_q_RNIFIH84Z0Z_5\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__10231\,
            I => \this_vga_signals.M_hstate_q_RNIFIH84Z0Z_5\
        );

    \I__1550\ : InMux
    port map (
            O => \N__10226\,
            I => \N__10223\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__10223\,
            I => \N__10220\
        );

    \I__1548\ : Span4Mux_h
    port map (
            O => \N__10220\,
            I => \N__10217\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__10217\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_16\
        );

    \I__1546\ : InMux
    port map (
            O => \N__10214\,
            I => \N__10211\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__10211\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_17\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10208\,
            I => \N__10205\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__10205\,
            I => \N__10199\
        );

    \I__1542\ : InMux
    port map (
            O => \N__10204\,
            I => \N__10196\
        );

    \I__1541\ : InMux
    port map (
            O => \N__10203\,
            I => \N__10193\
        );

    \I__1540\ : InMux
    port map (
            O => \N__10202\,
            I => \N__10190\
        );

    \I__1539\ : Odrv12
    port map (
            O => \N__10199\,
            I => \this_vga_signals.mult1_un54_sum_c3\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__10196\,
            I => \this_vga_signals.mult1_un54_sum_c3\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__10193\,
            I => \this_vga_signals.mult1_un54_sum_c3\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__10190\,
            I => \this_vga_signals.mult1_un54_sum_c3\
        );

    \I__1535\ : InMux
    port map (
            O => \N__10181\,
            I => \N__10178\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__10178\,
            I => \N__10171\
        );

    \I__1533\ : InMux
    port map (
            O => \N__10177\,
            I => \N__10166\
        );

    \I__1532\ : InMux
    port map (
            O => \N__10176\,
            I => \N__10166\
        );

    \I__1531\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10163\
        );

    \I__1530\ : InMux
    port map (
            O => \N__10174\,
            I => \N__10160\
        );

    \I__1529\ : Odrv12
    port map (
            O => \N__10171\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0_i\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__10166\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0_i\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__10163\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0_i\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__10160\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_0_i\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__10151\,
            I => \N__10148\
        );

    \I__1524\ : CascadeBuf
    port map (
            O => \N__10148\,
            I => \N__10145\
        );

    \I__1523\ : CascadeMux
    port map (
            O => \N__10145\,
            I => \N__10142\
        );

    \I__1522\ : CascadeBuf
    port map (
            O => \N__10142\,
            I => \N__10139\
        );

    \I__1521\ : CascadeMux
    port map (
            O => \N__10139\,
            I => \N__10136\
        );

    \I__1520\ : CascadeBuf
    port map (
            O => \N__10136\,
            I => \N__10133\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__10133\,
            I => \N__10130\
        );

    \I__1518\ : CascadeBuf
    port map (
            O => \N__10130\,
            I => \N__10127\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__10127\,
            I => \N__10124\
        );

    \I__1516\ : CascadeBuf
    port map (
            O => \N__10124\,
            I => \N__10121\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__10121\,
            I => \N__10118\
        );

    \I__1514\ : CascadeBuf
    port map (
            O => \N__10118\,
            I => \N__10115\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__10115\,
            I => \N__10112\
        );

    \I__1512\ : CascadeBuf
    port map (
            O => \N__10112\,
            I => \N__10109\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__10109\,
            I => \N__10106\
        );

    \I__1510\ : CascadeBuf
    port map (
            O => \N__10106\,
            I => \N__10103\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__10103\,
            I => \N__10100\
        );

    \I__1508\ : CascadeBuf
    port map (
            O => \N__10100\,
            I => \N__10097\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__10097\,
            I => \N__10094\
        );

    \I__1506\ : CascadeBuf
    port map (
            O => \N__10094\,
            I => \N__10091\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__10091\,
            I => \N__10088\
        );

    \I__1504\ : CascadeBuf
    port map (
            O => \N__10088\,
            I => \N__10085\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__10085\,
            I => \N__10082\
        );

    \I__1502\ : CascadeBuf
    port map (
            O => \N__10082\,
            I => \N__10079\
        );

    \I__1501\ : CascadeMux
    port map (
            O => \N__10079\,
            I => \N__10076\
        );

    \I__1500\ : CascadeBuf
    port map (
            O => \N__10076\,
            I => \N__10073\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__10073\,
            I => \N__10070\
        );

    \I__1498\ : CascadeBuf
    port map (
            O => \N__10070\,
            I => \N__10067\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__10067\,
            I => \N__10064\
        );

    \I__1496\ : CascadeBuf
    port map (
            O => \N__10064\,
            I => \N__10061\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__10061\,
            I => \N__10058\
        );

    \I__1494\ : InMux
    port map (
            O => \N__10058\,
            I => \N__10055\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__10055\,
            I => \N__10052\
        );

    \I__1492\ : Sp12to4
    port map (
            O => \N__10052\,
            I => \N__10049\
        );

    \I__1491\ : Span12Mux_h
    port map (
            O => \N__10049\,
            I => \N__10046\
        );

    \I__1490\ : Span12Mux_v
    port map (
            O => \N__10046\,
            I => \N__10043\
        );

    \I__1489\ : Odrv12
    port map (
            O => \N__10043\,
            I => this_vga_signals_un6_address_if_generate_plus_mult1_un54_sum_i_3
        );

    \I__1488\ : CascadeMux
    port map (
            O => \N__10040\,
            I => \this_vga_signals.g1_3_1_cascade_\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__10037\,
            I => \this_vga_signals.if_N_7_cascade_\
        );

    \I__1486\ : InMux
    port map (
            O => \N__10034\,
            I => \this_vga_signals.un1_M_haddress_q_cry_0\
        );

    \I__1485\ : InMux
    port map (
            O => \N__10031\,
            I => \N__10027\
        );

    \I__1484\ : InMux
    port map (
            O => \N__10030\,
            I => \N__10024\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__10027\,
            I => \N__10021\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__10024\,
            I => \this_vga_signals.M_haddress_qZ0Z_2\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__10021\,
            I => \this_vga_signals.M_haddress_qZ0Z_2\
        );

    \I__1480\ : InMux
    port map (
            O => \N__10016\,
            I => \this_vga_signals.un1_M_haddress_q_cry_1\
        );

    \I__1479\ : InMux
    port map (
            O => \N__10013\,
            I => \this_vga_signals.un1_M_haddress_q_cry_2\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10010\,
            I => \this_vga_signals.un1_M_haddress_q_cry_3\
        );

    \I__1477\ : InMux
    port map (
            O => \N__10007\,
            I => \N__10002\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__10006\,
            I => \N__9996\
        );

    \I__1475\ : CascadeMux
    port map (
            O => \N__10005\,
            I => \N__9992\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__10002\,
            I => \N__9988\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9985\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__10000\,
            I => \N__9981\
        );

    \I__1471\ : InMux
    port map (
            O => \N__9999\,
            I => \N__9978\
        );

    \I__1470\ : InMux
    port map (
            O => \N__9996\,
            I => \N__9975\
        );

    \I__1469\ : InMux
    port map (
            O => \N__9995\,
            I => \N__9968\
        );

    \I__1468\ : InMux
    port map (
            O => \N__9992\,
            I => \N__9968\
        );

    \I__1467\ : InMux
    port map (
            O => \N__9991\,
            I => \N__9968\
        );

    \I__1466\ : Span4Mux_h
    port map (
            O => \N__9988\,
            I => \N__9965\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__9985\,
            I => \N__9962\
        );

    \I__1464\ : InMux
    port map (
            O => \N__9984\,
            I => \N__9957\
        );

    \I__1463\ : InMux
    port map (
            O => \N__9981\,
            I => \N__9957\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__9978\,
            I => \this_vga_signals.M_haddress_qZ0Z_5\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__9975\,
            I => \this_vga_signals.M_haddress_qZ0Z_5\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__9968\,
            I => \this_vga_signals.M_haddress_qZ0Z_5\
        );

    \I__1459\ : Odrv4
    port map (
            O => \N__9965\,
            I => \this_vga_signals.M_haddress_qZ0Z_5\
        );

    \I__1458\ : Odrv4
    port map (
            O => \N__9962\,
            I => \this_vga_signals.M_haddress_qZ0Z_5\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__9957\,
            I => \this_vga_signals.M_haddress_qZ0Z_5\
        );

    \I__1456\ : InMux
    port map (
            O => \N__9944\,
            I => \this_vga_signals.un1_M_haddress_q_cry_4\
        );

    \I__1455\ : CascadeMux
    port map (
            O => \N__9941\,
            I => \N__9937\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__9940\,
            I => \N__9934\
        );

    \I__1453\ : InMux
    port map (
            O => \N__9937\,
            I => \N__9925\
        );

    \I__1452\ : InMux
    port map (
            O => \N__9934\,
            I => \N__9925\
        );

    \I__1451\ : InMux
    port map (
            O => \N__9933\,
            I => \N__9925\
        );

    \I__1450\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9917\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__9925\,
            I => \N__9914\
        );

    \I__1448\ : InMux
    port map (
            O => \N__9924\,
            I => \N__9911\
        );

    \I__1447\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9908\
        );

    \I__1446\ : InMux
    port map (
            O => \N__9922\,
            I => \N__9901\
        );

    \I__1445\ : InMux
    port map (
            O => \N__9921\,
            I => \N__9901\
        );

    \I__1444\ : InMux
    port map (
            O => \N__9920\,
            I => \N__9901\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__9917\,
            I => \this_vga_signals.M_haddress_qZ0Z_6\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__9914\,
            I => \this_vga_signals.M_haddress_qZ0Z_6\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__9911\,
            I => \this_vga_signals.M_haddress_qZ0Z_6\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__9908\,
            I => \this_vga_signals.M_haddress_qZ0Z_6\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__9901\,
            I => \this_vga_signals.M_haddress_qZ0Z_6\
        );

    \I__1438\ : InMux
    port map (
            O => \N__9890\,
            I => \this_vga_signals.un1_M_haddress_q_cry_5\
        );

    \I__1437\ : InMux
    port map (
            O => \N__9887\,
            I => \this_vga_signals.un1_M_haddress_q_cry_6\
        );

    \I__1436\ : InMux
    port map (
            O => \N__9884\,
            I => \bfn_18_16_0_\
        );

    \I__1435\ : InMux
    port map (
            O => \N__9881\,
            I => \this_vga_signals.un1_M_haddress_q_cry_8\
        );

    \I__1434\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9875\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__9875\,
            I => \N__9871\
        );

    \I__1432\ : InMux
    port map (
            O => \N__9874\,
            I => \N__9868\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__9871\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_3_1\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__9868\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_3_1\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__9863\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_1_0_cascade_\
        );

    \I__1428\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9857\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__9857\,
            I => \this_vga_signals.if_N_4_i\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__9854\,
            I => \this_vga_signals_un6_address_if_N_5_mux_0_cascade_\
        );

    \I__1425\ : CascadeMux
    port map (
            O => \N__9851\,
            I => \this_vga_signals.mult1_un47_sum_c3_cascade_\
        );

    \I__1424\ : InMux
    port map (
            O => \N__9848\,
            I => \N__9845\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__9845\,
            I => \this_vga_signals.if_m1_1\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__9842\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0_cascade_\
        );

    \I__1421\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9836\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__9836\,
            I => \this_vga_signals.if_m1_9_1\
        );

    \I__1419\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9828\
        );

    \I__1418\ : InMux
    port map (
            O => \N__9832\,
            I => \N__9825\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__9831\,
            I => \N__9820\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__9828\,
            I => \N__9817\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__9825\,
            I => \N__9813\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__9824\,
            I => \N__9810\
        );

    \I__1413\ : InMux
    port map (
            O => \N__9823\,
            I => \N__9807\
        );

    \I__1412\ : InMux
    port map (
            O => \N__9820\,
            I => \N__9804\
        );

    \I__1411\ : Sp12to4
    port map (
            O => \N__9817\,
            I => \N__9801\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__9816\,
            I => \N__9798\
        );

    \I__1409\ : Span4Mux_v
    port map (
            O => \N__9813\,
            I => \N__9795\
        );

    \I__1408\ : InMux
    port map (
            O => \N__9810\,
            I => \N__9792\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__9807\,
            I => \N__9787\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__9804\,
            I => \N__9787\
        );

    \I__1405\ : Span12Mux_v
    port map (
            O => \N__9801\,
            I => \N__9784\
        );

    \I__1404\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9781\
        );

    \I__1403\ : Span4Mux_h
    port map (
            O => \N__9795\,
            I => \N__9774\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__9792\,
            I => \N__9774\
        );

    \I__1401\ : Span4Mux_h
    port map (
            O => \N__9787\,
            I => \N__9774\
        );

    \I__1400\ : Odrv12
    port map (
            O => \N__9784\,
            I => \this_vga_signals.M_hstate_qZ0Z_1\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__9781\,
            I => \this_vga_signals.M_hstate_qZ0Z_1\
        );

    \I__1398\ : Odrv4
    port map (
            O => \N__9774\,
            I => \this_vga_signals.M_hstate_qZ0Z_1\
        );

    \I__1397\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9764\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__9764\,
            I => \this_vga_signals.M_haddress_qZ0Z_0\
        );

    \I__1395\ : InMux
    port map (
            O => \N__9761\,
            I => \N__9758\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__9758\,
            I => \this_vga_signals.M_haddress_qZ0Z_1\
        );

    \I__1393\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9752\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__9752\,
            I => \this_vga_signals.if_m2_0_1\
        );

    \I__1391\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9746\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__9746\,
            I => \this_vga_signals.if_N_3_0_i\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__9743\,
            I => \this_vga_signals.if_N_3_0_i_cascade_\
        );

    \I__1388\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9737\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__9737\,
            I => \this_vga_signals.mult1_un75_sum_c3_0\
        );

    \I__1386\ : InMux
    port map (
            O => \N__9734\,
            I => \N__9731\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__9731\,
            I => \this_vga_signals.if_i1_mux_0\
        );

    \I__1384\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9725\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__9725\,
            I => \this_vga_signals.if_m2\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__9722\,
            I => \this_vga_signals.M_haddress_q_RNILVKM8Z0Z_6_cascade_\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__9719\,
            I => \this_vga_signals.mult1_un54_sum_c3_cascade_\
        );

    \I__1380\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9713\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__9713\,
            I => \this_vga_signals.if_N_8_i\
        );

    \I__1378\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9707\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__9707\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_1_0\
        );

    \I__1376\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9701\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__9701\,
            I => \N__9698\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__9698\,
            I => \this_vga_signals.g1_2_1\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__9695\,
            I => \N__9692\
        );

    \I__1372\ : InMux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__9689\,
            I => \N__9686\
        );

    \I__1370\ : Odrv4
    port map (
            O => \N__9686\,
            I => \this_vga_signals.g2_5_0\
        );

    \I__1369\ : InMux
    port map (
            O => \N__9683\,
            I => \N__9680\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__9680\,
            I => \this_vga_signals.M_vaddress_q_RNI85LKP4Z0Z_2\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__9677\,
            I => \this_vga_signals.mult1_un54_sum_axb1_1_0_cascade_\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__9674\,
            I => \this_vga_signals.mult1_un61_sum_c3_1_1_0_cascade_\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__9671\,
            I => \this_vga_signals.g3_0_0_0_1_cascade_\
        );

    \I__1364\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9665\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__9665\,
            I => \this_vga_signals.g1_2\
        );

    \I__1362\ : InMux
    port map (
            O => \N__9662\,
            I => \N__9659\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__9659\,
            I => \this_vga_signals.g2\
        );

    \I__1360\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9653\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__9653\,
            I => \this_vga_signals.g1_0_1_0_0\
        );

    \I__1358\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9647\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__9647\,
            I => \this_vga_signals.N_4_i\
        );

    \I__1356\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__9641\,
            I => \this_vga_signals.g0_14_N_7L14_1\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__9638\,
            I => \this_vga_signals.g2_3_0_cascade_\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__9635\,
            I => \this_vga_signals.if_N_2_4_cascade_\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__9632\,
            I => \this_vga_signals.mult1_un61_sum_c3_2_cascade_\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__9629\,
            I => \this_vga_signals.g0_0_6_cascade_\
        );

    \I__1350\ : InMux
    port map (
            O => \N__9626\,
            I => \N__9623\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__9623\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3\
        );

    \I__1348\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9617\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__9617\,
            I => \this_vga_signals.g0_1_0\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__9614\,
            I => \this_vga_signals.mult1_un61_sum_c3_cascade_\
        );

    \I__1345\ : InMux
    port map (
            O => \N__9611\,
            I => \N__9608\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__9608\,
            I => \this_vga_signals.mult1_un68_sum_axb2_i\
        );

    \I__1343\ : CascadeMux
    port map (
            O => \N__9605\,
            I => \N__9602\
        );

    \I__1342\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9599\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__9599\,
            I => \this_vga_signals.g0_14_N_4L6\
        );

    \I__1340\ : InMux
    port map (
            O => \N__9596\,
            I => \N__9591\
        );

    \I__1339\ : InMux
    port map (
            O => \N__9595\,
            I => \N__9588\
        );

    \I__1338\ : InMux
    port map (
            O => \N__9594\,
            I => \N__9585\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__9591\,
            I => \N__9582\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__9588\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__9585\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1334\ : Odrv4
    port map (
            O => \N__9582\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1333\ : InMux
    port map (
            O => \N__9575\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__1332\ : InMux
    port map (
            O => \N__9572\,
            I => \N__9567\
        );

    \I__1331\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9564\
        );

    \I__1330\ : InMux
    port map (
            O => \N__9570\,
            I => \N__9561\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__9567\,
            I => \N__9558\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__9564\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__9561\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1326\ : Odrv4
    port map (
            O => \N__9558\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1325\ : InMux
    port map (
            O => \N__9551\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__1324\ : InMux
    port map (
            O => \N__9548\,
            I => \N__9542\
        );

    \I__1323\ : InMux
    port map (
            O => \N__9547\,
            I => \N__9537\
        );

    \I__1322\ : InMux
    port map (
            O => \N__9546\,
            I => \N__9537\
        );

    \I__1321\ : InMux
    port map (
            O => \N__9545\,
            I => \N__9534\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__9542\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__9537\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__9534\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1317\ : InMux
    port map (
            O => \N__9527\,
            I => \bfn_17_18_0_\
        );

    \I__1316\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9517\
        );

    \I__1315\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9512\
        );

    \I__1314\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9512\
        );

    \I__1313\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9507\
        );

    \I__1312\ : InMux
    port map (
            O => \N__9520\,
            I => \N__9507\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__9517\,
            I => \N__9499\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__9512\,
            I => \N__9499\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__9507\,
            I => \N__9499\
        );

    \I__1308\ : InMux
    port map (
            O => \N__9506\,
            I => \N__9496\
        );

    \I__1307\ : Span4Mux_v
    port map (
            O => \N__9499\,
            I => \N__9493\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__9496\,
            I => \this_vga_signals.M_hcounter_qZ0Z_10\
        );

    \I__1305\ : Odrv4
    port map (
            O => \N__9493\,
            I => \this_vga_signals.M_hcounter_qZ0Z_10\
        );

    \I__1304\ : InMux
    port map (
            O => \N__9488\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_9\
        );

    \I__1303\ : InMux
    port map (
            O => \N__9485\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_10\
        );

    \I__1302\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9477\
        );

    \I__1301\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9472\
        );

    \I__1300\ : InMux
    port map (
            O => \N__9480\,
            I => \N__9472\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__9477\,
            I => \this_vga_signals.M_hcounter_qZ0Z_11\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__9472\,
            I => \this_vga_signals.M_hcounter_qZ0Z_11\
        );

    \I__1297\ : InMux
    port map (
            O => \N__9467\,
            I => \N__9464\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__9464\,
            I => \this_vga_signals.g1_1_1\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__9461\,
            I => \this_vga_signals.g2_1_0_cascade_\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__9458\,
            I => \this_vga_signals.mult1_un40_sum_0_ac0_3_0_a1_0_cascade_\
        );

    \I__1293\ : InMux
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__9452\,
            I => \this_vga_signals.if_m3_0_0\
        );

    \I__1291\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__9446\,
            I => \this_vga_signals.mult1_un40_sum_0_ac0_3_1\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__9443\,
            I => \this_vga_signals.mult1_un40_sum_0_ac0_3_0_cascade_\
        );

    \I__1288\ : InMux
    port map (
            O => \N__9440\,
            I => \N__9437\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__9437\,
            I => \this_vga_signals.mult1_un40_sum_0_ac0_3_2\
        );

    \I__1286\ : InMux
    port map (
            O => \N__9434\,
            I => \N__9431\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__1284\ : Odrv4
    port map (
            O => \N__9428\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_14\
        );

    \I__1283\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9422\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__9422\,
            I => \N__9419\
        );

    \I__1281\ : Span4Mux_v
    port map (
            O => \N__9419\,
            I => \N__9416\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__9416\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_15\
        );

    \I__1279\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9404\
        );

    \I__1278\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9404\
        );

    \I__1277\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9401\
        );

    \I__1276\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9396\
        );

    \I__1275\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9396\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__9404\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__9401\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__9396\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__9389\,
            I => \N__9386\
        );

    \I__1270\ : InMux
    port map (
            O => \N__9386\,
            I => \N__9382\
        );

    \I__1269\ : InMux
    port map (
            O => \N__9385\,
            I => \N__9378\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__9382\,
            I => \N__9375\
        );

    \I__1267\ : InMux
    port map (
            O => \N__9381\,
            I => \N__9372\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__9378\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__9375\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__9372\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1263\ : InMux
    port map (
            O => \N__9365\,
            I => \N__9361\
        );

    \I__1262\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9358\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__9361\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__9358\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1259\ : InMux
    port map (
            O => \N__9353\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__1258\ : InMux
    port map (
            O => \N__9350\,
            I => \N__9346\
        );

    \I__1257\ : InMux
    port map (
            O => \N__9349\,
            I => \N__9343\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__9346\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__9343\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1254\ : InMux
    port map (
            O => \N__9338\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__9335\,
            I => \N__9331\
        );

    \I__1252\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9328\
        );

    \I__1251\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9325\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__9328\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__9325\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1248\ : InMux
    port map (
            O => \N__9320\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__1247\ : InMux
    port map (
            O => \N__9317\,
            I => \N__9312\
        );

    \I__1246\ : InMux
    port map (
            O => \N__9316\,
            I => \N__9309\
        );

    \I__1245\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9306\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__9312\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__9309\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__9306\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9299\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__1240\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9290\
        );

    \I__1239\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9283\
        );

    \I__1238\ : InMux
    port map (
            O => \N__9294\,
            I => \N__9283\
        );

    \I__1237\ : InMux
    port map (
            O => \N__9293\,
            I => \N__9283\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__9290\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__9283\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1234\ : InMux
    port map (
            O => \N__9278\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__1233\ : InMux
    port map (
            O => \N__9275\,
            I => \N__9272\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__9272\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_13\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__9269\,
            I => \this_vga_signals.mult1_un40_sum_0_ac0_3_2_1_cascade_\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__9266\,
            I => \this_vga_signals.if_N_2_6_cascade_\
        );

    \I__1229\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__9260\,
            I => \this_vga_signals.mult1_un61_sum_c3_0\
        );

    \I__1227\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__9254\,
            I => \this_vga_signals.g0_14_N_7L14\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__9251\,
            I => \this_vga_signals.if_N_9_0_cascade_\
        );

    \I__1224\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9245\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__9245\,
            I => \this_vga_signals.mult1_un61_sum_axb1\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__9242\,
            I => \this_vga_signals.mult1_un61_sum_axb1_cascade_\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__9239\,
            I => \this_vga_signals.if_m3_1_2_cascade_\
        );

    \I__1220\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9233\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__9233\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3_out\
        );

    \I__1218\ : InMux
    port map (
            O => \N__9230\,
            I => \N__9227\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__9227\,
            I => \this_vga_signals.if_i2_mux_0\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__9224\,
            I => \this_vga_signals.if_N_6_0_0_cascade_\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__9221\,
            I => \N__9218\
        );

    \I__1214\ : CascadeBuf
    port map (
            O => \N__9218\,
            I => \N__9215\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__9215\,
            I => \N__9212\
        );

    \I__1212\ : CascadeBuf
    port map (
            O => \N__9212\,
            I => \N__9209\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__9209\,
            I => \N__9206\
        );

    \I__1210\ : CascadeBuf
    port map (
            O => \N__9206\,
            I => \N__9203\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__1208\ : CascadeBuf
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__1206\ : CascadeBuf
    port map (
            O => \N__9194\,
            I => \N__9191\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__9191\,
            I => \N__9188\
        );

    \I__1204\ : CascadeBuf
    port map (
            O => \N__9188\,
            I => \N__9185\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__9185\,
            I => \N__9182\
        );

    \I__1202\ : CascadeBuf
    port map (
            O => \N__9182\,
            I => \N__9179\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__9179\,
            I => \N__9176\
        );

    \I__1200\ : CascadeBuf
    port map (
            O => \N__9176\,
            I => \N__9173\
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__9173\,
            I => \N__9170\
        );

    \I__1198\ : CascadeBuf
    port map (
            O => \N__9170\,
            I => \N__9167\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__9167\,
            I => \N__9164\
        );

    \I__1196\ : CascadeBuf
    port map (
            O => \N__9164\,
            I => \N__9161\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__9161\,
            I => \N__9158\
        );

    \I__1194\ : CascadeBuf
    port map (
            O => \N__9158\,
            I => \N__9155\
        );

    \I__1193\ : CascadeMux
    port map (
            O => \N__9155\,
            I => \N__9152\
        );

    \I__1192\ : CascadeBuf
    port map (
            O => \N__9152\,
            I => \N__9149\
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__9149\,
            I => \N__9146\
        );

    \I__1190\ : CascadeBuf
    port map (
            O => \N__9146\,
            I => \N__9143\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__9143\,
            I => \N__9140\
        );

    \I__1188\ : CascadeBuf
    port map (
            O => \N__9140\,
            I => \N__9137\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__9137\,
            I => \N__9134\
        );

    \I__1186\ : CascadeBuf
    port map (
            O => \N__9134\,
            I => \N__9131\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__1184\ : InMux
    port map (
            O => \N__9128\,
            I => \N__9125\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__9125\,
            I => \N__9122\
        );

    \I__1182\ : Span12Mux_h
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__1181\ : Span12Mux_v
    port map (
            O => \N__9119\,
            I => \N__9116\
        );

    \I__1180\ : Odrv12
    port map (
            O => \N__9116\,
            I => this_vga_signals_un6_address_if_generate_plus_mult1_un75_sum_i_3
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__9113\,
            I => \this_vga_signals.g2_2_cascade_\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__9110\,
            I => \this_vga_signals.g1_cascade_\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__9107\,
            I => \this_vga_signals.g2_5_cascade_\
        );

    \I__1176\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9101\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__9101\,
            I => \this_vga_signals.g1_1_4\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__9098\,
            I => \this_vga_signals.g0_14_N_8L16_cascade_\
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__9095\,
            I => \this_vga_signals.mult1_un75_sum_c3_0_0_cascade_\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__9092\,
            I => \N__9089\
        );

    \I__1171\ : CascadeBuf
    port map (
            O => \N__9089\,
            I => \N__9086\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__1169\ : CascadeBuf
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__1167\ : CascadeBuf
    port map (
            O => \N__9077\,
            I => \N__9074\
        );

    \I__1166\ : CascadeMux
    port map (
            O => \N__9074\,
            I => \N__9071\
        );

    \I__1165\ : CascadeBuf
    port map (
            O => \N__9071\,
            I => \N__9068\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__9068\,
            I => \N__9065\
        );

    \I__1163\ : CascadeBuf
    port map (
            O => \N__9065\,
            I => \N__9062\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__1161\ : CascadeBuf
    port map (
            O => \N__9059\,
            I => \N__9056\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__9056\,
            I => \N__9053\
        );

    \I__1159\ : CascadeBuf
    port map (
            O => \N__9053\,
            I => \N__9050\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__1157\ : CascadeBuf
    port map (
            O => \N__9047\,
            I => \N__9044\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__1155\ : CascadeBuf
    port map (
            O => \N__9041\,
            I => \N__9038\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__1153\ : CascadeBuf
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__1152\ : CascadeMux
    port map (
            O => \N__9032\,
            I => \N__9029\
        );

    \I__1151\ : CascadeBuf
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__9026\,
            I => \N__9023\
        );

    \I__1149\ : CascadeBuf
    port map (
            O => \N__9023\,
            I => \N__9020\
        );

    \I__1148\ : CascadeMux
    port map (
            O => \N__9020\,
            I => \N__9017\
        );

    \I__1147\ : CascadeBuf
    port map (
            O => \N__9017\,
            I => \N__9014\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__9014\,
            I => \N__9011\
        );

    \I__1145\ : CascadeBuf
    port map (
            O => \N__9011\,
            I => \N__9008\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__9008\,
            I => \N__9005\
        );

    \I__1143\ : CascadeBuf
    port map (
            O => \N__9005\,
            I => \N__9002\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__1141\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8996\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__8996\,
            I => \N__8993\
        );

    \I__1139\ : Span4Mux_v
    port map (
            O => \N__8993\,
            I => \N__8990\
        );

    \I__1138\ : Span4Mux_h
    port map (
            O => \N__8990\,
            I => \N__8987\
        );

    \I__1137\ : Span4Mux_h
    port map (
            O => \N__8987\,
            I => \N__8984\
        );

    \I__1136\ : Sp12to4
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__1135\ : Span12Mux_s11_v
    port map (
            O => \N__8981\,
            I => \N__8978\
        );

    \I__1134\ : Odrv12
    port map (
            O => \N__8978\,
            I => this_vga_signals_un14_address_if_generate_plus_mult1_un75_sum_i_3
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__8975\,
            I => \this_vga_signals.N_386_0_cascade_\
        );

    \I__1132\ : InMux
    port map (
            O => \N__8972\,
            I => \N__8968\
        );

    \I__1131\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8965\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__8968\,
            I => \N__8960\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__8965\,
            I => \N__8960\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__8960\,
            I => \this_vga_signals.M_hstate_q_srsts_0_o3_2_1\
        );

    \I__1127\ : InMux
    port map (
            O => \N__8957\,
            I => \N__8952\
        );

    \I__1126\ : InMux
    port map (
            O => \N__8956\,
            I => \N__8949\
        );

    \I__1125\ : InMux
    port map (
            O => \N__8955\,
            I => \N__8946\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__8952\,
            I => \this_vga_signals.N_388_0\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__8949\,
            I => \this_vga_signals.N_388_0\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__8946\,
            I => \this_vga_signals.N_388_0\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__1120\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8933\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__8933\,
            I => \this_vga_signals.M_hstate_q_srsts_0_o3_2_3_5\
        );

    \I__1118\ : InMux
    port map (
            O => \N__8930\,
            I => \N__8925\
        );

    \I__1117\ : InMux
    port map (
            O => \N__8929\,
            I => \N__8920\
        );

    \I__1116\ : InMux
    port map (
            O => \N__8928\,
            I => \N__8920\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__8925\,
            I => \this_vga_signals.N_393_0\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__8920\,
            I => \this_vga_signals.N_393_0\
        );

    \I__1113\ : InMux
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__8912\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__1111\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8897\
        );

    \I__1110\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8897\
        );

    \I__1109\ : InMux
    port map (
            O => \N__8907\,
            I => \N__8897\
        );

    \I__1108\ : InMux
    port map (
            O => \N__8906\,
            I => \N__8897\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__8897\,
            I => \N__8894\
        );

    \I__1106\ : Odrv12
    port map (
            O => \N__8894\,
            I => rst_n_c
        );

    \I__1105\ : InMux
    port map (
            O => \N__8891\,
            I => \N__8888\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__8888\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__1103\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8882\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__8882\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__8879\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa_cascade_\
        );

    \I__1100\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8873\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__8873\,
            I => \this_vga_signals.N_405_0\
        );

    \I__1098\ : InMux
    port map (
            O => \N__8870\,
            I => \N__8864\
        );

    \I__1097\ : InMux
    port map (
            O => \N__8869\,
            I => \N__8864\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__8864\,
            I => \this_vga_signals.M_hstate_qZ0Z_0\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__8861\,
            I => \this_vga_signals.N_405_0_cascade_\
        );

    \I__1094\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8855\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__8855\,
            I => \this_vga_signals.N_409\
        );

    \I__1092\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8847\
        );

    \I__1091\ : InMux
    port map (
            O => \N__8851\,
            I => \N__8842\
        );

    \I__1090\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8842\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__8847\,
            I => \this_vga_signals.N_397_0\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__8842\,
            I => \this_vga_signals.N_397_0\
        );

    \I__1087\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8832\
        );

    \I__1086\ : InMux
    port map (
            O => \N__8836\,
            I => \N__8829\
        );

    \I__1085\ : InMux
    port map (
            O => \N__8835\,
            I => \N__8826\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__8832\,
            I => \this_vga_signals.M_hstate_qZ0Z_5\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__8829\,
            I => \this_vga_signals.M_hstate_qZ0Z_5\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__8826\,
            I => \this_vga_signals.M_hstate_qZ0Z_5\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__8819\,
            I => \this_vga_signals.M_hstate_q_srsts_0_o3_2_3_5_cascade_\
        );

    \I__1080\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8810\
        );

    \I__1079\ : InMux
    port map (
            O => \N__8815\,
            I => \N__8810\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__8810\,
            I => \this_vga_signals.N_385_0\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__8807\,
            I => \this_vga_signals.N_385_0_cascade_\
        );

    \I__1076\ : InMux
    port map (
            O => \N__8804\,
            I => \N__8801\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__8801\,
            I => \N__8795\
        );

    \I__1074\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8792\
        );

    \I__1073\ : InMux
    port map (
            O => \N__8799\,
            I => \N__8787\
        );

    \I__1072\ : InMux
    port map (
            O => \N__8798\,
            I => \N__8787\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__8795\,
            I => \this_vga_signals.N_391_0\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__8792\,
            I => \this_vga_signals.N_391_0\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__8787\,
            I => \this_vga_signals.N_391_0\
        );

    \I__1068\ : InMux
    port map (
            O => \N__8780\,
            I => \N__8775\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__8779\,
            I => \N__8771\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__8778\,
            I => \N__8768\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__8775\,
            I => \N__8765\
        );

    \I__1064\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8762\
        );

    \I__1063\ : InMux
    port map (
            O => \N__8771\,
            I => \N__8759\
        );

    \I__1062\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8756\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__8765\,
            I => \this_vga_signals.N_386_0\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__8762\,
            I => \this_vga_signals.N_386_0\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__8759\,
            I => \this_vga_signals.N_386_0\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__8756\,
            I => \this_vga_signals.N_386_0\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__8747\,
            I => \this_vga_signals.N_390_0_cascade_\
        );

    \I__1056\ : InMux
    port map (
            O => \N__8744\,
            I => \N__8738\
        );

    \I__1055\ : InMux
    port map (
            O => \N__8743\,
            I => \N__8738\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__8738\,
            I => \this_vga_signals.N_390_0\
        );

    \I__1053\ : InMux
    port map (
            O => \N__8735\,
            I => \N__8731\
        );

    \I__1052\ : InMux
    port map (
            O => \N__8734\,
            I => \N__8728\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__8731\,
            I => \this_vga_signals.M_hstate_qZ0Z_2\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__8728\,
            I => \this_vga_signals.M_hstate_qZ0Z_2\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__8723\,
            I => \this_vga_signals.N_413_cascade_\
        );

    \I__1048\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8716\
        );

    \I__1047\ : InMux
    port map (
            O => \N__8719\,
            I => \N__8713\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__8716\,
            I => \this_vga_signals.N_398_0\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__8713\,
            I => \this_vga_signals.N_398_0\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__8708\,
            I => \N__8704\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__8707\,
            I => \N__8701\
        );

    \I__1042\ : InMux
    port map (
            O => \N__8704\,
            I => \N__8696\
        );

    \I__1041\ : InMux
    port map (
            O => \N__8701\,
            I => \N__8696\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__8696\,
            I => \this_vga_signals.M_hstate_qZ0Z_3\
        );

    \I__1039\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__8690\,
            I => \N__8687\
        );

    \I__1037\ : Odrv4
    port map (
            O => \N__8687\,
            I => \this_vga_signals.M_hstate_q_srsts_0_a3_0_4\
        );

    \I__1036\ : InMux
    port map (
            O => \N__8684\,
            I => \N__8681\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__8681\,
            I => \this_vga_signals.N_416\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__8678\,
            I => \this_vga_signals.M_hstate_q_srsts_0_a3_0_4_cascade_\
        );

    \I__1033\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__1031\ : Span4Mux_v
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__1030\ : Span4Mux_h
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__1029\ : Span4Mux_v
    port map (
            O => \N__8663\,
            I => \N__8659\
        );

    \I__1028\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8656\
        );

    \I__1027\ : Odrv4
    port map (
            O => \N__8659\,
            I => \this_vga_signals.M_hstate_qZ0Z_4\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__8656\,
            I => \this_vga_signals.M_hstate_qZ0Z_4\
        );

    \I__1025\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8648\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__8648\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_12\
        );

    \I__1023\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__8642\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_11\
        );

    \I__1021\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8636\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__8636\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_8\
        );

    \I__1019\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8630\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__8630\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_9\
        );

    \I__1017\ : InMux
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__8624\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_14\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__8621\,
            I => \this_vga_signals.N_417_cascade_\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__8618\,
            I => \this_vga_signals.N_412_cascade_\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__8615\,
            I => \N__8609\
        );

    \I__1012\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8606\
        );

    \I__1011\ : InMux
    port map (
            O => \N__8613\,
            I => \N__8603\
        );

    \I__1010\ : InMux
    port map (
            O => \N__8612\,
            I => \N__8600\
        );

    \I__1009\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8597\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__8606\,
            I => \N__8592\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__8603\,
            I => \N__8592\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__8600\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__8597\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1004\ : Odrv4
    port map (
            O => \N__8592\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1003\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8578\
        );

    \I__1002\ : InMux
    port map (
            O => \N__8584\,
            I => \N__8573\
        );

    \I__1001\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8573\
        );

    \I__1000\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8570\
        );

    \I__999\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8567\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__8578\,
            I => \N__8564\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__8573\,
            I => \N__8559\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__8570\,
            I => \N__8559\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__8567\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__8564\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__8559\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__992\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8548\
        );

    \I__991\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8545\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__8548\,
            I => \this_vga_signals.N_230_0\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__8545\,
            I => \this_vga_signals.N_230_0\
        );

    \I__988\ : CascadeMux
    port map (
            O => \N__8540\,
            I => \this_vga_signals.M_vstate_q_srsts_0_o2_2_5_cascade_\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__8537\,
            I => \N__8531\
        );

    \I__986\ : InMux
    port map (
            O => \N__8536\,
            I => \N__8527\
        );

    \I__985\ : InMux
    port map (
            O => \N__8535\,
            I => \N__8524\
        );

    \I__984\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8517\
        );

    \I__983\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8517\
        );

    \I__982\ : InMux
    port map (
            O => \N__8530\,
            I => \N__8517\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__8527\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__8524\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__8517\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__978\ : InMux
    port map (
            O => \N__8510\,
            I => \N__8503\
        );

    \I__977\ : InMux
    port map (
            O => \N__8509\,
            I => \N__8493\
        );

    \I__976\ : InMux
    port map (
            O => \N__8508\,
            I => \N__8493\
        );

    \I__975\ : InMux
    port map (
            O => \N__8507\,
            I => \N__8493\
        );

    \I__974\ : InMux
    port map (
            O => \N__8506\,
            I => \N__8493\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__8503\,
            I => \N__8490\
        );

    \I__972\ : InMux
    port map (
            O => \N__8502\,
            I => \N__8487\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__8493\,
            I => \this_vga_signals.N_248_0\
        );

    \I__970\ : Odrv4
    port map (
            O => \N__8490\,
            I => \this_vga_signals.N_248_0\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__8487\,
            I => \this_vga_signals.N_248_0\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__8480\,
            I => \this_vga_signals.N_248_0_cascade_\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__8477\,
            I => \N__8473\
        );

    \I__966\ : InMux
    port map (
            O => \N__8476\,
            I => \N__8467\
        );

    \I__965\ : InMux
    port map (
            O => \N__8473\,
            I => \N__8464\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__8472\,
            I => \N__8461\
        );

    \I__963\ : CascadeMux
    port map (
            O => \N__8471\,
            I => \N__8458\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__8470\,
            I => \N__8455\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__8467\,
            I => \N__8450\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__8464\,
            I => \N__8447\
        );

    \I__959\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8440\
        );

    \I__958\ : InMux
    port map (
            O => \N__8458\,
            I => \N__8440\
        );

    \I__957\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8440\
        );

    \I__956\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8437\
        );

    \I__955\ : InMux
    port map (
            O => \N__8453\,
            I => \N__8434\
        );

    \I__954\ : Odrv4
    port map (
            O => \N__8450\,
            I => \this_vga_signals.M_vstate_qZ0Z_5\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__8447\,
            I => \this_vga_signals.M_vstate_qZ0Z_5\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__8440\,
            I => \this_vga_signals.M_vstate_qZ0Z_5\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__8437\,
            I => \this_vga_signals.M_vstate_qZ0Z_5\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__8434\,
            I => \this_vga_signals.M_vstate_qZ0Z_5\
        );

    \I__949\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8420\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__8420\,
            I => \this_vga_signals.N_252\
        );

    \I__947\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8412\
        );

    \I__946\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8409\
        );

    \I__945\ : InMux
    port map (
            O => \N__8415\,
            I => \N__8403\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__8412\,
            I => \N__8398\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__8409\,
            I => \N__8398\
        );

    \I__942\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8395\
        );

    \I__941\ : InMux
    port map (
            O => \N__8407\,
            I => \N__8392\
        );

    \I__940\ : InMux
    port map (
            O => \N__8406\,
            I => \N__8389\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__8403\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__938\ : Odrv4
    port map (
            O => \N__8398\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__8395\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__8392\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__8389\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__8378\,
            I => \N__8373\
        );

    \I__933\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8368\
        );

    \I__932\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8365\
        );

    \I__931\ : InMux
    port map (
            O => \N__8373\,
            I => \N__8362\
        );

    \I__930\ : InMux
    port map (
            O => \N__8372\,
            I => \N__8359\
        );

    \I__929\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8356\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__8368\,
            I => \N__8353\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__8365\,
            I => \N__8350\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__8362\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__8359\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__8356\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__8353\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__8350\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__8339\,
            I => \N__8335\
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__8338\,
            I => \N__8332\
        );

    \I__919\ : InMux
    port map (
            O => \N__8335\,
            I => \N__8326\
        );

    \I__918\ : InMux
    port map (
            O => \N__8332\,
            I => \N__8323\
        );

    \I__917\ : InMux
    port map (
            O => \N__8331\,
            I => \N__8320\
        );

    \I__916\ : InMux
    port map (
            O => \N__8330\,
            I => \N__8317\
        );

    \I__915\ : InMux
    port map (
            O => \N__8329\,
            I => \N__8314\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__8326\,
            I => \N__8309\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__8323\,
            I => \N__8309\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__8320\,
            I => \N__8304\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__8317\,
            I => \N__8304\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__8314\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__8309\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__8304\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__907\ : InMux
    port map (
            O => \N__8297\,
            I => \N__8291\
        );

    \I__906\ : InMux
    port map (
            O => \N__8296\,
            I => \N__8287\
        );

    \I__905\ : InMux
    port map (
            O => \N__8295\,
            I => \N__8284\
        );

    \I__904\ : InMux
    port map (
            O => \N__8294\,
            I => \N__8281\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__8291\,
            I => \N__8278\
        );

    \I__902\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8275\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__8287\,
            I => \N__8272\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__8284\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__8281\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__898\ : Odrv4
    port map (
            O => \N__8278\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__8275\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__896\ : Odrv4
    port map (
            O => \N__8272\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__8261\,
            I => \this_vga_signals.M_vstate_q_srsts_0_o2_2_3_cascade_\
        );

    \I__894\ : InMux
    port map (
            O => \N__8258\,
            I => \N__8255\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__8255\,
            I => \N__8252\
        );

    \I__892\ : Odrv4
    port map (
            O => \N__8252\,
            I => \this_vga_signals.N_255\
        );

    \I__891\ : InMux
    port map (
            O => \N__8249\,
            I => \N__8246\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__8246\,
            I => \this_vga_signals.M_vstate_q_srsts_0_o2_2_3\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__8243\,
            I => \N__8239\
        );

    \I__888\ : InMux
    port map (
            O => \N__8242\,
            I => \N__8234\
        );

    \I__887\ : InMux
    port map (
            O => \N__8239\,
            I => \N__8234\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__8234\,
            I => \this_vga_signals.M_vstate_qZ0Z_3\
        );

    \I__885\ : InMux
    port map (
            O => \N__8231\,
            I => \N__8222\
        );

    \I__884\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8222\
        );

    \I__883\ : InMux
    port map (
            O => \N__8229\,
            I => \N__8217\
        );

    \I__882\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8217\
        );

    \I__881\ : InMux
    port map (
            O => \N__8227\,
            I => \N__8214\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__8222\,
            I => \this_vga_signals.N_226_0\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__8217\,
            I => \this_vga_signals.N_226_0\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__8214\,
            I => \this_vga_signals.N_226_0\
        );

    \I__877\ : InMux
    port map (
            O => \N__8207\,
            I => \N__8204\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__8204\,
            I => \this_vga_signals.N_256\
        );

    \I__875\ : InMux
    port map (
            O => \N__8201\,
            I => \N__8198\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__8198\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_7\
        );

    \I__873\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8192\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__8192\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_10\
        );

    \I__871\ : IoInMux
    port map (
            O => \N__8189\,
            I => \N__8186\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__8186\,
            I => \N__8183\
        );

    \I__869\ : Span12Mux_s11_h
    port map (
            O => \N__8183\,
            I => \N__8180\
        );

    \I__868\ : Odrv12
    port map (
            O => \N__8180\,
            I => \this_vga_signals.M_vstate_q_RNI3M6M4Z0Z_0\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__8177\,
            I => \this_vga_signals.N_251_cascade_\
        );

    \I__866\ : InMux
    port map (
            O => \N__8174\,
            I => \N__8170\
        );

    \I__865\ : InMux
    port map (
            O => \N__8173\,
            I => \N__8167\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__8170\,
            I => \N__8164\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__8167\,
            I => \this_vga_signals.N_237_0\
        );

    \I__862\ : Odrv4
    port map (
            O => \N__8164\,
            I => \this_vga_signals.N_237_0\
        );

    \I__861\ : InMux
    port map (
            O => \N__8159\,
            I => \N__8155\
        );

    \I__860\ : InMux
    port map (
            O => \N__8158\,
            I => \N__8151\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__8155\,
            I => \N__8148\
        );

    \I__858\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8145\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__8151\,
            I => \this_vga_signals.M_vstate_qZ0Z_0\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__8148\,
            I => \this_vga_signals.M_vstate_qZ0Z_0\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__8145\,
            I => \this_vga_signals.M_vstate_qZ0Z_0\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__8138\,
            I => \this_vga_signals.M_vstate_q_srsts_0_a4_0_4_cascade_\
        );

    \I__853\ : InMux
    port map (
            O => \N__8135\,
            I => \N__8132\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8132\,
            I => \this_vga_signals.M_vstate_q_srsts_0_a4_0_4\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__8129\,
            I => \this_vga_signals.N_230_0_cascade_\
        );

    \I__850\ : IoInMux
    port map (
            O => \N__8126\,
            I => \N__8123\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__8123\,
            I => \N__8120\
        );

    \I__848\ : IoSpan4Mux
    port map (
            O => \N__8120\,
            I => \N__8117\
        );

    \I__847\ : Span4Mux_s2_v
    port map (
            O => \N__8117\,
            I => \N__8114\
        );

    \I__846\ : Sp12to4
    port map (
            O => \N__8114\,
            I => \N__8110\
        );

    \I__845\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8107\
        );

    \I__844\ : Span12Mux_h
    port map (
            O => \N__8110\,
            I => \N__8104\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__8107\,
            I => \N__8101\
        );

    \I__842\ : Odrv12
    port map (
            O => \N__8104\,
            I => vsync_c
        );

    \I__841\ : Odrv4
    port map (
            O => \N__8101\,
            I => vsync_c
        );

    \I__840\ : InMux
    port map (
            O => \N__8096\,
            I => \N__8091\
        );

    \I__839\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8088\
        );

    \I__838\ : InMux
    port map (
            O => \N__8094\,
            I => \N__8085\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__8091\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__8088\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__8085\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__834\ : InMux
    port map (
            O => \N__8078\,
            I => \N__8073\
        );

    \I__833\ : InMux
    port map (
            O => \N__8077\,
            I => \N__8070\
        );

    \I__832\ : InMux
    port map (
            O => \N__8076\,
            I => \N__8067\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__8073\,
            I => \N__8064\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8070\,
            I => \N__8061\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__8067\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__828\ : Odrv4
    port map (
            O => \N__8064\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__827\ : Odrv4
    port map (
            O => \N__8061\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__8054\,
            I => \N__8050\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__8053\,
            I => \N__8046\
        );

    \I__824\ : InMux
    port map (
            O => \N__8050\,
            I => \N__8042\
        );

    \I__823\ : InMux
    port map (
            O => \N__8049\,
            I => \N__8037\
        );

    \I__822\ : InMux
    port map (
            O => \N__8046\,
            I => \N__8037\
        );

    \I__821\ : InMux
    port map (
            O => \N__8045\,
            I => \N__8034\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__8042\,
            I => \N__8031\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__8037\,
            I => \N__8028\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__8034\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__817\ : Odrv4
    port map (
            O => \N__8031\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__8028\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__815\ : InMux
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__813\ : Span4Mux_v
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__812\ : Odrv4
    port map (
            O => \N__8012\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_1\
        );

    \I__811\ : InMux
    port map (
            O => \N__8009\,
            I => \N__8006\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__8006\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_6\
        );

    \I__809\ : InMux
    port map (
            O => \N__8003\,
            I => \N__8000\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__8000\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_2\
        );

    \I__807\ : InMux
    port map (
            O => \N__7997\,
            I => \N__7994\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__7994\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_3\
        );

    \I__805\ : InMux
    port map (
            O => \N__7991\,
            I => \N__7988\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__7988\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_4\
        );

    \I__803\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7982\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__7982\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_5\
        );

    \I__801\ : InMux
    port map (
            O => \N__7979\,
            I => \N__7976\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__7976\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_13\
        );

    \I__799\ : InMux
    port map (
            O => \N__7973\,
            I => \N__7970\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__7970\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_11\
        );

    \I__797\ : InMux
    port map (
            O => \N__7967\,
            I => \N__7964\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__7964\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_12\
        );

    \I__795\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__7958\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_9\
        );

    \I__793\ : InMux
    port map (
            O => \N__7955\,
            I => \N__7952\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__7952\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_10\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__7949\,
            I => \this_vga_signals.N_237_0_cascade_\
        );

    \I__790\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7943\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__7943\,
            I => \this_vga_signals.M_vstate_d_0_sqmuxa\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__7940\,
            I => \N__7937\
        );

    \I__787\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7931\
        );

    \I__786\ : InMux
    port map (
            O => \N__7936\,
            I => \N__7931\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__7931\,
            I => \this_vga_signals.N_221_0\
        );

    \I__784\ : InMux
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__7925\,
            I => \this_vga_signals.N_225_0\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__7922\,
            I => \this_vga_signals.N_225_0_cascade_\
        );

    \I__781\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__7916\,
            I => \this_vga_signals.N_239_0\
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__7913\,
            I => \this_vga_signals.N_239_0_cascade_\
        );

    \I__778\ : IoInMux
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__7907\,
            I => \N__7904\
        );

    \I__776\ : Span4Mux_s0_h
    port map (
            O => \N__7904\,
            I => \N__7900\
        );

    \I__775\ : InMux
    port map (
            O => \N__7903\,
            I => \N__7897\
        );

    \I__774\ : Sp12to4
    port map (
            O => \N__7900\,
            I => \N__7894\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__7897\,
            I => \N__7891\
        );

    \I__772\ : Span12Mux_v
    port map (
            O => \N__7894\,
            I => \N__7887\
        );

    \I__771\ : Sp12to4
    port map (
            O => \N__7891\,
            I => \N__7884\
        );

    \I__770\ : InMux
    port map (
            O => \N__7890\,
            I => \N__7881\
        );

    \I__769\ : Span12Mux_h
    port map (
            O => \N__7887\,
            I => \N__7876\
        );

    \I__768\ : Span12Mux_v
    port map (
            O => \N__7884\,
            I => \N__7873\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__7881\,
            I => \N__7870\
        );

    \I__766\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7867\
        );

    \I__765\ : InMux
    port map (
            O => \N__7879\,
            I => \N__7864\
        );

    \I__764\ : Odrv12
    port map (
            O => \N__7876\,
            I => port_nmib_c
        );

    \I__763\ : Odrv12
    port map (
            O => \N__7873\,
            I => port_nmib_c
        );

    \I__762\ : Odrv4
    port map (
            O => \N__7870\,
            I => port_nmib_c
        );

    \I__761\ : LocalMux
    port map (
            O => \N__7867\,
            I => port_nmib_c
        );

    \I__760\ : LocalMux
    port map (
            O => \N__7864\,
            I => port_nmib_c
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__7853\,
            I => \this_vga_signals.N_258_cascade_\
        );

    \I__758\ : InMux
    port map (
            O => \N__7850\,
            I => \N__7847\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__7847\,
            I => \this_vga_signals.N_238_0\
        );

    \I__756\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7838\
        );

    \I__755\ : InMux
    port map (
            O => \N__7843\,
            I => \N__7838\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__7838\,
            I => \this_vga_signals.M_vstate_qZ0Z_2\
        );

    \I__753\ : InMux
    port map (
            O => \N__7835\,
            I => \bfn_13_18_0_\
        );

    \I__752\ : InMux
    port map (
            O => \N__7832\,
            I => \this_vga_signals.un1_M_vcounter_q_10_cry_8\
        );

    \I__751\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__7826\,
            I => \this_vga_signals.un1_M_vcounter_q_10_cry_2_THRU_CO\
        );

    \I__749\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7820\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__7820\,
            I => \this_vga_signals.un1_M_vcounter_q_10_cry_1_THRU_CO\
        );

    \I__747\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7814\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__7814\,
            I => \this_vga_signals.un1_M_vcounter_q_10_cry_0_THRU_CO\
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__7811\,
            I => \this_vga_signals.N_238_0_cascade_\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__7808\,
            I => \this_vga_signals.N_221_0_cascade_\
        );

    \I__743\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7799\
        );

    \I__742\ : InMux
    port map (
            O => \N__7804\,
            I => \N__7799\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__7799\,
            I => \this_vga_signals.N_232_0\
        );

    \I__740\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7793\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__7793\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_3\
        );

    \I__738\ : InMux
    port map (
            O => \N__7790\,
            I => \N__7787\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__7787\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_4\
        );

    \I__736\ : InMux
    port map (
            O => \N__7784\,
            I => \this_vga_signals.un1_M_vcounter_q_10_cry_0\
        );

    \I__735\ : InMux
    port map (
            O => \N__7781\,
            I => \this_vga_signals.un1_M_vcounter_q_10_cry_1\
        );

    \I__734\ : InMux
    port map (
            O => \N__7778\,
            I => \this_vga_signals.un1_M_vcounter_q_10_cry_2\
        );

    \I__733\ : InMux
    port map (
            O => \N__7775\,
            I => \this_vga_signals.un1_M_vcounter_q_10_cry_3\
        );

    \I__732\ : InMux
    port map (
            O => \N__7772\,
            I => \this_vga_signals.un1_M_vcounter_q_10_cry_4\
        );

    \I__731\ : InMux
    port map (
            O => \N__7769\,
            I => \this_vga_signals.un1_M_vcounter_q_10_cry_5\
        );

    \I__730\ : InMux
    port map (
            O => \N__7766\,
            I => \this_vga_signals.un1_M_vcounter_q_10_cry_6\
        );

    \I__729\ : InMux
    port map (
            O => \N__7763\,
            I => \N__7756\
        );

    \I__728\ : InMux
    port map (
            O => \N__7762\,
            I => \N__7756\
        );

    \I__727\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7753\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__7756\,
            I => \N__7748\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__7753\,
            I => \N__7748\
        );

    \I__724\ : Span4Mux_v
    port map (
            O => \N__7748\,
            I => \N__7745\
        );

    \I__723\ : Span4Mux_v
    port map (
            O => \N__7745\,
            I => \N__7742\
        );

    \I__722\ : Sp12to4
    port map (
            O => \N__7742\,
            I => \N__7739\
        );

    \I__721\ : Span12Mux_h
    port map (
            O => \N__7739\,
            I => \N__7736\
        );

    \I__720\ : Odrv12
    port map (
            O => \N__7736\,
            I => port_clk_c
        );

    \I__719\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7729\
        );

    \I__718\ : InMux
    port map (
            O => \N__7732\,
            I => \N__7726\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__7729\,
            I => \this_start_data_delay_this_edge_detector_M_last_q\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__7726\,
            I => \this_start_data_delay_this_edge_detector_M_last_q\
        );

    \I__715\ : InMux
    port map (
            O => \N__7721\,
            I => \N__7718\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__7718\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_0\
        );

    \I__713\ : InMux
    port map (
            O => \N__7715\,
            I => \N__7712\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__7712\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_1\
        );

    \I__711\ : InMux
    port map (
            O => \N__7709\,
            I => \N__7706\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__7706\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_2\
        );

    \I__709\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7700\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__7700\,
            I => m16
        );

    \I__707\ : InMux
    port map (
            O => \N__7697\,
            I => \N__7694\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__7694\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_8\
        );

    \I__705\ : InMux
    port map (
            O => \N__7691\,
            I => \N__7688\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__7688\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_6\
        );

    \I__703\ : InMux
    port map (
            O => \N__7685\,
            I => \N__7682\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__7682\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_7\
        );

    \I__701\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7676\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__7676\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_5\
        );

    \I__699\ : InMux
    port map (
            O => \N__7673\,
            I => \N__7670\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__7670\,
            I => \N__7667\
        );

    \I__697\ : Span4Mux_v
    port map (
            O => \N__7667\,
            I => \N__7664\
        );

    \I__696\ : Odrv4
    port map (
            O => \N__7664\,
            I => \rgb_2_5_0__i2_mux_0\
        );

    \I__695\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7658\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__7658\,
            I => \N__7655\
        );

    \I__693\ : Odrv12
    port map (
            O => \N__7655\,
            I => \rgb_2_5_0__i2_mux\
        );

    \I__692\ : InMux
    port map (
            O => \N__7652\,
            I => \N__7649\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__690\ : Span4Mux_v
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__7643\,
            I => m19
        );

    \I__688\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7634\
        );

    \I__687\ : InMux
    port map (
            O => \N__7639\,
            I => \N__7631\
        );

    \I__686\ : InMux
    port map (
            O => \N__7638\,
            I => \N__7628\
        );

    \I__685\ : InMux
    port map (
            O => \N__7637\,
            I => \N__7625\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__7634\,
            I => \N__7622\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__7631\,
            I => \N__7618\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__7628\,
            I => \N__7615\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__7625\,
            I => \N__7612\
        );

    \I__680\ : Span4Mux_v
    port map (
            O => \N__7622\,
            I => \N__7608\
        );

    \I__679\ : InMux
    port map (
            O => \N__7621\,
            I => \N__7605\
        );

    \I__678\ : Span4Mux_v
    port map (
            O => \N__7618\,
            I => \N__7600\
        );

    \I__677\ : Span4Mux_v
    port map (
            O => \N__7615\,
            I => \N__7600\
        );

    \I__676\ : Span4Mux_v
    port map (
            O => \N__7612\,
            I => \N__7597\
        );

    \I__675\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7594\
        );

    \I__674\ : Span4Mux_v
    port map (
            O => \N__7608\,
            I => \N__7589\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__7605\,
            I => \N__7589\
        );

    \I__672\ : Odrv4
    port map (
            O => \N__7600\,
            I => rgb72
        );

    \I__671\ : Odrv4
    port map (
            O => \N__7597\,
            I => rgb72
        );

    \I__670\ : LocalMux
    port map (
            O => \N__7594\,
            I => rgb72
        );

    \I__669\ : Odrv4
    port map (
            O => \N__7589\,
            I => rgb72
        );

    \I__668\ : IoInMux
    port map (
            O => \N__7580\,
            I => \N__7577\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__7577\,
            I => \N__7574\
        );

    \I__666\ : IoSpan4Mux
    port map (
            O => \N__7574\,
            I => \N__7571\
        );

    \I__665\ : Sp12to4
    port map (
            O => \N__7571\,
            I => \N__7568\
        );

    \I__664\ : Span12Mux_s6_h
    port map (
            O => \N__7568\,
            I => \N__7565\
        );

    \I__663\ : Odrv12
    port map (
            O => \N__7565\,
            I => rgb_c_3
        );

    \I__662\ : InMux
    port map (
            O => \N__7562\,
            I => \N__7559\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__7559\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_0\
        );

    \I__660\ : IoInMux
    port map (
            O => \N__7556\,
            I => \N__7553\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__7553\,
            I => \N__7550\
        );

    \I__658\ : Span4Mux_s1_v
    port map (
            O => \N__7550\,
            I => \N__7547\
        );

    \I__657\ : Span4Mux_v
    port map (
            O => \N__7547\,
            I => \N__7544\
        );

    \I__656\ : Span4Mux_v
    port map (
            O => \N__7544\,
            I => \N__7541\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__7541\,
            I => \this_vga_signals_M_hstate_q_i_1\
        );

    \I__654\ : IoInMux
    port map (
            O => \N__7538\,
            I => \N__7535\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__7535\,
            I => \N__7532\
        );

    \I__652\ : Span12Mux_s2_v
    port map (
            O => \N__7532\,
            I => \N__7529\
        );

    \I__651\ : Odrv12
    port map (
            O => \N__7529\,
            I => port_nmib_c_i
        );

    \I__650\ : IoInMux
    port map (
            O => \N__7526\,
            I => \N__7523\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__7523\,
            I => \N__7520\
        );

    \I__648\ : Odrv12
    port map (
            O => \N__7520\,
            I => rgb_c_2
        );

    \I__647\ : IoInMux
    port map (
            O => \N__7517\,
            I => \N__7514\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__7514\,
            I => \N__7511\
        );

    \I__645\ : Span4Mux_s2_h
    port map (
            O => \N__7511\,
            I => \N__7508\
        );

    \I__644\ : Span4Mux_h
    port map (
            O => \N__7508\,
            I => \N__7505\
        );

    \I__643\ : Span4Mux_v
    port map (
            O => \N__7505\,
            I => \N__7502\
        );

    \I__642\ : Odrv4
    port map (
            O => \N__7502\,
            I => rgb_c_5
        );

    \I__641\ : IoInMux
    port map (
            O => \N__7499\,
            I => \N__7496\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__7496\,
            I => \N__7493\
        );

    \I__639\ : IoSpan4Mux
    port map (
            O => \N__7493\,
            I => \N__7490\
        );

    \I__638\ : Span4Mux_s1_v
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__637\ : Span4Mux_v
    port map (
            O => \N__7487\,
            I => \N__7484\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__7484\,
            I => \this_vga_signals_M_hstate_q_i_4\
        );

    \I__635\ : IoInMux
    port map (
            O => \N__7481\,
            I => \N__7478\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__7478\,
            I => \N__7475\
        );

    \I__633\ : Span12Mux_s8_h
    port map (
            O => \N__7475\,
            I => \N__7472\
        );

    \I__632\ : Odrv12
    port map (
            O => \N__7472\,
            I => rgb_c_4
        );

    \I__631\ : IoInMux
    port map (
            O => \N__7469\,
            I => \N__7466\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__7466\,
            I => \N__7463\
        );

    \I__629\ : IoSpan4Mux
    port map (
            O => \N__7463\,
            I => \N__7460\
        );

    \I__628\ : IoSpan4Mux
    port map (
            O => \N__7460\,
            I => \N__7457\
        );

    \I__627\ : Span4Mux_s3_h
    port map (
            O => \N__7457\,
            I => \N__7454\
        );

    \I__626\ : Span4Mux_h
    port map (
            O => \N__7454\,
            I => \N__7451\
        );

    \I__625\ : Odrv4
    port map (
            O => \N__7451\,
            I => rgb_c_0
        );

    \I__624\ : InMux
    port map (
            O => \N__7448\,
            I => \N__7445\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__7445\,
            I => \N__7442\
        );

    \I__622\ : Odrv4
    port map (
            O => \N__7442\,
            I => m5
        );

    \I__621\ : IoInMux
    port map (
            O => \N__7439\,
            I => \N__7436\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__7436\,
            I => \N__7433\
        );

    \I__619\ : Span12Mux_s9_h
    port map (
            O => \N__7433\,
            I => \N__7430\
        );

    \I__618\ : Odrv12
    port map (
            O => \N__7430\,
            I => rgb_c_1
        );

    \I__617\ : IoInMux
    port map (
            O => \N__7427\,
            I => \N__7424\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__7424\,
            I => port_rw_c_i
        );

    \I__615\ : SRMux
    port map (
            O => \N__7421\,
            I => \N__7418\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__7418\,
            I => \N__7413\
        );

    \I__613\ : SRMux
    port map (
            O => \N__7417\,
            I => \N__7410\
        );

    \I__612\ : SRMux
    port map (
            O => \N__7416\,
            I => \N__7407\
        );

    \I__611\ : Span4Mux_v
    port map (
            O => \N__7413\,
            I => \N__7397\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__7410\,
            I => \N__7397\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__7407\,
            I => \N__7397\
        );

    \I__608\ : SRMux
    port map (
            O => \N__7406\,
            I => \N__7394\
        );

    \I__607\ : SRMux
    port map (
            O => \N__7405\,
            I => \N__7391\
        );

    \I__606\ : SRMux
    port map (
            O => \N__7404\,
            I => \N__7386\
        );

    \I__605\ : Span4Mux_v
    port map (
            O => \N__7397\,
            I => \N__7377\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__7394\,
            I => \N__7377\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__7391\,
            I => \N__7377\
        );

    \I__602\ : SRMux
    port map (
            O => \N__7390\,
            I => \N__7374\
        );

    \I__601\ : SRMux
    port map (
            O => \N__7389\,
            I => \N__7370\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__7386\,
            I => \N__7367\
        );

    \I__599\ : SRMux
    port map (
            O => \N__7385\,
            I => \N__7364\
        );

    \I__598\ : SRMux
    port map (
            O => \N__7384\,
            I => \N__7361\
        );

    \I__597\ : Span4Mux_v
    port map (
            O => \N__7377\,
            I => \N__7354\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__7374\,
            I => \N__7354\
        );

    \I__595\ : SRMux
    port map (
            O => \N__7373\,
            I => \N__7351\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__7370\,
            I => \N__7346\
        );

    \I__593\ : Span4Mux_s1_v
    port map (
            O => \N__7367\,
            I => \N__7339\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__7364\,
            I => \N__7339\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__7361\,
            I => \N__7339\
        );

    \I__590\ : SRMux
    port map (
            O => \N__7360\,
            I => \N__7336\
        );

    \I__589\ : SRMux
    port map (
            O => \N__7359\,
            I => \N__7333\
        );

    \I__588\ : Span4Mux_h
    port map (
            O => \N__7354\,
            I => \N__7324\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__7351\,
            I => \N__7324\
        );

    \I__586\ : SRMux
    port map (
            O => \N__7350\,
            I => \N__7321\
        );

    \I__585\ : SRMux
    port map (
            O => \N__7349\,
            I => \N__7317\
        );

    \I__584\ : Span4Mux_v
    port map (
            O => \N__7346\,
            I => \N__7305\
        );

    \I__583\ : Span4Mux_v
    port map (
            O => \N__7339\,
            I => \N__7305\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__7336\,
            I => \N__7305\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__7333\,
            I => \N__7305\
        );

    \I__580\ : SRMux
    port map (
            O => \N__7332\,
            I => \N__7302\
        );

    \I__579\ : SRMux
    port map (
            O => \N__7331\,
            I => \N__7299\
        );

    \I__578\ : IoInMux
    port map (
            O => \N__7330\,
            I => \N__7295\
        );

    \I__577\ : SRMux
    port map (
            O => \N__7329\,
            I => \N__7292\
        );

    \I__576\ : Span4Mux_v
    port map (
            O => \N__7324\,
            I => \N__7287\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__7321\,
            I => \N__7287\
        );

    \I__574\ : SRMux
    port map (
            O => \N__7320\,
            I => \N__7284\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__7317\,
            I => \N__7278\
        );

    \I__572\ : SRMux
    port map (
            O => \N__7316\,
            I => \N__7275\
        );

    \I__571\ : SRMux
    port map (
            O => \N__7315\,
            I => \N__7270\
        );

    \I__570\ : SRMux
    port map (
            O => \N__7314\,
            I => \N__7266\
        );

    \I__569\ : Span4Mux_v
    port map (
            O => \N__7305\,
            I => \N__7259\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__7302\,
            I => \N__7259\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__7299\,
            I => \N__7259\
        );

    \I__566\ : SRMux
    port map (
            O => \N__7298\,
            I => \N__7256\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__7295\,
            I => \N__7252\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__7292\,
            I => \N__7245\
        );

    \I__563\ : Span4Mux_h
    port map (
            O => \N__7287\,
            I => \N__7245\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__7284\,
            I => \N__7245\
        );

    \I__561\ : SRMux
    port map (
            O => \N__7283\,
            I => \N__7242\
        );

    \I__560\ : SRMux
    port map (
            O => \N__7282\,
            I => \N__7239\
        );

    \I__559\ : SRMux
    port map (
            O => \N__7281\,
            I => \N__7236\
        );

    \I__558\ : Span4Mux_v
    port map (
            O => \N__7278\,
            I => \N__7231\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__7275\,
            I => \N__7231\
        );

    \I__556\ : SRMux
    port map (
            O => \N__7274\,
            I => \N__7228\
        );

    \I__555\ : SRMux
    port map (
            O => \N__7273\,
            I => \N__7225\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__7270\,
            I => \N__7222\
        );

    \I__553\ : SRMux
    port map (
            O => \N__7269\,
            I => \N__7219\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__7266\,
            I => \N__7215\
        );

    \I__551\ : Span4Mux_v
    port map (
            O => \N__7259\,
            I => \N__7210\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__7256\,
            I => \N__7210\
        );

    \I__549\ : SRMux
    port map (
            O => \N__7255\,
            I => \N__7206\
        );

    \I__548\ : IoSpan4Mux
    port map (
            O => \N__7252\,
            I => \N__7203\
        );

    \I__547\ : Span4Mux_v
    port map (
            O => \N__7245\,
            I => \N__7198\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__7242\,
            I => \N__7198\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__7239\,
            I => \N__7195\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__7236\,
            I => \N__7192\
        );

    \I__543\ : Span4Mux_v
    port map (
            O => \N__7231\,
            I => \N__7185\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__7228\,
            I => \N__7185\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__7225\,
            I => \N__7185\
        );

    \I__540\ : Span4Mux_v
    port map (
            O => \N__7222\,
            I => \N__7180\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__7219\,
            I => \N__7180\
        );

    \I__538\ : SRMux
    port map (
            O => \N__7218\,
            I => \N__7177\
        );

    \I__537\ : Span12Mux_h
    port map (
            O => \N__7215\,
            I => \N__7174\
        );

    \I__536\ : Span4Mux_v
    port map (
            O => \N__7210\,
            I => \N__7171\
        );

    \I__535\ : SRMux
    port map (
            O => \N__7209\,
            I => \N__7168\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__7206\,
            I => \N__7165\
        );

    \I__533\ : Span4Mux_s2_h
    port map (
            O => \N__7203\,
            I => \N__7162\
        );

    \I__532\ : Span4Mux_h
    port map (
            O => \N__7198\,
            I => \N__7159\
        );

    \I__531\ : Span4Mux_s3_v
    port map (
            O => \N__7195\,
            I => \N__7156\
        );

    \I__530\ : Span4Mux_s3_v
    port map (
            O => \N__7192\,
            I => \N__7147\
        );

    \I__529\ : Span4Mux_v
    port map (
            O => \N__7185\,
            I => \N__7147\
        );

    \I__528\ : Span4Mux_s3_v
    port map (
            O => \N__7180\,
            I => \N__7147\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__7177\,
            I => \N__7147\
        );

    \I__526\ : Span12Mux_h
    port map (
            O => \N__7174\,
            I => \N__7144\
        );

    \I__525\ : Sp12to4
    port map (
            O => \N__7171\,
            I => \N__7139\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__7168\,
            I => \N__7139\
        );

    \I__523\ : Span12Mux_h
    port map (
            O => \N__7165\,
            I => \N__7136\
        );

    \I__522\ : Span4Mux_h
    port map (
            O => \N__7162\,
            I => \N__7133\
        );

    \I__521\ : Span4Mux_v
    port map (
            O => \N__7159\,
            I => \N__7126\
        );

    \I__520\ : Span4Mux_h
    port map (
            O => \N__7156\,
            I => \N__7126\
        );

    \I__519\ : Span4Mux_h
    port map (
            O => \N__7147\,
            I => \N__7126\
        );

    \I__518\ : Span12Mux_v
    port map (
            O => \N__7144\,
            I => \N__7123\
        );

    \I__517\ : Span12Mux_h
    port map (
            O => \N__7139\,
            I => \N__7120\
        );

    \I__516\ : Span12Mux_h
    port map (
            O => \N__7136\,
            I => \N__7115\
        );

    \I__515\ : Sp12to4
    port map (
            O => \N__7133\,
            I => \N__7115\
        );

    \I__514\ : Sp12to4
    port map (
            O => \N__7126\,
            I => \N__7112\
        );

    \I__513\ : Span12Mux_v
    port map (
            O => \N__7123\,
            I => \N__7109\
        );

    \I__512\ : Span12Mux_h
    port map (
            O => \N__7120\,
            I => \N__7104\
        );

    \I__511\ : Span12Mux_v
    port map (
            O => \N__7115\,
            I => \N__7104\
        );

    \I__510\ : Span12Mux_h
    port map (
            O => \N__7112\,
            I => \N__7101\
        );

    \I__509\ : Odrv12
    port map (
            O => \N__7109\,
            I => \CONSTANT_ONE_NET\
        );

    \I__508\ : Odrv12
    port map (
            O => \N__7104\,
            I => \CONSTANT_ONE_NET\
        );

    \I__507\ : Odrv12
    port map (
            O => \N__7101\,
            I => \CONSTANT_ONE_NET\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_10_cry_7\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_23_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_9_0_\
        );

    \IN_MUX_bfv_23_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vaddress_q_cry_7\,
            carryinitout => \bfn_23_10_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_haddress_q_cry_7\,
            carryinitout => \bfn_18_16_0_\
        );

    \this_vga_signals.M_vstate_q_RNI3M6M4_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8189\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_583_g\
        );

    \this_reset_cond.M_stage_q_RNI6VB7_3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19510\,
            GLOBALBUFFEROUTPUT => \N_631_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \port_data_rw_obuf_RNO_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18859\,
            lcout => port_rw_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNI1DID_1_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9833\,
            lcout => \this_vga_signals_M_hstate_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNIFPC1_1_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7903\,
            lcout => port_nmib_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_obuf_RNO_2_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7661\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7639\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_obuf_RNO_5_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7673\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7638\,
            lcout => rgb_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNI4GID_4_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8675\,
            lcout => \this_vga_signals_M_hstate_q_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_obuf_RNO_4_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7652\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7637\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_obuf_RNO_0_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000000000"
        )
    port map (
            in0 => \N__15566\,
            in1 => \N__11939\,
            in2 => \N__11458\,
            in3 => \N__7640\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m5_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__11940\,
            in1 => \N__15584\,
            in2 => \_gnd_net_\,
            in3 => \N__15856\,
            lcout => m5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_obuf_RNO_1_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__15865\,
            in1 => \N__7448\,
            in2 => \N__11495\,
            in3 => \N__7611\,
            lcout => rgb_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m22_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100001001111"
        )
    port map (
            in0 => \N__11941\,
            in1 => \N__15590\,
            in2 => \N__15869\,
            in3 => \N__11493\,
            lcout => \rgb_2_5_0__i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m10_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101001111"
        )
    port map (
            in0 => \N__15588\,
            in1 => \N__11958\,
            in2 => \N__15855\,
            in3 => \N__11485\,
            lcout => \rgb_2_5_0__i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNIG6VE_1_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9832\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7890\,
            lcout => rgb72,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m19_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100001011011"
        )
    port map (
            in0 => \N__15589\,
            in1 => \N__11962\,
            in2 => \N__15863\,
            in3 => \N__11492\,
            lcout => m19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_obuf_RNO_3_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__7621\,
            in1 => \N__7703\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rgb_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_1_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7562\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19139\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_last_q_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7763\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13168\,
            lcout => \this_start_data_delay_this_edge_detector_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19139\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_0_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__13167\,
            in1 => \N__7762\,
            in2 => \_gnd_net_\,
            in3 => \N__7732\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19139\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_3_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7709\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_0_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__13166\,
            in1 => \N__7761\,
            in2 => \_gnd_net_\,
            in3 => \N__7733\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_1_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7721\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_2_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7715\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m16_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100100011111"
        )
    port map (
            in0 => \N__15565\,
            in1 => \N__15864\,
            in2 => \N__11966\,
            in3 => \N__11494\,
            lcout => m16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_6_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7679\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_8_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7685\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_9_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7697\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_7_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7691\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_5_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7790\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_4_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7796\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19140\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_10_cry_0_c_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14099\,
            in2 => \N__8615\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_10_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_10_cry_0_THRU_LUT4_0_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8408\,
            in2 => \_gnd_net_\,
            in3 => \N__7784\,
            lcout => \this_vga_signals.un1_M_vcounter_q_10_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_10_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_10_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_10_cry_1_THRU_LUT4_0_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8372\,
            in2 => \_gnd_net_\,
            in3 => \N__7781\,
            lcout => \this_vga_signals.un1_M_vcounter_q_10_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_10_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_10_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_10_cry_2_THRU_LUT4_0_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8294\,
            in2 => \_gnd_net_\,
            in3 => \N__7778\,
            lcout => \this_vga_signals.un1_M_vcounter_q_10_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_10_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_10_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8329\,
            in2 => \_gnd_net_\,
            in3 => \N__7775\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_10_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_10_cry_4\,
            clk => \N__19153\,
            ce => 'H',
            sr => \N__17803\
        );

    \this_vga_signals.M_vcounter_q_5_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8076\,
            in2 => \_gnd_net_\,
            in3 => \N__7772\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_10_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_10_cry_5\,
            clk => \N__19153\,
            ce => 'H',
            sr => \N__17803\
        );

    \this_vga_signals.M_vcounter_q_6_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8045\,
            in2 => \_gnd_net_\,
            in3 => \N__7769\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_10_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_10_cry_6\,
            clk => \N__19153\,
            ce => 'H',
            sr => \N__17803\
        );

    \this_vga_signals.M_vcounter_q_7_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8581\,
            in2 => \_gnd_net_\,
            in3 => \N__7766\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_10_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_10_cry_7\,
            clk => \N__19153\,
            ce => 'H',
            sr => \N__17803\
        );

    \this_vga_signals.M_vcounter_q_8_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8536\,
            in2 => \_gnd_net_\,
            in3 => \N__7835\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_10_cry_8\,
            clk => \N__19160\,
            ce => 'H',
            sr => \N__17800\
        );

    \this_vga_signals.M_vcounter_q_9_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__8509\,
            in1 => \N__8096\,
            in2 => \N__8470\,
            in3 => \N__7832\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19160\,
            ce => 'H',
            sr => \N__17800\
        );

    \this_vga_signals.M_vcounter_q_3_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__8508\,
            in1 => \N__8295\,
            in2 => \N__8472\,
            in3 => \N__7829\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19160\,
            ce => 'H',
            sr => \N__17800\
        );

    \this_vga_signals.M_vcounter_q_2_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011101110000"
        )
    port map (
            in0 => \N__8476\,
            in1 => \N__8507\,
            in2 => \N__8378\,
            in3 => \N__7823\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19160\,
            ce => 'H',
            sr => \N__17800\
        );

    \this_vga_signals.M_vcounter_q_1_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__8506\,
            in1 => \N__8415\,
            in2 => \N__8471\,
            in3 => \N__7817\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19160\,
            ce => 'H',
            sr => \N__17800\
        );

    \this_vga_signals.M_vcounter_q_RNIHOM62_6_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__8330\,
            in1 => \N__8406\,
            in2 => \N__8053\,
            in3 => \N__7928\,
            lcout => \this_vga_signals.N_232_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIFUDD4_7_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7805\,
            in1 => \N__8534\,
            in2 => \N__7940\,
            in3 => \N__8584\,
            lcout => \this_vga_signals.N_238_0\,
            ltout => \this_vga_signals.N_238_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_1_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000010"
        )
    port map (
            in0 => \N__7879\,
            in1 => \N__19476\,
            in2 => \N__7811\,
            in3 => \N__7946\,
            lcout => port_nmib_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19164\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNILPDA1_9_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__8094\,
            in1 => \N__8077\,
            in2 => \_gnd_net_\,
            in3 => \N__8613\,
            lcout => \this_vga_signals.N_221_0\,
            ltout => \this_vga_signals.N_221_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIFUDD4_1_7_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8530\,
            in1 => \N__8582\,
            in2 => \N__7808\,
            in3 => \N__7804\,
            lcout => \this_vga_signals.N_237_0\,
            ltout => \this_vga_signals.N_237_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNO_0_1_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7949\,
            in3 => \N__8159\,
            lcout => \this_vga_signals.M_vstate_d_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIHQRK2_6_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8583\,
            in1 => \N__7936\,
            in2 => \N__8537\,
            in3 => \N__8049\,
            lcout => \this_vga_signals.N_226_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_3_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010101010"
        )
    port map (
            in0 => \N__8207\,
            in1 => \N__7844\,
            in2 => \N__19509\,
            in3 => \N__7919\,
            lcout => \this_vga_signals.M_vstate_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIV19S_2_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8296\,
            in2 => \_gnd_net_\,
            in3 => \N__8376\,
            lcout => \this_vga_signals.N_225_0\,
            ltout => \this_vga_signals.N_225_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIFUDD4_1_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8227\,
            in1 => \N__8331\,
            in2 => \N__7922\,
            in3 => \N__8417\,
            lcout => \this_vga_signals.N_239_0\,
            ltout => \this_vga_signals.N_239_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNO_0_2_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7843\,
            in2 => \N__7913\,
            in3 => \N__19479\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_258_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_2_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__19480\,
            in1 => \N__7880\,
            in2 => \N__7853\,
            in3 => \N__7850\,
            lcout => \this_vga_signals.M_vstate_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_7_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8009\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_2_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8021\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_6_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7985\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_3_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8003\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_4_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7997\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_5_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7991\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_14_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7979\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_11_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7955\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_13_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7967\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_12_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7973\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_10_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7961\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNI3M6M4_0_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__8154\,
            in1 => \N__19468\,
            in2 => \_gnd_net_\,
            in3 => \N__8174\,
            lcout => \this_vga_signals.M_vstate_q_RNI3M6M4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__8510\,
            in1 => \N__8612\,
            in2 => \N__8477\,
            in3 => \N__14100\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19147\,
            ce => 'H',
            sr => \N__17801\
        );

    \this_vga_signals.M_vstate_q_RNO_0_0_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8454\,
            in2 => \_gnd_net_\,
            in3 => \N__8502\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_251_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_0_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__19481\,
            in1 => \N__8158\,
            in2 => \N__8177\,
            in3 => \N__8173\,
            lcout => \this_vga_signals.M_vstate_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19154\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNIORO8_4_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__19474\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8113\,
            lcout => \this_vga_signals.M_vstate_q_srsts_0_a4_0_4\,
            ltout => \this_vga_signals.M_vstate_q_srsts_0_a4_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_5_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__8552\,
            in1 => \N__8423\,
            in2 => \N__8138\,
            in3 => \N__8231\,
            lcout => \this_vga_signals.M_vstate_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19161\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIU3IO1_2_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__8407\,
            in1 => \N__8290\,
            in2 => \N__8338\,
            in3 => \N__8371\,
            lcout => \this_vga_signals.N_230_0\,
            ltout => \this_vga_signals.N_230_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_4_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011101110"
        )
    port map (
            in0 => \N__8135\,
            in1 => \N__8258\,
            in2 => \N__8129\,
            in3 => \N__8230\,
            lcout => vsync_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19161\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI8EIO1_9_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__8095\,
            in1 => \N__8078\,
            in2 => \N__8054\,
            in3 => \N__8614\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vstate_q_srsts_0_o2_2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIFUDD4_0_7_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__8585\,
            in1 => \N__8551\,
            in2 => \N__8540\,
            in3 => \N__8535\,
            lcout => \this_vga_signals.N_248_0\,
            ltout => \this_vga_signals.N_248_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNO_0_5_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__19475\,
            in1 => \_gnd_net_\,
            in2 => \N__8480\,
            in3 => \N__8453\,
            lcout => \this_vga_signals.N_252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIU3IO1_0_2_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__8416\,
            in1 => \N__8377\,
            in2 => \N__8339\,
            in3 => \N__8297\,
            lcout => \this_vga_signals.M_vstate_q_srsts_0_o2_2_3\,
            ltout => \this_vga_signals.M_vstate_q_srsts_0_o2_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNO_0_4_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8242\,
            in1 => \N__19477\,
            in2 => \N__8261\,
            in3 => \N__8229\,
            lcout => \this_vga_signals.N_255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNO_0_3_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__8249\,
            in1 => \N__19478\,
            in2 => \N__8243\,
            in3 => \N__8228\,
            lcout => \this_vga_signals.N_256\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_8_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8201\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_11_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8195\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_10_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8633\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_12_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8645\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_9_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8639\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_15_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8627\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_0_5_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__19445\,
            in1 => \N__8837\,
            in2 => \_gnd_net_\,
            in3 => \N__8852\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_5_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__8693\,
            in1 => \N__8774\,
            in2 => \N__8621\,
            in3 => \N__8800\,
            lcout => \this_vga_signals.M_hstate_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI42JJ3_1_10_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8816\,
            in1 => \N__9521\,
            in2 => \N__8778\,
            in3 => \N__8956\,
            lcout => \this_vga_signals.N_398_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_16_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9425\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_0_2_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8972\,
            in1 => \N__8930\,
            in2 => \N__9824\,
            in3 => \N__19469\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_2_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__19470\,
            in1 => \N__8734\,
            in2 => \N__8618\,
            in3 => \N__8719\,
            lcout => \this_vga_signals.M_hstate_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIDR6I_0_7_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9572\,
            in2 => \_gnd_net_\,
            in3 => \N__9596\,
            lcout => \this_vga_signals.N_390_0\,
            ltout => \this_vga_signals.N_390_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI42JJ3_10_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9520\,
            in1 => \N__8955\,
            in2 => \N__8747\,
            in3 => \N__8815\,
            lcout => \this_vga_signals.N_397_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_0_4_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8743\,
            in1 => \N__19533\,
            in2 => \N__8707\,
            in3 => \N__8798\,
            lcout => \this_vga_signals.N_416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_0_3_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__8744\,
            in1 => \N__19534\,
            in2 => \N__8708\,
            in3 => \N__8799\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_3_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__19535\,
            in1 => \N__8735\,
            in2 => \N__8723\,
            in3 => \N__8720\,
            lcout => \this_vga_signals.M_hstate_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNIAFUK_4_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8662\,
            in2 => \_gnd_net_\,
            in3 => \N__19473\,
            lcout => \this_vga_signals.M_hstate_q_srsts_0_a3_0_4\,
            ltout => \this_vga_signals.M_hstate_q_srsts_0_a3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_4_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011111100"
        )
    port map (
            in0 => \N__8804\,
            in1 => \N__8684\,
            in2 => \N__8678\,
            in3 => \N__8780\,
            lcout => \this_vga_signals.M_hstate_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19155\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_13_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8651\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_0_1_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__8929\,
            in1 => \N__8971\,
            in2 => \N__9816\,
            in3 => \N__19376\,
            lcout => \this_vga_signals.N_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNI9J514_5_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8835\,
            in2 => \_gnd_net_\,
            in3 => \N__8850\,
            lcout => \this_vga_signals.M_hstate_d_0_sqmuxa\,
            ltout => \this_vga_signals.M_hstate_d_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_0_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__8870\,
            in1 => \N__8876\,
            in2 => \N__8879\,
            in3 => \N__19378\,
            lcout => \this_vga_signals.M_hstate_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI42JJ3_0_10_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8928\,
            in1 => \N__9524\,
            in2 => \N__8779\,
            in3 => \N__8957\,
            lcout => \this_vga_signals.N_405_0\,
            ltout => \this_vga_signals.N_405_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_1_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__19377\,
            in1 => \N__8869\,
            in2 => \N__8861\,
            in3 => \N__8858\,
            lcout => \this_vga_signals.M_hstate_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNIFIH84_5_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__8851\,
            in1 => \N__19375\,
            in2 => \_gnd_net_\,
            in3 => \N__8836\,
            lcout => \this_vga_signals.M_hstate_q_RNIFIH84Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9349\,
            in1 => \N__9364\,
            in2 => \N__9335\,
            in3 => \N__9381\,
            lcout => \this_vga_signals.M_hstate_q_srsts_0_o3_2_3_5\,
            ltout => \this_vga_signals.M_hstate_q_srsts_0_o3_2_3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9480\,
            in1 => \N__9409\,
            in2 => \N__8819\,
            in3 => \N__9315\,
            lcout => \this_vga_signals.N_385_0\,
            ltout => \this_vga_signals.N_385_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIN6C13_6_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__9295\,
            in1 => \N__9523\,
            in2 => \N__8807\,
            in3 => \N__9547\,
            lcout => \this_vga_signals.N_391_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIDR6I_7_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9570\,
            in2 => \_gnd_net_\,
            in3 => \N__9594\,
            lcout => \this_vga_signals.N_386_0\,
            ltout => \this_vga_signals.N_386_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIAIMG1_6_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9294\,
            in1 => \N__9522\,
            in2 => \N__8975\,
            in3 => \N__9546\,
            lcout => \this_vga_signals.M_hstate_q_srsts_0_o3_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIDR6I_6_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9545\,
            in2 => \_gnd_net_\,
            in3 => \N__9293\,
            lcout => \this_vga_signals.N_388_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIQFS22_0_11_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9410\,
            in1 => \N__9481\,
            in2 => \N__8939\,
            in3 => \N__9316\,
            lcout => \this_vga_signals.N_393_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_0_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9412\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19138\,
            ce => 'H',
            sr => \N__17795\
        );

    \this_vga_signals.M_hcounter_q_1_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__9413\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9385\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19138\,
            ce => 'H',
            sr => \N__17795\
        );

    \this_reset_cond.M_stage_q_2_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8908\,
            in2 => \_gnd_net_\,
            in3 => \N__8885\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8909\,
            in2 => \_gnd_net_\,
            in3 => \N__8915\,
            lcout => \M_this_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8906\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__8907\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8891\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g2_2_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15353\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12357\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g1_4_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__15124\,
            in1 => \N__14502\,
            in2 => \N__9113\,
            in3 => \N__12677\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g1_1_4_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9467\,
            in1 => \N__10274\,
            in2 => \N__9110\,
            in3 => \N__17658\,
            lcout => \this_vga_signals.g1_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g2_4_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12356\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15352\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g1_6_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__14501\,
            in1 => \N__15123\,
            in2 => \N__9107\,
            in3 => \N__11240\,
            lcout => \this_vga_signals.g1_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_14_N_8L16_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000001001"
        )
    port map (
            in0 => \N__9257\,
            in1 => \N__17662\,
            in2 => \N__11516\,
            in3 => \N__9263\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_14_N_8L16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_14_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011011110110"
        )
    port map (
            in0 => \N__12659\,
            in1 => \N__9104\,
            in2 => \N__9098\,
            in3 => \N__9683\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_c3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9620\,
            in1 => \N__9611\,
            in2 => \N__9095\,
            in3 => \N__9662\,
            lcout => this_vga_signals_un14_address_if_generate_plus_mult1_un75_sum_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_1_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011110001"
        )
    port map (
            in0 => \N__12362\,
            in1 => \N__12630\,
            in2 => \N__15389\,
            in3 => \N__14906\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_0_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011101100"
        )
    port map (
            in0 => \N__13963\,
            in1 => \N__11264\,
            in2 => \N__9266\,
            in3 => \N__14507\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_14_N_7L14_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011100001"
        )
    port map (
            in0 => \N__12363\,
            in1 => \N__12631\,
            in2 => \N__9605\,
            in3 => \N__9644\,
            lcout => \this_vga_signals.g0_14_N_7L14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m5_e_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__11699\,
            in1 => \_gnd_net_\,
            in2 => \N__11373\,
            in3 => \N__9248\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m5_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__19852\,
            in1 => \N__11366\,
            in2 => \N__9251\,
            in3 => \N__19904\,
            lcout => \this_vga_signals.if_i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_3_s_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11437\,
            in1 => \N__11408\,
            in2 => \_gnd_net_\,
            in3 => \N__19851\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_3_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axb1_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__10007\,
            in1 => \N__10202\,
            in2 => \_gnd_net_\,
            in3 => \N__10175\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1\,
            ltout => \this_vga_signals.mult1_un61_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m3_1_2_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11362\,
            in1 => \N__11430\,
            in2 => \N__9242\,
            in3 => \N__19850\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m3_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m5_i_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__11409\,
            in1 => \N__10031\,
            in2 => \N__9239\,
            in3 => \N__9749\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_6_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un75_sum_i_3_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__9236\,
            in1 => \N__9230\,
            in2 => \N__9224\,
            in3 => \N__9740\,
            lcout => this_vga_signals_un6_address_if_generate_plus_mult1_un75_sum_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m2_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000010100"
        )
    port map (
            in0 => \N__10874\,
            in1 => \N__9924\,
            in2 => \N__10000\,
            in3 => \N__10577\,
            lcout => \this_vga_signals.if_m2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m3_3_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__10578\,
            in1 => \N__9923\,
            in2 => \_gnd_net_\,
            in3 => \N__10873\,
            lcout => \this_vga_signals.if_i1_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10177\,
            in1 => \N__11677\,
            in2 => \N__10006\,
            in3 => \N__10204\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_c2_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101110001110"
        )
    port map (
            in0 => \N__9984\,
            in1 => \N__10203\,
            in2 => \N__11694\,
            in3 => \N__10176\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_14_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9275\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m3_0_0_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__13470\,
            in1 => \N__13659\,
            in2 => \_gnd_net_\,
            in3 => \N__13578\,
            lcout => \this_vga_signals.if_m3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_1_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011001110"
        )
    port map (
            in0 => \N__13657\,
            in1 => \N__13576\,
            in2 => \N__13503\,
            in3 => \N__13380\,
            lcout => \this_vga_signals.mult1_un40_sum_0_ac0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_2_1_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13575\,
            in2 => \_gnd_net_\,
            in3 => \N__13379\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_0_ac0_3_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_2_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110111"
        )
    port map (
            in0 => \N__10861\,
            in1 => \N__13483\,
            in2 => \N__9269\,
            in3 => \N__13658\,
            lcout => \this_vga_signals.mult1_un40_sum_0_ac0_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_0_a1_0_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13471\,
            in2 => \_gnd_net_\,
            in3 => \N__10860\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_0_ac0_3_0_a1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_ac0_3_0_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101111111"
        )
    port map (
            in0 => \N__13381\,
            in1 => \N__13656\,
            in2 => \N__9458\,
            in3 => \N__13577\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_0_ac0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m3_0_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__9455\,
            in1 => \N__9449\,
            in2 => \N__9443\,
            in3 => \N__9440\,
            lcout => \this_vga_signals.if_N_4_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_15_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9434\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19134\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9411\,
            in2 => \N__9389\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9365\,
            in2 => \_gnd_net_\,
            in3 => \N__9353\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__19142\,
            ce => 'H',
            sr => \N__17798\
        );

    \this_vga_signals.M_hcounter_q_3_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9350\,
            in2 => \_gnd_net_\,
            in3 => \N__9338\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__19142\,
            ce => 'H',
            sr => \N__17798\
        );

    \this_vga_signals.M_hcounter_q_4_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9334\,
            in2 => \_gnd_net_\,
            in3 => \N__9320\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__19142\,
            ce => 'H',
            sr => \N__17798\
        );

    \this_vga_signals.M_hcounter_q_5_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9317\,
            in2 => \_gnd_net_\,
            in3 => \N__9299\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \N__19142\,
            ce => 'H',
            sr => \N__17798\
        );

    \this_vga_signals.M_hcounter_q_6_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9296\,
            in2 => \_gnd_net_\,
            in3 => \N__9278\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \N__19142\,
            ce => 'H',
            sr => \N__17798\
        );

    \this_vga_signals.M_hcounter_q_7_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14082\,
            in1 => \N__9595\,
            in2 => \_gnd_net_\,
            in3 => \N__9575\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \N__19142\,
            ce => 'H',
            sr => \N__17798\
        );

    \this_vga_signals.M_hcounter_q_8_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9571\,
            in2 => \_gnd_net_\,
            in3 => \N__9551\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \N__19142\,
            ce => 'H',
            sr => \N__17798\
        );

    \this_vga_signals.M_hcounter_q_9_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9548\,
            in2 => \_gnd_net_\,
            in3 => \N__9527\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_9\,
            clk => \N__19149\,
            ce => 'H',
            sr => \N__17796\
        );

    \this_vga_signals.M_hcounter_q_10_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__14093\,
            in1 => \N__9506\,
            in2 => \_gnd_net_\,
            in3 => \N__9488\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_10\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_9\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_10\,
            clk => \N__19149\,
            ce => 'H',
            sr => \N__17796\
        );

    \this_vga_signals.M_hcounter_q_11_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__9482\,
            in1 => \N__14092\,
            in2 => \_gnd_net_\,
            in3 => \N__9485\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19149\,
            ce => 'H',
            sr => \N__17796\
        );

    \this_vga_signals.un14_address_g1_1_1_0_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13895\,
            in1 => \N__14027\,
            in2 => \_gnd_net_\,
            in3 => \N__15348\,
            lcout => \this_vga_signals.g1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g2_1_0_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15105\,
            in2 => \_gnd_net_\,
            in3 => \N__16369\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g2_3_0_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13894\,
            in1 => \N__14505\,
            in2 => \N__9461\,
            in3 => \N__15214\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g2_5_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001101001"
        )
    port map (
            in0 => \N__15347\,
            in1 => \N__12628\,
            in2 => \N__9638\,
            in3 => \N__12358\,
            lcout => \this_vga_signals.g2_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__17724\,
            in1 => \N__17683\,
            in2 => \_gnd_net_\,
            in3 => \N__17638\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_11_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__12620\,
            in1 => \N__12455\,
            in2 => \N__12427\,
            in3 => \N__12367\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_10_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111101000"
        )
    port map (
            in0 => \N__14500\,
            in1 => \N__13958\,
            in2 => \N__9635\,
            in3 => \N__10343\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_0_6_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17639\,
            in1 => \N__10280\,
            in2 => \N__9632\,
            in3 => \N__10289\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_1_0_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101111010010"
        )
    port map (
            in0 => \N__14036\,
            in1 => \N__13959\,
            in2 => \N__9629\,
            in3 => \N__9626\,
            lcout => \this_vga_signals.g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m5_1_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001100100"
        )
    port map (
            in0 => \N__14503\,
            in1 => \N__10734\,
            in2 => \N__13974\,
            in3 => \N__10349\,
            lcout => \this_vga_signals.mult1_un61_sum_c3\,
            ltout => \this_vga_signals.mult1_un61_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un68_sum_axb2_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17725\,
            in1 => \N__13960\,
            in2 => \N__9614\,
            in3 => \N__14504\,
            lcout => \this_vga_signals.mult1_un68_sum_axb2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_14_N_4L6_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15111\,
            in1 => \N__16370\,
            in2 => \N__13973\,
            in3 => \N__15215\,
            lcout => \this_vga_signals.g0_14_N_4L6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g1_2_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \N__10265\,
            in1 => \N__9704\,
            in2 => \N__9695\,
            in3 => \N__10775\,
            lcout => \this_vga_signals.g1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_RNI85LKP4_2_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011111100001"
        )
    port map (
            in0 => \N__17644\,
            in1 => \N__13965\,
            in2 => \N__10325\,
            in3 => \N__14498\,
            lcout => \this_vga_signals.M_vaddress_q_RNI85LKP4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_30_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001101001"
        )
    port map (
            in0 => \N__12629\,
            in1 => \N__15351\,
            in2 => \N__15125\,
            in3 => \N__12348\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_axb1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_33_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100001011110"
        )
    port map (
            in0 => \N__14506\,
            in1 => \N__13964\,
            in2 => \N__9677\,
            in3 => \N__10760\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c3_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_32_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9656\,
            in1 => \N__11015\,
            in2 => \N__9674\,
            in3 => \N__17643\,
            lcout => OPEN,
            ltout => \this_vga_signals.g3_0_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_17_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011001"
        )
    port map (
            in0 => \N__13975\,
            in1 => \N__9650\,
            in2 => \N__9671\,
            in3 => \N__9668\,
            lcout => \this_vga_signals.g2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_29_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010010101101"
        )
    port map (
            in0 => \N__15350\,
            in1 => \N__14497\,
            in2 => \N__10769\,
            in3 => \N__15117\,
            lcout => \this_vga_signals.g1_0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_0_x2_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17654\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14499\,
            lcout => \this_vga_signals.N_4_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_14_N_7L14_1_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101100110001"
        )
    port map (
            in0 => \N__15112\,
            in1 => \N__10331\,
            in2 => \N__14516\,
            in3 => \N__15349\,
            lcout => \this_vga_signals.g0_14_N_7L14_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m2_0_1_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__10702\,
            in1 => \N__9874\,
            in2 => \_gnd_net_\,
            in3 => \N__10883\,
            lcout => \this_vga_signals.if_m2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m2_0_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9755\,
            in1 => \N__19849\,
            in2 => \N__11701\,
            in3 => \N__9710\,
            lcout => \this_vga_signals.if_N_3_0_i\,
            ltout => \this_vga_signals.if_N_3_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m4_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010110000101"
        )
    port map (
            in0 => \N__11374\,
            in1 => \N__9839\,
            in2 => \N__9743\,
            in3 => \N__11413\,
            lcout => \this_vga_signals.mult1_un75_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m7_0_x4_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011010010011"
        )
    port map (
            in0 => \N__10882\,
            in1 => \N__10387\,
            in2 => \N__9940\,
            in3 => \N__10575\,
            lcout => \this_vga_signals.if_N_8_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_axbxc3_0_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10701\,
            in1 => \N__9734\,
            in2 => \N__10388\,
            in3 => \N__10522\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_3_1_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011111010100"
        )
    port map (
            in0 => \N__10524\,
            in1 => \N__10001\,
            in2 => \N__9941\,
            in3 => \N__10547\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_1_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_haddress_q_RNILVKM8_6_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__10576\,
            in1 => \N__9933\,
            in2 => \_gnd_net_\,
            in3 => \N__10881\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_haddress_q_RNILVKM8Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_ac0_3_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101101000111"
        )
    port map (
            in0 => \N__10523\,
            in1 => \N__9728\,
            in2 => \N__9722\,
            in3 => \N__10546\,
            lcout => \this_vga_signals.mult1_un54_sum_c3\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9719\,
            in3 => \N__10174\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_1_0_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110110010"
        )
    port map (
            in0 => \N__9991\,
            in1 => \N__9716\,
            in2 => \N__11698\,
            in3 => \N__9848\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_1_1_0\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10706\,
            in1 => \N__9878\,
            in2 => \N__9863\,
            in3 => \N__10867\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m3_2_ns_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10367\,
            in1 => \N__9860\,
            in2 => \_gnd_net_\,
            in3 => \N__10889\,
            lcout => \this_vga_signals_un6_address_if_N_5_mux_0\,
            ltout => \this_vga_signals_un6_address_if_N_5_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_ac0_3_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011101100"
        )
    port map (
            in0 => \N__9920\,
            in1 => \N__10383\,
            in2 => \N__9854\,
            in3 => \N__10866\,
            lcout => \this_vga_signals.mult1_un47_sum_c3\,
            ltout => \this_vga_signals.mult1_un47_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m1_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__10544\,
            in1 => \_gnd_net_\,
            in2 => \N__9851\,
            in3 => \N__9921\,
            lcout => \this_vga_signals.if_m1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axb1_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001110010100"
        )
    port map (
            in0 => \N__13673\,
            in1 => \N__13595\,
            in2 => \N__13515\,
            in3 => \N__13404\,
            lcout => \this_vga_signals.mult1_un40_sum_1_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10545\,
            in1 => \N__9922\,
            in2 => \N__10005\,
            in3 => \N__10525\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_0\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_m1_9_1_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9842\,
            in3 => \N__9995\,
            lcout => \this_vga_signals.if_m1_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_haddress_q_0_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9767\,
            in2 => \N__9831\,
            in3 => \N__9823\,
            lcout => \this_vga_signals.M_haddress_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \this_vga_signals.un1_M_haddress_q_cry_0\,
            clk => \N__19135\,
            ce => 'H',
            sr => \N__10252\
        );

    \this_vga_signals.M_haddress_q_1_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9761\,
            in2 => \_gnd_net_\,
            in3 => \N__10034\,
            lcout => \this_vga_signals.M_haddress_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_haddress_q_cry_0\,
            carryout => \this_vga_signals.un1_M_haddress_q_cry_1\,
            clk => \N__19135\,
            ce => 'H',
            sr => \N__10252\
        );

    \this_vga_signals.M_haddress_q_2_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10030\,
            in2 => \_gnd_net_\,
            in3 => \N__10016\,
            lcout => \this_vga_signals.M_haddress_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_haddress_q_cry_1\,
            carryout => \this_vga_signals.un1_M_haddress_q_cry_2\,
            clk => \N__19135\,
            ce => 'H',
            sr => \N__10252\
        );

    \this_vga_signals.M_haddress_q_3_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11361\,
            in2 => \_gnd_net_\,
            in3 => \N__10013\,
            lcout => \this_vga_signals.M_haddress_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_haddress_q_cry_2\,
            carryout => \this_vga_signals.un1_M_haddress_q_cry_3\,
            clk => \N__19135\,
            ce => 'H',
            sr => \N__10252\
        );

    \this_vga_signals.M_haddress_q_4_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11678\,
            in2 => \_gnd_net_\,
            in3 => \N__10010\,
            lcout => \this_vga_signals.M_haddress_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_haddress_q_cry_3\,
            carryout => \this_vga_signals.un1_M_haddress_q_cry_4\,
            clk => \N__19135\,
            ce => 'H',
            sr => \N__10252\
        );

    \this_vga_signals.M_haddress_q_5_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9999\,
            in2 => \_gnd_net_\,
            in3 => \N__9944\,
            lcout => \this_vga_signals.M_haddress_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_haddress_q_cry_4\,
            carryout => \this_vga_signals.un1_M_haddress_q_cry_5\,
            clk => \N__19135\,
            ce => 'H',
            sr => \N__10252\
        );

    \this_vga_signals.M_haddress_q_6_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9932\,
            in2 => \_gnd_net_\,
            in3 => \N__9890\,
            lcout => \this_vga_signals.M_haddress_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_haddress_q_cry_5\,
            carryout => \this_vga_signals.un1_M_haddress_q_cry_6\,
            clk => \N__19135\,
            ce => 'H',
            sr => \N__10252\
        );

    \this_vga_signals.M_haddress_q_7_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10878\,
            in2 => \_gnd_net_\,
            in3 => \N__9887\,
            lcout => \this_vga_signals.M_haddress_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_haddress_q_cry_6\,
            carryout => \this_vga_signals.un1_M_haddress_q_cry_7\,
            clk => \N__19135\,
            ce => 'H',
            sr => \N__10252\
        );

    \this_vga_signals.M_haddress_q_8_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13591\,
            in2 => \_gnd_net_\,
            in3 => \N__9884\,
            lcout => \this_vga_signals.M_haddress_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \this_vga_signals.un1_M_haddress_q_cry_8\,
            clk => \N__19143\,
            ce => 'H',
            sr => \N__10253\
        );

    \this_vga_signals.M_haddress_q_9_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13669\,
            in2 => \_gnd_net_\,
            in3 => \N__9881\,
            lcout => \this_vga_signals.M_haddress_qZ0Z_9\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_haddress_q_cry_8\,
            carryout => \this_vga_signals.un1_M_haddress_q_cry_9\,
            clk => \N__19143\,
            ce => 'H',
            sr => \N__10253\
        );

    \this_vga_signals.M_haddress_q_10_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13493\,
            in2 => \_gnd_net_\,
            in3 => \N__10259\,
            lcout => \this_vga_signals.M_haddress_qZ0Z_10\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_haddress_q_cry_9\,
            carryout => \this_vga_signals.un1_M_haddress_q_cry_10\,
            clk => \N__19143\,
            ce => 'H',
            sr => \N__10253\
        );

    \this_vga_signals.M_haddress_q_11_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13398\,
            in2 => \_gnd_net_\,
            in3 => \N__10256\,
            lcout => \this_vga_signals.CO0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19143\,
            ce => 'H',
            sr => \N__10253\
        );

    \this_start_address_delay.this_delay.M_pipe_q_17_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10226\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19156\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_18_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10214\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19156\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un54_sum_i_3_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10208\,
            in2 => \_gnd_net_\,
            in3 => \N__10181\,
            lcout => this_vga_signals_un6_address_if_generate_plus_mult1_un54_sum_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m12_bm_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001011110"
        )
    port map (
            in0 => \N__10745\,
            in1 => \N__14030\,
            in2 => \N__10310\,
            in3 => \N__14476\,
            lcout => \this_vga_signals.if_m12_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m6_0_N_2L1_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__12398\,
            in1 => \N__12594\,
            in2 => \_gnd_net_\,
            in3 => \N__12353\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m6_0_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001000100100"
        )
    port map (
            in0 => \N__14494\,
            in1 => \N__14028\,
            in2 => \N__10040\,
            in3 => \N__12456\,
            lcout => \this_vga_signals.if_N_7\,
            ltout => \this_vga_signals.if_N_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m8_bm_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14495\,
            in2 => \N__10037\,
            in3 => \N__10743\,
            lcout => \this_vga_signals.if_m8_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m1_3_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100100110110"
        )
    port map (
            in0 => \N__12354\,
            in1 => \N__12399\,
            in2 => \N__12623\,
            in3 => \N__12457\,
            lcout => \this_vga_signals.if_m1_3\,
            ltout => \this_vga_signals.if_m1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m8_am_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111110110001"
        )
    port map (
            in0 => \N__14029\,
            in1 => \N__14496\,
            in2 => \N__10301\,
            in3 => \N__10744\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m8_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m13_ns_1_LC_19_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__13944\,
            in1 => \N__17720\,
            in2 => \N__10298\,
            in3 => \N__10295\,
            lcout => \this_vga_signals.if_m13_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g1_3_LC_19_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100010001"
        )
    port map (
            in0 => \N__13961\,
            in1 => \N__14493\,
            in2 => \_gnd_net_\,
            in3 => \N__17637\,
            lcout => \this_vga_signals.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_0_2_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001101001"
        )
    port map (
            in0 => \N__12312\,
            in1 => \N__11278\,
            in2 => \N__11294\,
            in3 => \N__12587\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_0_1_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101111000"
        )
    port map (
            in0 => \N__14492\,
            in1 => \N__10342\,
            in2 => \N__10283\,
            in3 => \N__11194\,
            lcout => \this_vga_signals.g0_0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g1_1_1_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010011001"
        )
    port map (
            in0 => \N__12311\,
            in1 => \N__12738\,
            in2 => \_gnd_net_\,
            in3 => \N__12586\,
            lcout => \this_vga_signals.g3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_39_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101001011110"
        )
    port map (
            in0 => \N__11239\,
            in1 => \N__13962\,
            in2 => \N__14515\,
            in3 => \N__11216\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010111101010"
        )
    port map (
            in0 => \N__11195\,
            in1 => \N__10733\,
            in2 => \N__14509\,
            in3 => \N__11279\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m5_0_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12737\,
            in1 => \N__12718\,
            in2 => \_gnd_net_\,
            in3 => \N__12699\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m1_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__12309\,
            in1 => \N__12412\,
            in2 => \N__10352\,
            in3 => \N__12585\,
            lcout => \this_vga_signals.if_m1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_19_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001101001"
        )
    port map (
            in0 => \N__12584\,
            in1 => \N__12454\,
            in2 => \N__12420\,
            in3 => \N__12310\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_26_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001100100"
        )
    port map (
            in0 => \N__14477\,
            in1 => \N__10732\,
            in2 => \N__13972\,
            in3 => \N__11201\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_12_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011001001"
        )
    port map (
            in0 => \N__12315\,
            in1 => \N__15090\,
            in2 => \N__12605\,
            in3 => \N__15328\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g1_N_2L1_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100101"
        )
    port map (
            in0 => \N__15089\,
            in1 => \N__12559\,
            in2 => \N__14510\,
            in3 => \N__12314\,
            lcout => \this_vga_signals.g1_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_RNI8GTIA1_4_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__12316\,
            in1 => \N__15329\,
            in2 => \N__15120\,
            in3 => \N__12598\,
            lcout => \this_vga_signals.G_5_0_x2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axb1_LC_19_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011100001"
        )
    port map (
            in0 => \N__12288\,
            in1 => \N__12558\,
            in2 => \N__15119\,
            in3 => \N__15322\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1\,
            ltout => \this_vga_signals.mult1_un54_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g2_3_LC_19_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10316\,
            in3 => \N__14481\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g1_0_1_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__13948\,
            in1 => \N__11277\,
            in2 => \N__10313\,
            in3 => \N__11193\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_0_0_LC_19_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__14032\,
            in1 => \N__17636\,
            in2 => \N__10784\,
            in3 => \N__10781\,
            lcout => \this_vga_signals.g0_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_29_1_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000100011"
        )
    port map (
            in0 => \N__12607\,
            in1 => \N__12317\,
            in2 => \N__14511\,
            in3 => \N__15093\,
            lcout => \this_vga_signals.g0_29_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_34_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__12318\,
            in1 => \N__11501\,
            in2 => \N__11252\,
            in3 => \N__12608\,
            lcout => \this_vga_signals.N_3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m12_am_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__14475\,
            in1 => \N__10754\,
            in2 => \_gnd_net_\,
            in3 => \N__10742\,
            lcout => \this_vga_signals.if_m12_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_m_2_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__10912\,
            in1 => \N__10369\,
            in2 => \_gnd_net_\,
            in3 => \N__10927\,
            lcout => \this_vga_signals.mult1_un40_sum_m_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111010100001"
        )
    port map (
            in0 => \N__10928\,
            in1 => \N__10370\,
            in2 => \N__10916\,
            in3 => \N__10579\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_0\,
            ltout => \this_vga_signals.mult1_un47_sum_axbxc3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un47_sum_i_3_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10529\,
            in3 => \N__10526\,
            lcout => this_vga_signals_un6_address_if_generate_plus_mult1_un47_sum_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_m_1_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111100010"
        )
    port map (
            in0 => \N__10940\,
            in1 => \N__10368\,
            in2 => \N__12833\,
            in3 => \N__10880\,
            lcout => \this_vga_signals.mult1_un40_sum_m_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_haddress_q_RNID85Q_11_LC_19_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13497\,
            in2 => \_gnd_net_\,
            in3 => \N__13402\,
            lcout => \this_vga_signals.CO1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_c2_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__10939\,
            in1 => \N__11003\,
            in2 => \_gnd_net_\,
            in3 => \N__10862\,
            lcout => \this_vga_signals.mult1_un40_sum_1_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc2_0_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011110011100"
        )
    port map (
            in0 => \N__13403\,
            in1 => \N__13677\,
            in2 => \N__13514\,
            in3 => \N__13599\,
            lcout => \this_vga_signals.mult1_un40_sum_1_axbxc2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a1_1_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__13651\,
            in1 => \N__13573\,
            in2 => \_gnd_net_\,
            in3 => \N__13382\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_0_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110101111"
        )
    port map (
            in0 => \N__10858\,
            in1 => \_gnd_net_\,
            in2 => \N__10904\,
            in3 => \N__13476\,
            lcout => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a4_LC_19_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__13652\,
            in1 => \N__10854\,
            in2 => \N__13502\,
            in3 => \N__13385\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_1_axbxc3_a4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__10859\,
            in1 => \N__13654\,
            in2 => \N__10901\,
            in3 => \N__13580\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__10790\,
            in1 => \N__10796\,
            in2 => \N__10898\,
            in3 => \N__10895\,
            lcout => \this_vga_signals.mult1_un40_sum1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a5_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__13383\,
            in1 => \N__13475\,
            in2 => \N__10879\,
            in3 => \N__13579\,
            lcout => \this_vga_signals.mult1_un40_sum_1_axbxc3_a5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_1_1_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101000010"
        )
    port map (
            in0 => \N__13653\,
            in1 => \N__13574\,
            in2 => \N__13501\,
            in3 => \N__13384\,
            lcout => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_1_ac0_2_LC_19_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100101"
        )
    port map (
            in0 => \N__13386\,
            in1 => \N__13655\,
            in2 => \N__13507\,
            in3 => \N__13581\,
            lcout => \this_vga_signals.mult1_un40_sum_1_ac0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_16_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10997\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19150\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_18_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10973\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19150\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_19_LC_19_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10985\,
            lcout => \M_this_start_data_delay_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19150\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_17_LC_19_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10979\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19150\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_o3_0_0_0_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__13045\,
            in1 => \N__19471\,
            in2 => \_gnd_net_\,
            in3 => \N__13184\,
            lcout => \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_o3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_5_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110001111"
        )
    port map (
            in0 => \N__11312\,
            in1 => \N__13046\,
            in2 => \N__10961\,
            in3 => \N__11390\,
            lcout => \M_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19157\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_o4_5_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010001"
        )
    port map (
            in0 => \N__17160\,
            in1 => \N__10967\,
            in2 => \N__13187\,
            in3 => \N__19531\,
            lcout => \this_start_data_delay.this_edge_detector.N_252_0\,
            ltout => \this_start_data_delay.this_edge_detector.N_252_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_0_0_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000110000"
        )
    port map (
            in0 => \N__13091\,
            in1 => \N__10952\,
            in2 => \N__10943\,
            in3 => \N__11389\,
            lcout => \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_19_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11180\,
            lcout => \M_this_start_address_delay_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a2_0_5_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__13185\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19511\,
            lcout => \this_start_data_delay.this_edge_detector.N_267\,
            ltout => \this_start_data_delay.this_edge_detector.N_267_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_4_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13094\,
            in2 => \N__11174\,
            in3 => \N__13062\,
            lcout => debug_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m13_ns_LC_19_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__11171\,
            in1 => \N__11156\,
            in2 => \N__13976\,
            in3 => \N__11135\,
            lcout => if_m13_ns,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_11_LC_20_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010011001"
        )
    port map (
            in0 => \N__15346\,
            in1 => \N__12627\,
            in2 => \_gnd_net_\,
            in3 => \N__12355\,
            lcout => \this_vram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_6_3_i_o3_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15046\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15345\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_9_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_4_2_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001101001"
        )
    port map (
            in0 => \N__11972\,
            in1 => \N__12593\,
            in2 => \N__11018\,
            in3 => \N__12352\,
            lcout => \this_vga_signals.g0_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000110001110"
        )
    port map (
            in0 => \N__15205\,
            in1 => \N__15045\,
            in2 => \N__16382\,
            in3 => \N__11897\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_x_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__15044\,
            in1 => \N__16378\,
            in2 => \_gnd_net_\,
            in3 => \N__15204\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1_1_x\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_44_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011100001"
        )
    port map (
            in0 => \N__12556\,
            in1 => \N__12285\,
            in2 => \N__15122\,
            in3 => \N__15297\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_0_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_ac0_3_d_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000010000"
        )
    port map (
            in0 => \N__16371\,
            in1 => \N__12804\,
            in2 => \N__15118\,
            in3 => \N__15179\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_d\,
            ltout => \this_vga_signals.mult1_un47_sum_ac0_3_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_37_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12286\,
            in2 => \N__11225\,
            in3 => \N__15298\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_36_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100001010101"
        )
    port map (
            in0 => \N__15082\,
            in1 => \N__14471\,
            in2 => \N__11222\,
            in3 => \N__12026\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_c3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_42_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000100011110"
        )
    port map (
            in0 => \N__12557\,
            in1 => \N__12287\,
            in2 => \N__11219\,
            in3 => \N__11903\,
            lcout => \this_vga_signals.N_3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_3_0_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__12284\,
            in1 => \N__11210\,
            in2 => \N__11896\,
            in3 => \N__12555\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_18_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011010010"
        )
    port map (
            in0 => \N__12739\,
            in1 => \N__12717\,
            in2 => \N__11204\,
            in3 => \N__12700\,
            lcout => \this_vga_signals.if_N_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_ac0_2_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__15100\,
            in1 => \N__15299\,
            in2 => \_gnd_net_\,
            in3 => \N__12289\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m2_3_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__14609\,
            in1 => \N__16347\,
            in2 => \_gnd_net_\,
            in3 => \N__15185\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\,
            ltout => \this_vga_signals.mult1_un47_sum_ac0_3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m1_0_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100101010110"
        )
    port map (
            in0 => \N__15186\,
            in1 => \N__12554\,
            in2 => \N__11297\,
            in3 => \N__12055\,
            lcout => \this_vga_signals.if_m1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m5_0_s_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001001000"
        )
    port map (
            in0 => \N__15083\,
            in1 => \N__16348\,
            in2 => \N__14508\,
            in3 => \N__15188\,
            lcout => \this_vga_signals.if_m5_0_s\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_0_4_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15085\,
            in2 => \_gnd_net_\,
            in3 => \N__15301\,
            lcout => \this_vga_signals.g0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_0_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__15084\,
            in1 => \N__16349\,
            in2 => \_gnd_net_\,
            in3 => \N__15187\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_axbxc3_1_2_0_0_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001101001"
        )
    port map (
            in0 => \N__12563\,
            in1 => \N__15300\,
            in2 => \N__11282\,
            in3 => \N__12290\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_1_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_9_LC_20_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001101001"
        )
    port map (
            in0 => \N__12291\,
            in1 => \N__15101\,
            in2 => \N__15333\,
            in3 => \N__12564\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_c2_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011011101"
        )
    port map (
            in0 => \N__15091\,
            in1 => \N__16365\,
            in2 => \_gnd_net_\,
            in3 => \N__15200\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_3_1_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12809\,
            in2 => \N__11255\,
            in3 => \N__12056\,
            lcout => \this_vga_signals.g0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_19_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011001"
        )
    port map (
            in0 => \N__15314\,
            in1 => \N__12606\,
            in2 => \_gnd_net_\,
            in3 => \N__12313\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_35_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100000110011"
        )
    port map (
            in0 => \N__14482\,
            in1 => \N__15092\,
            in2 => \N__11243\,
            in3 => \N__11981\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIMTEJ4_11_LC_20_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16187\,
            in1 => \N__15628\,
            in2 => \_gnd_net_\,
            in3 => \N__16778\,
            lcout => \M_this_vram_read_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_axbxc3_0_1_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__11438\,
            in1 => \N__11414\,
            in2 => \_gnd_net_\,
            in3 => \N__19908\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_o3_5_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12645\,
            in2 => \_gnd_net_\,
            in3 => \N__13208\,
            lcout => \this_start_data_delay.this_edge_detector.N_253_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_i_1_3_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__11700\,
            in1 => \N__19915\,
            in2 => \N__11378\,
            in3 => \N__19864\,
            lcout => \this_vga_signals.mult1_un68_sum_i_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_2_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__11849\,
            in1 => \N__11862\,
            in2 => \N__11812\,
            in3 => \N__11764\,
            lcout => OPEN,
            ltout => \this_start_data_delay.this_edge_detector.N_261_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_2_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__12646\,
            in1 => \N__13052\,
            in2 => \N__11327\,
            in3 => \N__19472\,
            lcout => \M_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_0_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000011001100"
        )
    port map (
            in0 => \N__11848\,
            in1 => \N__11324\,
            in2 => \N__11811\,
            in3 => \N__11765\,
            lcout => \M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_0_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14222\,
            in1 => \N__11318\,
            in2 => \N__18848\,
            in3 => \N__11311\,
            lcout => \this_start_data_delay.this_edge_detector.N_275\,
            ltout => \this_start_data_delay.this_edge_detector.N_275_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_1_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__11841\,
            in1 => \N__11807\,
            in2 => \N__11300\,
            in3 => \N__11863\,
            lcout => OPEN,
            ltout => \this_start_data_delay.this_edge_detector.N_263_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_1_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__13063\,
            in1 => \N__13213\,
            in2 => \N__11867\,
            in3 => \N__19519\,
            lcout => \M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19165\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_state_q_srsts_0_a4_0_3_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__11864\,
            in1 => \N__11842\,
            in2 => \N__11813\,
            in3 => \N__11763\,
            lcout => OPEN,
            ltout => \this_start_data_delay.this_edge_detector.N_259_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_3_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__19518\,
            in1 => \N__13092\,
            in2 => \N__11750\,
            in3 => \N__13064\,
            lcout => \M_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19165\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un68_sum_i_3_LC_20_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101111010100"
        )
    port map (
            in0 => \N__11747\,
            in1 => \N__11726\,
            in2 => \N__11714\,
            in3 => \N__11630\,
            lcout => this_vga_signals_un6_address_if_generate_plus_mult1_un68_sum_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_12_LC_21_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__12893\,
            in1 => \N__11995\,
            in2 => \_gnd_net_\,
            in3 => \N__15468\,
            lcout => \this_vram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_14_N_8L16_sx_LC_21_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14051\,
            in2 => \_gnd_net_\,
            in3 => \N__14031\,
            lcout => \this_vga_signals.g0_14_N_8L16_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a1_1_0_LC_21_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12994\,
            in3 => \N__12065\,
            lcout => \this_vga_signals.N_2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_LC_21_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12082\,
            in1 => \N__12044\,
            in2 => \_gnd_net_\,
            in3 => \N__12763\,
            lcout => \this_vga_signals.mult1_un40_sum1_3\,
            ltout => \this_vga_signals.mult1_un40_sum1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_4_0_LC_21_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000111100"
        )
    port map (
            in0 => \N__12892\,
            in1 => \N__16356\,
            in2 => \N__11975\,
            in3 => \N__15467\,
            lcout => \this_vga_signals.g0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIETEJ4_11_LC_21_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15611\,
            in1 => \N__16418\,
            in2 => \_gnd_net_\,
            in3 => \N__15998\,
            lcout => \M_this_vram_read_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_1_1_1_LC_21_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000001111"
        )
    port map (
            in0 => \N__12935\,
            in1 => \N__12920\,
            in2 => \N__12020\,
            in3 => \N__15459\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_3_2_LC_21_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__14749\,
            in1 => \N__11873\,
            in2 => \N__11906\,
            in3 => \N__12861\,
            lcout => \this_vga_signals.g0_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_axbxc3_1_1_1_LC_21_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001011010"
        )
    port map (
            in0 => \N__12015\,
            in1 => \N__12919\,
            in2 => \N__12808\,
            in3 => \N__15458\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_1_1_LC_21_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14707\,
            in2 => \_gnd_net_\,
            in3 => \N__12860\,
            lcout => \this_vga_signals.mult1_un40_sum_m_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_6_LC_21_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14593\,
            lcout => \this_vga_signals.M_vaddress_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19124\,
            ce => 'H',
            sr => \N__16240\
        );

    \this_vga_signals.M_vaddress_q_fast_6_LC_21_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14594\,
            lcout => \this_vga_signals.M_vaddress_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19124\,
            ce => 'H',
            sr => \N__16240\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_3_LC_21_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111111"
        )
    port map (
            in0 => \N__14831\,
            in1 => \N__12859\,
            in2 => \N__12782\,
            in3 => \N__11879\,
            lcout => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_3_2_1_LC_21_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100110011100"
        )
    port map (
            in0 => \N__16363\,
            in1 => \N__13706\,
            in2 => \N__15121\,
            in3 => \N__15189\,
            lcout => \this_vga_signals.g0_3_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_am_x_2_LC_21_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110001000"
        )
    port map (
            in0 => \N__13704\,
            in1 => \N__14753\,
            in2 => \_gnd_net_\,
            in3 => \N__12862\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_m_am_x_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_ns_2_LC_21_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000010100"
        )
    port map (
            in0 => \N__15456\,
            in1 => \N__13828\,
            in2 => \N__12059\,
            in3 => \N__12917\,
            lcout => \this_vga_signals.mult1_un40_sum_m_ns_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_x1_3_LC_21_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__15454\,
            in1 => \N__12043\,
            in2 => \N__12764\,
            in3 => \N__12881\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_m_x1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_ns_3_LC_21_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__12882\,
            in1 => \N__15455\,
            in2 => \N__12032\,
            in3 => \N__12083\,
            lcout => \this_vga_signals.mult1_un40_sum_m_ns_3\,
            ltout => \this_vga_signals.mult1_un40_sum_m_ns_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_21_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111000011"
        )
    port map (
            in0 => \N__12918\,
            in1 => \N__12019\,
            in2 => \N__12029\,
            in3 => \N__15457\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g1_3_i_o3_LC_21_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16364\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15190\,
            lcout => \this_vga_signals.N_6_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_am_2_LC_21_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000101111000"
        )
    port map (
            in0 => \N__13705\,
            in1 => \N__14754\,
            in2 => \N__13829\,
            in3 => \N__12863\,
            lcout => \this_vga_signals.mult1_un40_sum_m_am_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_28_LC_21_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001011010"
        )
    port map (
            in0 => \N__11999\,
            in1 => \N__12886\,
            in2 => \N__16377\,
            in3 => \N__15470\,
            lcout => \this_vga_signals.N_6_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_16_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001101001"
        )
    port map (
            in0 => \N__15321\,
            in1 => \N__12621\,
            in2 => \N__15113\,
            in3 => \N__12322\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_8_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12740\,
            in1 => \N__12719\,
            in2 => \_gnd_net_\,
            in3 => \N__12701\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_5_LC_21_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__12416\,
            in1 => \N__12622\,
            in2 => \N__12683\,
            in3 => \N__12323\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_15_LC_21_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111101000"
        )
    port map (
            in0 => \N__14448\,
            in1 => \N__13932\,
            in2 => \N__12680\,
            in3 => \N__12673\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_0_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__13065\,
            in1 => \N__12647\,
            in2 => \N__13186\,
            in3 => \N__13209\,
            lcout => \M_current_address_qZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un54_sum_i_3_LC_21_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__12632\,
            in1 => \N__12467\,
            in2 => \N__12431\,
            in3 => \N__12368\,
            lcout => this_vga_signals_un14_address_if_generate_plus_mult1_un54_sum_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_4_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001111"
        )
    port map (
            in0 => \N__13816\,
            in1 => \N__13748\,
            in2 => \N__12749\,
            in3 => \N__14672\,
            lcout => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_7_rep1_LC_22_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14566\,
            lcout => \this_vga_signals.M_vaddress_q_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19125\,
            ce => 'H',
            sr => \N__16241\
        );

    \this_vga_signals.M_vaddress_q_fast_7_LC_22_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14567\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vaddress_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19125\,
            ce => 'H',
            sr => \N__16241\
        );

    \this_vga_signals.M_vaddress_q_fast_9_LC_22_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14543\,
            lcout => \this_vga_signals.M_vaddress_q_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19125\,
            ce => 'H',
            sr => \N__16241\
        );

    \this_vga_signals.M_vaddress_q_7_LC_22_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14565\,
            lcout => \this_vga_signals.M_vaddress_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19125\,
            ce => 'H',
            sr => \N__16241\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un40_sum_0_axb1_LC_22_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001001101101"
        )
    port map (
            in0 => \N__13682\,
            in1 => \N__13604\,
            in2 => \N__13520\,
            in3 => \N__13409\,
            lcout => \this_vga_signals.mult1_un40_sum_0_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_fast_RNI08841_0_8_LC_22_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010001100001"
        )
    port map (
            in0 => \N__12961\,
            in1 => \N__12990\,
            in2 => \N__13761\,
            in3 => \N__13811\,
            lcout => \this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8\,
            ltout => \this_vga_signals.M_vaddress_q_fast_RNI08841_0Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_1_LC_22_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010011001"
        )
    port map (
            in0 => \N__12818\,
            in1 => \N__13703\,
            in2 => \N__12812\,
            in3 => \N__15453\,
            lcout => \this_vga_signals.mult1_un40_sum_m_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_2_0_LC_22_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000111"
        )
    port map (
            in0 => \N__12778\,
            in1 => \N__13004\,
            in2 => \N__12965\,
            in3 => \N__12989\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_5_2_LC_22_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011011011"
        )
    port map (
            in0 => \N__13747\,
            in1 => \N__13810\,
            in2 => \N__12767\,
            in3 => \N__15452\,
            lcout => \this_vga_signals.mult1_un40_sum_1_axbxc3_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_fast_RNIHLHA_8_LC_22_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12988\,
            in2 => \N__12964\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.CO1_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_fast_8_LC_22_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14528\,
            lcout => \this_vga_signals.M_vaddress_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19128\,
            ce => 'H',
            sr => \N__16238\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_1_axbxc3_a4_1_0_LC_22_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12963\,
            in3 => \N__13003\,
            lcout => \this_vga_signals.mult1_un40_sum_1_axbxc3_a4_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_fast_5_LC_22_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16401\,
            lcout => \this_vga_signals.M_vaddress_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19128\,
            ce => 'H',
            sr => \N__16238\
        );

    \this_vga_signals.M_vaddress_q_fast_RNI08841_8_LC_22_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111000011"
        )
    port map (
            in0 => \N__12995\,
            in1 => \N__13804\,
            in2 => \N__13763\,
            in3 => \N__12962\,
            lcout => \this_vga_signals.N_353_0\,
            ltout => \this_vga_signals.N_353_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_m_bm_2_LC_22_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111010000111"
        )
    port map (
            in0 => \N__12858\,
            in1 => \N__12934\,
            in2 => \N__12923\,
            in3 => \N__14723\,
            lcout => \this_vga_signals.mult1_un40_sum_m_bm_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_6_rep1_LC_22_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14592\,
            lcout => \this_vga_signals.M_vaddress_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19136\,
            ce => 'H',
            sr => \N__16236\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_3_LC_22_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011100011"
        )
    port map (
            in0 => \N__14800\,
            in1 => \N__14656\,
            in2 => \N__13815\,
            in3 => \N__13752\,
            lcout => \this_vga_signals.mult1_un40_sum_0_axbxc3_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_1_0_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001011100"
        )
    port map (
            in0 => \N__13809\,
            in1 => \N__14664\,
            in2 => \N__13762\,
            in3 => \N__12857\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_0_axbxc3_5_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un40_sum_0_axbxc3_5_LC_22_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110100000000"
        )
    port map (
            in0 => \N__14871\,
            in1 => \N__14828\,
            in2 => \N__12902\,
            in3 => \N__12899\,
            lcout => \this_vga_signals.mult1_un40_sum0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_9_LC_22_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14539\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.CO0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19136\,
            ce => 'H',
            sr => \N__16236\
        );

    \this_vga_signals.M_vaddress_q_5_rep1_LC_22_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16406\,
            lcout => \this_vga_signals.M_vaddress_q_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19136\,
            ce => 'H',
            sr => \N__16236\
        );

    \this_vga_signals.M_vaddress_q_7_rep1_RNI65F81_LC_22_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001001011"
        )
    port map (
            in0 => \N__14825\,
            in1 => \N__14660\,
            in2 => \N__13817\,
            in3 => \N__13760\,
            lcout => \this_vga_signals.N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_7_rep1_RNI65F81_0_LC_22_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110111000011"
        )
    port map (
            in0 => \N__13805\,
            in1 => \N__14824\,
            in2 => \N__14671\,
            in3 => \N__13759\,
            lcout => \this_vga_signals.N_15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_RNIA1HT_1_7_LC_22_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001010001001"
        )
    port map (
            in0 => \N__14872\,
            in1 => \N__14826\,
            in2 => \N__14756\,
            in3 => \N__14665\,
            lcout => \this_vga_signals.N_355_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_31_LC_22_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15000\,
            in1 => \N__16346\,
            in2 => \_gnd_net_\,
            in3 => \N__15191\,
            lcout => \this_vga_signals.N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_RNIA1HT_0_7_LC_22_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110010011011"
        )
    port map (
            in0 => \N__14873\,
            in1 => \N__14827\,
            in2 => \N__14755\,
            in3 => \N__14666\,
            lcout => \this_vga_signals.N_15_0_0\,
            ltout => \this_vga_signals.N_15_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_1_N_2L1_LC_22_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101011010"
        )
    port map (
            in0 => \N__14765\,
            in1 => \N__14894\,
            in2 => \N__13685\,
            in3 => \N__15469\,
            lcout => \this_vga_signals.g0_1_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_haddress_q_RNI8ARU_11_LC_22_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111001011000"
        )
    port map (
            in0 => \N__13678\,
            in1 => \N__13600\,
            in2 => \N__13516\,
            in3 => \N__13405\,
            lcout => \M_haddress_q_RNI8ARU_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_RNI4EAV_1_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__13066\,
            in1 => \N__17816\,
            in2 => \N__13180\,
            in3 => \N__13217\,
            lcout => \M_current_address_q_0_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_data_d_0_sqmuxa_0_a4_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__13165\,
            in1 => \N__13093\,
            in2 => \_gnd_net_\,
            in3 => \N__13067\,
            lcout => \M_current_data_d_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_6_0_wclke_3_LC_22_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__17348\,
            in1 => \N__16972\,
            in2 => \N__17297\,
            in3 => \N__17178\,
            lcout => \this_vram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_3_0_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__14261\,
            in1 => \N__14249\,
            in2 => \_gnd_net_\,
            in3 => \N__14237\,
            lcout => \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_data_q_1_LC_22_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__14126\,
            in1 => \N__19601\,
            in2 => \N__18032\,
            in3 => \N__19505\,
            lcout => \M_current_data_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_0_LC_23_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14050\,
            in2 => \N__14111\,
            in3 => \N__14110\,
            lcout => \this_vga_signals.M_vaddress_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_23_9_0_\,
            carryout => \this_vga_signals.un1_M_vaddress_q_cry_0\,
            clk => \N__19129\,
            ce => 'H',
            sr => \N__16239\
        );

    \this_vga_signals.M_vaddress_q_1_LC_23_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14020\,
            in2 => \_gnd_net_\,
            in3 => \N__13979\,
            lcout => \this_vga_signals.M_vaddress_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vaddress_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vaddress_q_cry_1\,
            clk => \N__19129\,
            ce => 'H',
            sr => \N__16239\
        );

    \this_vga_signals.M_vaddress_q_2_LC_23_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13878\,
            in2 => \_gnd_net_\,
            in3 => \N__13838\,
            lcout => \this_vga_signals.M_vaddress_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vaddress_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vaddress_q_cry_2\,
            clk => \N__19129\,
            ce => 'H',
            sr => \N__16239\
        );

    \this_vga_signals.M_vaddress_q_3_LC_23_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14339\,
            in2 => \_gnd_net_\,
            in3 => \N__13835\,
            lcout => \this_vga_signals.M_vaddress_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vaddress_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vaddress_q_cry_3\,
            clk => \N__19129\,
            ce => 'H',
            sr => \N__16239\
        );

    \this_vga_signals.M_vaddress_q_4_LC_23_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14999\,
            in2 => \_gnd_net_\,
            in3 => \N__13832\,
            lcout => \this_vga_signals.M_vaddress_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vaddress_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vaddress_q_cry_4\,
            clk => \N__19129\,
            ce => 'H',
            sr => \N__16239\
        );

    \this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKME_LC_23_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16345\,
            in2 => \_gnd_net_\,
            in3 => \N__14597\,
            lcout => \this_vga_signals.un1_M_vaddress_q_cry_4_c_RNIOKMEZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vaddress_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vaddress_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNE_LC_23_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14766\,
            in2 => \_gnd_net_\,
            in3 => \N__14570\,
            lcout => \this_vga_signals.un1_M_vaddress_q_cry_5_c_RNIQNNEZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vaddress_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vaddress_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vaddress_q_cry_6_c_RNISQOE_LC_23_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14870\,
            in2 => \_gnd_net_\,
            in3 => \N__14552\,
            lcout => \this_vga_signals.un1_M_vaddress_q_cry_6_c_RNISQOEZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vaddress_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vaddress_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPE_LC_23_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14823\,
            in2 => \_gnd_net_\,
            in3 => \N__14549\,
            lcout => \this_vga_signals.un1_M_vaddress_q_cry_7_c_RNIUTPEZ0\,
            ltout => OPEN,
            carryin => \bfn_23_10_0_\,
            carryout => \this_vga_signals.un1_M_vaddress_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01RE_LC_23_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14670\,
            in2 => \_gnd_net_\,
            in3 => \N__14546\,
            lcout => \this_vga_signals.un1_M_vaddress_q_cry_8_c_RNI01REZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_8_LC_23_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14527\,
            lcout => \this_vga_signals.M_vaddress_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19137\,
            ce => 'H',
            sr => \N__16237\
        );

    \this_vga_signals.un14_address_g0_i_0_LC_23_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000101000"
        )
    port map (
            in0 => \N__16309\,
            in1 => \N__15001\,
            in2 => \N__14436\,
            in3 => \N__15206\,
            lcout => \this_vga_signals.N_1253_0\,
            ltout => \this_vga_signals.N_1253_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_1_N_5L7_x1_LC_23_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__15397\,
            in1 => \N__15404\,
            in2 => \N__14288\,
            in3 => \N__15361\,
            lcout => \this_vga_signals.g0_1_N_5L7_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_RNIHQ4M_7_LC_23_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011011101"
        )
    port map (
            in0 => \N__14876\,
            in1 => \N__14822\,
            in2 => \_gnd_net_\,
            in3 => \N__14669\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_2_LC_23_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100000011110"
        )
    port map (
            in0 => \N__14757\,
            in1 => \N__16308\,
            in2 => \N__15488\,
            in3 => \N__15485\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_3520_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_7_LC_23_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__15479\,
            in1 => \N__14882\,
            in2 => \N__15473\,
            in3 => \N__15466\,
            lcout => \this_vga_signals.mult1_un40_sum_0_2\,
            ltout => \this_vga_signals.mult1_un40_sum_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_1_N_5L7_x0_LC_23_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101011010"
        )
    port map (
            in0 => \N__15398\,
            in1 => \N__15376\,
            in2 => \N__15365\,
            in3 => \N__15362\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_N_5L7_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_1_N_5L7_ns_LC_23_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15334\,
            in2 => \N__15224\,
            in3 => \N__15221\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_N_5L7_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g0_1_1_0_LC_23_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011100001"
        )
    port map (
            in0 => \N__15207\,
            in1 => \N__15064\,
            in2 => \N__14909\,
            in3 => \N__16310\,
            lcout => \this_vga_signals.g0_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_13_LC_23_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001000111101000"
        )
    port map (
            in0 => \N__14668\,
            in1 => \N__14875\,
            in2 => \N__14767\,
            in3 => \N__14830\,
            lcout => \this_vram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19151\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_g1_0_LC_23_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110111011"
        )
    port map (
            in0 => \N__16293\,
            in1 => \N__14758\,
            in2 => \_gnd_net_\,
            in3 => \N__14893\,
            lcout => \this_vga_signals.g1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un14_address_if_m6_LC_23_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010010100"
        )
    port map (
            in0 => \N__14874\,
            in1 => \N__14829\,
            in2 => \N__14768\,
            in3 => \N__14667\,
            lcout => \this_vga_signals.if_i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_23_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15632\,
            in1 => \N__16685\,
            in2 => \_gnd_net_\,
            in3 => \N__15926\,
            lcout => \M_this_vram_read_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_4_0_wclke_3_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__17330\,
            in1 => \N__16968\,
            in2 => \N__17284\,
            in3 => \N__17194\,
            lcout => \this_vram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_RNIBHE21_3_LC_23_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15779\,
            in2 => \_gnd_net_\,
            in3 => \N__17815\,
            lcout => \M_current_address_q_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_esr_0_LC_23_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18156\,
            lcout => \M_current_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19188\,
            ce => \N__18325\,
            sr => \N__17792\
        );

    \this_vram.mem_mem_1_0_RNISSK11_LC_24_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16519\,
            in1 => \N__15662\,
            in2 => \_gnd_net_\,
            in3 => \N__15644\,
            lcout => \this_vram.mem_mem_1_0_RNISSKZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI5OL72_0_12_LC_24_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16652\,
            in1 => \N__15638\,
            in2 => \_gnd_net_\,
            in3 => \N__16731\,
            lcout => OPEN,
            ltout => \this_vram.mem_N_109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIETEJ4_0_11_LC_24_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__15621\,
            in1 => \_gnd_net_\,
            in2 => \N__15593\,
            in3 => \N__15494\,
            lcout => \M_this_vram_read_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_RNIQOI11_LC_24_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15524\,
            in1 => \N__15512\,
            in2 => \_gnd_net_\,
            in3 => \N__16520\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_0_0_RNIQOIZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16034\,
            in2 => \N__15497\,
            in3 => \N__16730\,
            lcout => \this_vram.mem_N_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_RNIU0N11_LC_24_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__16513\,
            in1 => \_gnd_net_\,
            in2 => \N__16061\,
            in3 => \N__16052\,
            lcout => \this_vram.mem_mem_2_0_RNIU0NZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16512\,
            in1 => \N__16028\,
            in2 => \_gnd_net_\,
            in3 => \N__16016\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_1_0_RNISSK11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI5OL72_12_LC_24_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__16097\,
            in1 => \_gnd_net_\,
            in2 => \N__16001\,
            in3 => \N__16711\,
            lcout => \this_vram.mem_N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_1_RNISOI11_LC_24_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15989\,
            in1 => \N__15974\,
            in2 => \_gnd_net_\,
            in3 => \N__16506\,
            lcout => \this_vram.mem_mem_0_1_RNISOIZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_1_RNI01N11_LC_24_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16508\,
            in1 => \N__15962\,
            in2 => \_gnd_net_\,
            in3 => \N__15944\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_2_1_RNI01NZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15935\,
            in2 => \N__15929\,
            in3 => \N__16733\,
            lcout => \this_vram.mem_N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_RNIU0N11_0_LC_24_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15917\,
            in1 => \N__15902\,
            in2 => \_gnd_net_\,
            in3 => \N__16507\,
            lcout => \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_RNIQOI11_0_LC_24_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15896\,
            in1 => \N__15884\,
            in2 => \_gnd_net_\,
            in3 => \N__16505\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI1GH72_12_LC_24_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__16732\,
            in1 => \_gnd_net_\,
            in2 => \N__16427\,
            in3 => \N__16424\,
            lcout => \this_vram.mem_N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vaddress_q_5_LC_24_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16405\,
            lcout => \this_vga_signals.M_vaddress_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19152\,
            ce => 'H',
            sr => \N__16235\
        );

    \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16475\,
            in1 => \N__16214\,
            in2 => \_gnd_net_\,
            in3 => \N__16196\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_2_1_RNI01N11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI5GH72_12_LC_24_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16734\,
            in1 => \_gnd_net_\,
            in2 => \N__16190\,
            in3 => \N__16148\,
            lcout => \this_vram.mem_N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_1_RNISOI11_0_LC_24_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16175\,
            in1 => \N__16160\,
            in2 => \_gnd_net_\,
            in3 => \N__16474\,
            lcout => \this_vram.mem_mem_0_1_RNISOI11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_0_wclke_3_LC_24_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__17347\,
            in1 => \N__16973\,
            in2 => \N__17291\,
            in3 => \N__17218\,
            lcout => \this_vram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16478\,
            in1 => \N__16121\,
            in2 => \_gnd_net_\,
            in3 => \N__16103\,
            lcout => \this_vram.mem_mem_3_0_RNI05P11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16088\,
            in1 => \N__16073\,
            in2 => \_gnd_net_\,
            in3 => \N__16476\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_1_1_RNIUSK11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI9OL72_12_LC_24_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__16736\,
            in1 => \N__16553\,
            in2 => \N__16781\,
            in3 => \_gnd_net_\,
            lcout => \this_vram.mem_N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_1_RNIUSK11_LC_24_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16766\,
            in1 => \N__16751\,
            in2 => \_gnd_net_\,
            in3 => \N__16477\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_1_1_RNIUSKZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__16735\,
            in1 => \_gnd_net_\,
            in2 => \N__16688\,
            in3 => \N__16436\,
            lcout => \this_vram.mem_N_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_RNI05P11_LC_24_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16679\,
            in1 => \N__16667\,
            in2 => \_gnd_net_\,
            in3 => \N__16479\,
            lcout => \this_vram.mem_mem_3_0_RNI05PZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_wclke_3_LC_24_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__17345\,
            in1 => \N__16966\,
            in2 => \N__17289\,
            in3 => \N__17214\,
            lcout => \this_vram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_wclke_3_LC_24_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__17346\,
            in1 => \N__16967\,
            in2 => \N__17290\,
            in3 => \N__17215\,
            lcout => \this_vram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_wclke_3_LC_24_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__17344\,
            in1 => \N__16965\,
            in2 => \N__17288\,
            in3 => \N__17213\,
            lcout => \this_vram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_1_RNI25P11_0_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16577\,
            in1 => \N__16559\,
            in2 => \_gnd_net_\,
            in3 => \N__16514\,
            lcout => \this_vram.mem_mem_3_1_RNI25P11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_1_RNI25P11_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16544\,
            in1 => \N__16538\,
            in2 => \_gnd_net_\,
            in3 => \N__16515\,
            lcout => \this_vram.mem_mem_3_1_RNI25PZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_esr_13_LC_24_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17491\,
            lcout => \M_current_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19169\,
            ce => \N__17868\,
            sr => \N__17808\
        );

    \M_current_address_q_esr_6_LC_24_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17492\,
            lcout => \M_current_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19172\,
            ce => \N__18301\,
            sr => \N__17807\
        );

    \M_current_address_q_esr_12_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17101\,
            lcout => \M_current_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19175\,
            ce => \N__17869\,
            sr => \N__17806\
        );

    \this_vram.mem_mem_5_0_wclke_3_LC_24_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__17317\,
            in1 => \N__16954\,
            in2 => \N__17292\,
            in3 => \N__17216\,
            lcout => \this_vram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_7_0_wclke_3_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17318\,
            in1 => \N__16955\,
            in2 => \N__17293\,
            in3 => \N__17217\,
            lcout => \this_vram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_esr_5_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17108\,
            lcout => \M_current_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19178\,
            ce => \N__18316\,
            sr => \N__17805\
        );

    \M_current_address_q_esr_11_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16916\,
            lcout => \M_current_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19179\,
            ce => \N__17880\,
            sr => \N__17804\
        );

    \M_current_address_q_esr_4_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16912\,
            lcout => \M_current_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19182\,
            ce => \N__18317\,
            sr => \N__17802\
        );

    \M_current_address_q_esr_2_LC_24_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19730\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_current_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19183\,
            ce => \N__18318\,
            sr => \N__17799\
        );

    \M_current_address_q_esr_9_LC_24_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19723\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_current_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19186\,
            ce => \N__17881\,
            sr => \N__17797\
        );

    \M_current_data_q_0_LC_24_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__18554\,
            in1 => \N__19609\,
            in2 => \N__18173\,
            in3 => \N__19532\,
            lcout => \M_current_data_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19189\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_esr_1_LC_24_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18021\,
            lcout => \M_current_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19193\,
            ce => \N__18326\,
            sr => \N__17794\
        );

    \M_current_address_q_esr_3_LC_24_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19566\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_current_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19193\,
            ce => \N__18326\,
            sr => \N__17794\
        );

    \M_current_address_q_esr_10_LC_24_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19571\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_current_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19194\,
            ce => \N__17879\,
            sr => \N__17793\
        );

    \M_current_address_q_esr_7_LC_24_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18169\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_current_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19194\,
            ce => \N__17879\,
            sr => \N__17793\
        );

    \M_current_address_q_esr_8_LC_24_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18031\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_current_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19197\,
            ce => \N__17885\,
            sr => \N__17791\
        );

    \this_vga_signals.un14_address_if_generate_plus_mult1_un61_sum_i_3_LC_24_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17738\,
            in1 => \N__17699\,
            in2 => \_gnd_net_\,
            in3 => \N__17672\,
            lcout => this_vga_signals_un14_address_if_generate_plus_mult1_un61_sum_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un6_address_if_generate_plus_mult1_un61_sum_axbxc3_LC_24_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19922\,
            in2 => \_gnd_net_\,
            in3 => \N__19880\,
            lcout => this_vga_signals_un6_address_if_generate_plus_mult1_un61_sum_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_data_q_2_LC_26_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__19639\,
            in1 => \N__19613\,
            in2 => \N__19523\,
            in3 => \N__19722\,
            lcout => \M_current_data_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_data_q_3_LC_26_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__19220\,
            in1 => \N__19608\,
            in2 => \N__19570\,
            in3 => \N__19504\,
            lcout => \M_current_data_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19198\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_4_0_LC_32_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18917\,
            in1 => \N__18905\,
            in2 => \N__18884\,
            in3 => \N__18869\,
            lcout => \this_start_data_delay.this_edge_detector.M_state_q_srsts_i_a2_1_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
